magic
tech sky130A
magscale 1 2
timestamp 1655506426
<< obsli1 >>
rect 51104 505159 534800 650401
<< obsm1 >>
rect 566 3408 580414 700528
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 580778 703610
rect 572 536 580778 703464
rect 710 480 1590 536
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6374 536
rect 6598 480 7570 536
rect 7794 480 8674 536
rect 8898 480 9870 536
rect 10094 480 11066 536
rect 11290 480 12262 536
rect 12486 480 13458 536
rect 13682 480 14654 536
rect 14878 480 15850 536
rect 16074 480 16954 536
rect 17178 480 18150 536
rect 18374 480 19346 536
rect 19570 480 20542 536
rect 20766 480 21738 536
rect 21962 480 22934 536
rect 23158 480 24130 536
rect 24354 480 25234 536
rect 25458 480 26430 536
rect 26654 480 27626 536
rect 27850 480 28822 536
rect 29046 480 30018 536
rect 30242 480 31214 536
rect 31438 480 32318 536
rect 32542 480 33514 536
rect 33738 480 34710 536
rect 34934 480 35906 536
rect 36130 480 37102 536
rect 37326 480 38298 536
rect 38522 480 39494 536
rect 39718 480 40598 536
rect 40822 480 41794 536
rect 42018 480 42990 536
rect 43214 480 44186 536
rect 44410 480 45382 536
rect 45606 480 46578 536
rect 46802 480 47774 536
rect 47998 480 48878 536
rect 49102 480 50074 536
rect 50298 480 51270 536
rect 51494 480 52466 536
rect 52690 480 53662 536
rect 53886 480 54858 536
rect 55082 480 55962 536
rect 56186 480 57158 536
rect 57382 480 58354 536
rect 58578 480 59550 536
rect 59774 480 60746 536
rect 60970 480 61942 536
rect 62166 480 63138 536
rect 63362 480 64242 536
rect 64466 480 65438 536
rect 65662 480 66634 536
rect 66858 480 67830 536
rect 68054 480 69026 536
rect 69250 480 70222 536
rect 70446 480 71418 536
rect 71642 480 72522 536
rect 72746 480 73718 536
rect 73942 480 74914 536
rect 75138 480 76110 536
rect 76334 480 77306 536
rect 77530 480 78502 536
rect 78726 480 79606 536
rect 79830 480 80802 536
rect 81026 480 81998 536
rect 82222 480 83194 536
rect 83418 480 84390 536
rect 84614 480 85586 536
rect 85810 480 86782 536
rect 87006 480 87886 536
rect 88110 480 89082 536
rect 89306 480 90278 536
rect 90502 480 91474 536
rect 91698 480 92670 536
rect 92894 480 93866 536
rect 94090 480 95062 536
rect 95286 480 96166 536
rect 96390 480 97362 536
rect 97586 480 98558 536
rect 98782 480 99754 536
rect 99978 480 100950 536
rect 101174 480 102146 536
rect 102370 480 103250 536
rect 103474 480 104446 536
rect 104670 480 105642 536
rect 105866 480 106838 536
rect 107062 480 108034 536
rect 108258 480 109230 536
rect 109454 480 110426 536
rect 110650 480 111530 536
rect 111754 480 112726 536
rect 112950 480 113922 536
rect 114146 480 115118 536
rect 115342 480 116314 536
rect 116538 480 117510 536
rect 117734 480 118706 536
rect 118930 480 119810 536
rect 120034 480 121006 536
rect 121230 480 122202 536
rect 122426 480 123398 536
rect 123622 480 124594 536
rect 124818 480 125790 536
rect 126014 480 126894 536
rect 127118 480 128090 536
rect 128314 480 129286 536
rect 129510 480 130482 536
rect 130706 480 131678 536
rect 131902 480 132874 536
rect 133098 480 134070 536
rect 134294 480 135174 536
rect 135398 480 136370 536
rect 136594 480 137566 536
rect 137790 480 138762 536
rect 138986 480 139958 536
rect 140182 480 141154 536
rect 141378 480 142350 536
rect 142574 480 143454 536
rect 143678 480 144650 536
rect 144874 480 145846 536
rect 146070 480 147042 536
rect 147266 480 148238 536
rect 148462 480 149434 536
rect 149658 480 150538 536
rect 150762 480 151734 536
rect 151958 480 152930 536
rect 153154 480 154126 536
rect 154350 480 155322 536
rect 155546 480 156518 536
rect 156742 480 157714 536
rect 157938 480 158818 536
rect 159042 480 160014 536
rect 160238 480 161210 536
rect 161434 480 162406 536
rect 162630 480 163602 536
rect 163826 480 164798 536
rect 165022 480 165994 536
rect 166218 480 167098 536
rect 167322 480 168294 536
rect 168518 480 169490 536
rect 169714 480 170686 536
rect 170910 480 171882 536
rect 172106 480 173078 536
rect 173302 480 174182 536
rect 174406 480 175378 536
rect 175602 480 176574 536
rect 176798 480 177770 536
rect 177994 480 178966 536
rect 179190 480 180162 536
rect 180386 480 181358 536
rect 181582 480 182462 536
rect 182686 480 183658 536
rect 183882 480 184854 536
rect 185078 480 186050 536
rect 186274 480 187246 536
rect 187470 480 188442 536
rect 188666 480 189638 536
rect 189862 480 190742 536
rect 190966 480 191938 536
rect 192162 480 193134 536
rect 193358 480 194330 536
rect 194554 480 195526 536
rect 195750 480 196722 536
rect 196946 480 197826 536
rect 198050 480 199022 536
rect 199246 480 200218 536
rect 200442 480 201414 536
rect 201638 480 202610 536
rect 202834 480 203806 536
rect 204030 480 205002 536
rect 205226 480 206106 536
rect 206330 480 207302 536
rect 207526 480 208498 536
rect 208722 480 209694 536
rect 209918 480 210890 536
rect 211114 480 212086 536
rect 212310 480 213282 536
rect 213506 480 214386 536
rect 214610 480 215582 536
rect 215806 480 216778 536
rect 217002 480 217974 536
rect 218198 480 219170 536
rect 219394 480 220366 536
rect 220590 480 221470 536
rect 221694 480 222666 536
rect 222890 480 223862 536
rect 224086 480 225058 536
rect 225282 480 226254 536
rect 226478 480 227450 536
rect 227674 480 228646 536
rect 228870 480 229750 536
rect 229974 480 230946 536
rect 231170 480 232142 536
rect 232366 480 233338 536
rect 233562 480 234534 536
rect 234758 480 235730 536
rect 235954 480 236926 536
rect 237150 480 238030 536
rect 238254 480 239226 536
rect 239450 480 240422 536
rect 240646 480 241618 536
rect 241842 480 242814 536
rect 243038 480 244010 536
rect 244234 480 245114 536
rect 245338 480 246310 536
rect 246534 480 247506 536
rect 247730 480 248702 536
rect 248926 480 249898 536
rect 250122 480 251094 536
rect 251318 480 252290 536
rect 252514 480 253394 536
rect 253618 480 254590 536
rect 254814 480 255786 536
rect 256010 480 256982 536
rect 257206 480 258178 536
rect 258402 480 259374 536
rect 259598 480 260570 536
rect 260794 480 261674 536
rect 261898 480 262870 536
rect 263094 480 264066 536
rect 264290 480 265262 536
rect 265486 480 266458 536
rect 266682 480 267654 536
rect 267878 480 268758 536
rect 268982 480 269954 536
rect 270178 480 271150 536
rect 271374 480 272346 536
rect 272570 480 273542 536
rect 273766 480 274738 536
rect 274962 480 275934 536
rect 276158 480 277038 536
rect 277262 480 278234 536
rect 278458 480 279430 536
rect 279654 480 280626 536
rect 280850 480 281822 536
rect 282046 480 283018 536
rect 283242 480 284214 536
rect 284438 480 285318 536
rect 285542 480 286514 536
rect 286738 480 287710 536
rect 287934 480 288906 536
rect 289130 480 290102 536
rect 290326 480 291298 536
rect 291522 480 292494 536
rect 292718 480 293598 536
rect 293822 480 294794 536
rect 295018 480 295990 536
rect 296214 480 297186 536
rect 297410 480 298382 536
rect 298606 480 299578 536
rect 299802 480 300682 536
rect 300906 480 301878 536
rect 302102 480 303074 536
rect 303298 480 304270 536
rect 304494 480 305466 536
rect 305690 480 306662 536
rect 306886 480 307858 536
rect 308082 480 308962 536
rect 309186 480 310158 536
rect 310382 480 311354 536
rect 311578 480 312550 536
rect 312774 480 313746 536
rect 313970 480 314942 536
rect 315166 480 316138 536
rect 316362 480 317242 536
rect 317466 480 318438 536
rect 318662 480 319634 536
rect 319858 480 320830 536
rect 321054 480 322026 536
rect 322250 480 323222 536
rect 323446 480 324326 536
rect 324550 480 325522 536
rect 325746 480 326718 536
rect 326942 480 327914 536
rect 328138 480 329110 536
rect 329334 480 330306 536
rect 330530 480 331502 536
rect 331726 480 332606 536
rect 332830 480 333802 536
rect 334026 480 334998 536
rect 335222 480 336194 536
rect 336418 480 337390 536
rect 337614 480 338586 536
rect 338810 480 339782 536
rect 340006 480 340886 536
rect 341110 480 342082 536
rect 342306 480 343278 536
rect 343502 480 344474 536
rect 344698 480 345670 536
rect 345894 480 346866 536
rect 347090 480 347970 536
rect 348194 480 349166 536
rect 349390 480 350362 536
rect 350586 480 351558 536
rect 351782 480 352754 536
rect 352978 480 353950 536
rect 354174 480 355146 536
rect 355370 480 356250 536
rect 356474 480 357446 536
rect 357670 480 358642 536
rect 358866 480 359838 536
rect 360062 480 361034 536
rect 361258 480 362230 536
rect 362454 480 363426 536
rect 363650 480 364530 536
rect 364754 480 365726 536
rect 365950 480 366922 536
rect 367146 480 368118 536
rect 368342 480 369314 536
rect 369538 480 370510 536
rect 370734 480 371614 536
rect 371838 480 372810 536
rect 373034 480 374006 536
rect 374230 480 375202 536
rect 375426 480 376398 536
rect 376622 480 377594 536
rect 377818 480 378790 536
rect 379014 480 379894 536
rect 380118 480 381090 536
rect 381314 480 382286 536
rect 382510 480 383482 536
rect 383706 480 384678 536
rect 384902 480 385874 536
rect 386098 480 387070 536
rect 387294 480 388174 536
rect 388398 480 389370 536
rect 389594 480 390566 536
rect 390790 480 391762 536
rect 391986 480 392958 536
rect 393182 480 394154 536
rect 394378 480 395258 536
rect 395482 480 396454 536
rect 396678 480 397650 536
rect 397874 480 398846 536
rect 399070 480 400042 536
rect 400266 480 401238 536
rect 401462 480 402434 536
rect 402658 480 403538 536
rect 403762 480 404734 536
rect 404958 480 405930 536
rect 406154 480 407126 536
rect 407350 480 408322 536
rect 408546 480 409518 536
rect 409742 480 410714 536
rect 410938 480 411818 536
rect 412042 480 413014 536
rect 413238 480 414210 536
rect 414434 480 415406 536
rect 415630 480 416602 536
rect 416826 480 417798 536
rect 418022 480 418902 536
rect 419126 480 420098 536
rect 420322 480 421294 536
rect 421518 480 422490 536
rect 422714 480 423686 536
rect 423910 480 424882 536
rect 425106 480 426078 536
rect 426302 480 427182 536
rect 427406 480 428378 536
rect 428602 480 429574 536
rect 429798 480 430770 536
rect 430994 480 431966 536
rect 432190 480 433162 536
rect 433386 480 434358 536
rect 434582 480 435462 536
rect 435686 480 436658 536
rect 436882 480 437854 536
rect 438078 480 439050 536
rect 439274 480 440246 536
rect 440470 480 441442 536
rect 441666 480 442546 536
rect 442770 480 443742 536
rect 443966 480 444938 536
rect 445162 480 446134 536
rect 446358 480 447330 536
rect 447554 480 448526 536
rect 448750 480 449722 536
rect 449946 480 450826 536
rect 451050 480 452022 536
rect 452246 480 453218 536
rect 453442 480 454414 536
rect 454638 480 455610 536
rect 455834 480 456806 536
rect 457030 480 458002 536
rect 458226 480 459106 536
rect 459330 480 460302 536
rect 460526 480 461498 536
rect 461722 480 462694 536
rect 462918 480 463890 536
rect 464114 480 465086 536
rect 465310 480 466190 536
rect 466414 480 467386 536
rect 467610 480 468582 536
rect 468806 480 469778 536
rect 470002 480 470974 536
rect 471198 480 472170 536
rect 472394 480 473366 536
rect 473590 480 474470 536
rect 474694 480 475666 536
rect 475890 480 476862 536
rect 477086 480 478058 536
rect 478282 480 479254 536
rect 479478 480 480450 536
rect 480674 480 481646 536
rect 481870 480 482750 536
rect 482974 480 483946 536
rect 484170 480 485142 536
rect 485366 480 486338 536
rect 486562 480 487534 536
rect 487758 480 488730 536
rect 488954 480 489834 536
rect 490058 480 491030 536
rect 491254 480 492226 536
rect 492450 480 493422 536
rect 493646 480 494618 536
rect 494842 480 495814 536
rect 496038 480 497010 536
rect 497234 480 498114 536
rect 498338 480 499310 536
rect 499534 480 500506 536
rect 500730 480 501702 536
rect 501926 480 502898 536
rect 503122 480 504094 536
rect 504318 480 505290 536
rect 505514 480 506394 536
rect 506618 480 507590 536
rect 507814 480 508786 536
rect 509010 480 509982 536
rect 510206 480 511178 536
rect 511402 480 512374 536
rect 512598 480 513478 536
rect 513702 480 514674 536
rect 514898 480 515870 536
rect 516094 480 517066 536
rect 517290 480 518262 536
rect 518486 480 519458 536
rect 519682 480 520654 536
rect 520878 480 521758 536
rect 521982 480 522954 536
rect 523178 480 524150 536
rect 524374 480 525346 536
rect 525570 480 526542 536
rect 526766 480 527738 536
rect 527962 480 528934 536
rect 529158 480 530038 536
rect 530262 480 531234 536
rect 531458 480 532430 536
rect 532654 480 533626 536
rect 533850 480 534822 536
rect 535046 480 536018 536
rect 536242 480 537122 536
rect 537346 480 538318 536
rect 538542 480 539514 536
rect 539738 480 540710 536
rect 540934 480 541906 536
rect 542130 480 543102 536
rect 543326 480 544298 536
rect 544522 480 545402 536
rect 545626 480 546598 536
rect 546822 480 547794 536
rect 548018 480 548990 536
rect 549214 480 550186 536
rect 550410 480 551382 536
rect 551606 480 552578 536
rect 552802 480 553682 536
rect 553906 480 554878 536
rect 555102 480 556074 536
rect 556298 480 557270 536
rect 557494 480 558466 536
rect 558690 480 559662 536
rect 559886 480 560766 536
rect 560990 480 561962 536
rect 562186 480 563158 536
rect 563382 480 564354 536
rect 564578 480 565550 536
rect 565774 480 566746 536
rect 566970 480 567942 536
rect 568166 480 569046 536
rect 569270 480 570242 536
rect 570466 480 571438 536
rect 571662 480 572634 536
rect 572858 480 573830 536
rect 574054 480 575026 536
rect 575250 480 576222 536
rect 576446 480 577326 536
rect 577550 480 578522 536
rect 578746 480 579718 536
rect 579942 480 580778 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 560 684084 583520 684317
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19588 583440 19988
rect 480 19580 583520 19588
rect 560 19180 583520 19580
rect 480 6796 583520 19180
rect 480 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 480 3299 583520 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 -5734 9854 709670
rect 12294 -1894 12914 705830
rect 12954 -7654 13574 711590
rect 16014 -3814 16634 707750
rect 19734 -5734 20354 709670
rect 22794 -1894 23414 705830
rect 23454 -7654 24074 711590
rect 26514 -3814 27134 707750
rect 30234 -5734 30854 709670
rect 33294 -1894 33914 705830
rect 33954 -7654 34574 711590
rect 37014 -3814 37634 707750
rect 40734 -5734 41354 709670
rect 43794 -1894 44414 705830
rect 44454 -7654 45074 711590
rect 47514 653033 48134 707750
rect 51234 653033 51854 709670
rect 54294 653033 54914 705830
rect 54954 653033 55574 711590
rect 58014 653033 58634 707750
rect 61734 653033 62354 709670
rect 64794 653033 65414 705830
rect 65454 653033 66074 711590
rect 68514 653033 69134 707750
rect 72234 653033 72854 709670
rect 75294 653033 75914 705830
rect 75954 653033 76574 711590
rect 79014 653033 79634 707750
rect 82734 653033 83354 709670
rect 85794 653033 86414 705830
rect 86454 653033 87074 711590
rect 89514 653033 90134 707750
rect 93234 653033 93854 709670
rect 96294 653033 96914 705830
rect 96954 653033 97574 711590
rect 100014 653033 100634 707750
rect 103734 653033 104354 709670
rect 106794 653033 107414 705830
rect 107454 653033 108074 711590
rect 110514 653033 111134 707750
rect 114234 653033 114854 709670
rect 117294 653033 117914 705830
rect 117954 653033 118574 711590
rect 121014 653033 121634 707750
rect 124734 653033 125354 709670
rect 127794 653033 128414 705830
rect 128454 653033 129074 711590
rect 131514 653033 132134 707750
rect 135234 653033 135854 709670
rect 138294 653033 138914 705830
rect 138954 653033 139574 711590
rect 142014 653033 142634 707750
rect 145734 653033 146354 709670
rect 148794 653033 149414 705830
rect 149454 653033 150074 711590
rect 152514 653033 153134 707750
rect 156234 653033 156854 709670
rect 159294 653033 159914 705830
rect 159954 653033 160574 711590
rect 47514 465308 48134 538000
rect 51234 465308 51854 538000
rect 54294 465308 54914 538000
rect 54954 465308 55574 538000
rect 58014 465308 58634 538000
rect 61734 465308 62354 538000
rect 64794 465308 65414 538000
rect 65454 465308 66074 538000
rect 68514 465308 69134 538000
rect 72234 465308 72854 538000
rect 75294 465308 75914 538000
rect 75954 465308 76574 538000
rect 79014 465308 79634 538000
rect 82734 465308 83354 538000
rect 85794 465308 86414 538000
rect 86454 465308 87074 538000
rect 89514 465308 90134 538000
rect 93234 465308 93854 538000
rect 96294 465308 96914 538000
rect 96954 465308 97574 538000
rect 100014 465308 100634 538000
rect 103734 465308 104354 538000
rect 106794 465308 107414 538000
rect 107454 465308 108074 538000
rect 110514 465308 111134 538000
rect 114234 465308 114854 538000
rect 117294 465308 117914 538000
rect 117954 465308 118574 538000
rect 121014 465308 121634 538000
rect 124734 465308 125354 538000
rect 127794 465308 128414 538000
rect 128454 465308 129074 538000
rect 131514 465308 132134 538000
rect 135234 465308 135854 538000
rect 138294 465308 138914 538000
rect 138954 465308 139574 538000
rect 142014 465308 142634 538000
rect 145734 465308 146354 538000
rect 148794 465308 149414 538000
rect 149454 465308 150074 538000
rect 152514 465308 153134 538000
rect 156234 465308 156854 538000
rect 159294 465308 159914 538000
rect 159954 465308 160574 538000
rect 163014 465308 163634 707750
rect 166734 465308 167354 709670
rect 169794 465308 170414 705830
rect 170454 465308 171074 711590
rect 173514 465308 174134 707750
rect 177234 465308 177854 709670
rect 180294 465308 180914 705830
rect 180954 465308 181574 711590
rect 184014 465308 184634 707750
rect 187734 465308 188354 709670
rect 47514 355308 48134 378000
rect 51234 355308 51854 378000
rect 54294 355308 54914 378000
rect 54954 355308 55574 378000
rect 58014 355308 58634 378000
rect 61734 355308 62354 378000
rect 64794 355308 65414 378000
rect 65454 355308 66074 378000
rect 68514 355308 69134 378000
rect 72234 355308 72854 378000
rect 75294 355308 75914 378000
rect 75954 355308 76574 378000
rect 79014 355308 79634 378000
rect 82734 355308 83354 378000
rect 85794 355308 86414 378000
rect 86454 355308 87074 378000
rect 89514 355308 90134 378000
rect 93234 355308 93854 378000
rect 96294 355308 96914 378000
rect 96954 355308 97574 378000
rect 100014 355308 100634 378000
rect 103734 355308 104354 378000
rect 106794 355308 107414 378000
rect 107454 355308 108074 378000
rect 110514 355308 111134 378000
rect 114234 355308 114854 378000
rect 117294 355308 117914 378000
rect 117954 355308 118574 378000
rect 121014 355308 121634 378000
rect 124734 355308 125354 378000
rect 127794 355308 128414 378000
rect 128454 355308 129074 378000
rect 131514 355308 132134 378000
rect 135234 355308 135854 378000
rect 138294 355308 138914 378000
rect 138954 355308 139574 378000
rect 142014 355308 142634 378000
rect 145734 355308 146354 378000
rect 148794 355308 149414 378000
rect 149454 355308 150074 378000
rect 152514 355308 153134 378000
rect 156234 355308 156854 378000
rect 159294 355308 159914 378000
rect 159954 355308 160574 378000
rect 163014 355308 163634 378000
rect 166734 355308 167354 378000
rect 169794 355308 170414 378000
rect 170454 355308 171074 378000
rect 173514 355308 174134 378000
rect 177234 355308 177854 378000
rect 180294 355308 180914 378000
rect 180954 355308 181574 378000
rect 184014 355308 184634 378000
rect 187734 355308 188354 378000
rect 47514 245308 48134 268000
rect 51234 245308 51854 268000
rect 54294 245308 54914 268000
rect 54954 245308 55574 268000
rect 58014 245308 58634 268000
rect 61734 245308 62354 268000
rect 64794 245308 65414 268000
rect 65454 245308 66074 268000
rect 68514 245308 69134 268000
rect 72234 245308 72854 268000
rect 75294 245308 75914 268000
rect 75954 245308 76574 268000
rect 79014 245308 79634 268000
rect 82734 245308 83354 268000
rect 85794 245308 86414 268000
rect 86454 245308 87074 268000
rect 89514 245308 90134 268000
rect 93234 245308 93854 268000
rect 96294 245308 96914 268000
rect 96954 245308 97574 268000
rect 100014 245308 100634 268000
rect 103734 245308 104354 268000
rect 106794 245308 107414 268000
rect 107454 245308 108074 268000
rect 110514 245308 111134 268000
rect 114234 245308 114854 268000
rect 117294 245308 117914 268000
rect 117954 245308 118574 268000
rect 121014 245308 121634 268000
rect 124734 245308 125354 268000
rect 127794 245308 128414 268000
rect 128454 245308 129074 268000
rect 131514 245308 132134 268000
rect 135234 245308 135854 268000
rect 138294 245308 138914 268000
rect 138954 245308 139574 268000
rect 142014 245308 142634 268000
rect 145734 245308 146354 268000
rect 148794 245308 149414 268000
rect 149454 245308 150074 268000
rect 152514 245308 153134 268000
rect 156234 245308 156854 268000
rect 159294 245308 159914 268000
rect 159954 245308 160574 268000
rect 163014 245308 163634 268000
rect 166734 245308 167354 268000
rect 169794 245308 170414 268000
rect 170454 245308 171074 268000
rect 173514 245308 174134 268000
rect 177234 245308 177854 268000
rect 180294 245308 180914 268000
rect 180954 245308 181574 268000
rect 184014 245308 184634 268000
rect 187734 245308 188354 268000
rect 47514 135308 48134 158000
rect 51234 135308 51854 158000
rect 54294 135308 54914 158000
rect 54954 135308 55574 158000
rect 58014 135308 58634 158000
rect 61734 135308 62354 158000
rect 64794 135308 65414 158000
rect 65454 135308 66074 158000
rect 68514 135308 69134 158000
rect 72234 135308 72854 158000
rect 75294 135308 75914 158000
rect 75954 135308 76574 158000
rect 79014 135308 79634 158000
rect 82734 135308 83354 158000
rect 85794 135308 86414 158000
rect 86454 135308 87074 158000
rect 89514 135308 90134 158000
rect 93234 135308 93854 158000
rect 96294 135308 96914 158000
rect 96954 135308 97574 158000
rect 100014 135308 100634 158000
rect 103734 135308 104354 158000
rect 106794 135308 107414 158000
rect 107454 135308 108074 158000
rect 110514 135308 111134 158000
rect 114234 135308 114854 158000
rect 117294 135308 117914 158000
rect 117954 135308 118574 158000
rect 121014 135308 121634 158000
rect 124734 135308 125354 158000
rect 127794 135308 128414 158000
rect 128454 135308 129074 158000
rect 131514 135308 132134 158000
rect 135234 135308 135854 158000
rect 138294 135308 138914 158000
rect 138954 135308 139574 158000
rect 142014 135308 142634 158000
rect 145734 135308 146354 158000
rect 148794 135308 149414 158000
rect 149454 135308 150074 158000
rect 152514 135308 153134 158000
rect 156234 135308 156854 158000
rect 159294 135308 159914 158000
rect 159954 135308 160574 158000
rect 163014 135308 163634 158000
rect 166734 135308 167354 158000
rect 169794 135308 170414 158000
rect 170454 135308 171074 158000
rect 173514 135308 174134 158000
rect 177234 135308 177854 158000
rect 180294 135308 180914 158000
rect 180954 135308 181574 158000
rect 184014 135308 184634 158000
rect 187734 135308 188354 158000
rect 47514 -3814 48134 48000
rect 51234 -5734 51854 48000
rect 54294 -1894 54914 48000
rect 54954 -7654 55574 48000
rect 58014 -3814 58634 48000
rect 61734 -5734 62354 48000
rect 64794 -1894 65414 48000
rect 65454 -7654 66074 48000
rect 68514 -3814 69134 48000
rect 72234 -5734 72854 48000
rect 75294 -1894 75914 48000
rect 75954 -7654 76574 48000
rect 79014 -3814 79634 48000
rect 82734 -5734 83354 48000
rect 85794 -1894 86414 48000
rect 86454 -7654 87074 48000
rect 89514 -3814 90134 48000
rect 93234 -5734 93854 48000
rect 96294 -1894 96914 48000
rect 96954 -7654 97574 48000
rect 100014 -3814 100634 48000
rect 103734 -5734 104354 48000
rect 106794 -1894 107414 48000
rect 107454 -7654 108074 48000
rect 110514 -3814 111134 48000
rect 114234 -5734 114854 48000
rect 117294 -1894 117914 48000
rect 117954 -7654 118574 48000
rect 121014 -3814 121634 48000
rect 124734 -5734 125354 48000
rect 127794 -1894 128414 48000
rect 128454 -7654 129074 48000
rect 131514 -3814 132134 48000
rect 135234 -5734 135854 48000
rect 138294 -1894 138914 48000
rect 138954 -7654 139574 48000
rect 142014 -3814 142634 48000
rect 145734 -5734 146354 48000
rect 148794 -1894 149414 48000
rect 149454 -7654 150074 48000
rect 152514 -3814 153134 48000
rect 156234 -5734 156854 48000
rect 159294 -1894 159914 48000
rect 159954 -7654 160574 48000
rect 163014 -3814 163634 48000
rect 166734 -5734 167354 48000
rect 169794 -1894 170414 48000
rect 170454 -7654 171074 48000
rect 173514 -3814 174134 48000
rect 177234 -5734 177854 48000
rect 180294 -1894 180914 48000
rect 180954 -7654 181574 48000
rect 184014 -3814 184634 48000
rect 187734 -5734 188354 48000
rect 190794 -1894 191414 705830
rect 191454 -7654 192074 711590
rect 194514 -3814 195134 707750
rect 198234 -5734 198854 709670
rect 201294 -1894 201914 705830
rect 201954 -7654 202574 711590
rect 205014 -3814 205634 707750
rect 208734 652000 209354 709670
rect 211794 652000 212414 705830
rect 212454 652000 213074 711590
rect 215514 652000 216134 707750
rect 219234 652000 219854 709670
rect 222294 652000 222914 705830
rect 222954 652000 223574 711590
rect 226014 652000 226634 707750
rect 229734 652000 230354 709670
rect 232794 652000 233414 705830
rect 233454 652000 234074 711590
rect 236514 652000 237134 707750
rect 240234 652000 240854 709670
rect 243294 652000 243914 705830
rect 243954 652000 244574 711590
rect 247014 652000 247634 707750
rect 250734 652000 251354 709670
rect 253794 652000 254414 705830
rect 254454 652000 255074 711590
rect 257514 652000 258134 707750
rect 261234 652000 261854 709670
rect 264294 652000 264914 705830
rect 264954 652000 265574 711590
rect 268014 652000 268634 707750
rect 271734 652000 272354 709670
rect 274794 652000 275414 705830
rect 275454 652000 276074 711590
rect 278514 652000 279134 707750
rect 282234 652000 282854 709670
rect 285294 652000 285914 705830
rect 285954 652000 286574 711590
rect 289014 652000 289634 707750
rect 292734 652000 293354 709670
rect 295794 652000 296414 705830
rect 296454 652000 297074 711590
rect 299514 652000 300134 707750
rect 303234 652000 303854 709670
rect 306294 652000 306914 705830
rect 306954 652000 307574 711590
rect 310014 652000 310634 707750
rect 313734 652000 314354 709670
rect 316794 652000 317414 705830
rect 317454 652000 318074 711590
rect 320514 652000 321134 707750
rect 324234 652000 324854 709670
rect 327294 652000 327914 705830
rect 327954 652000 328574 711590
rect 331014 652000 331634 707750
rect 208734 -5734 209354 501000
rect 211794 -1894 212414 501000
rect 212454 -7654 213074 501000
rect 215514 -3814 216134 501000
rect 219234 -5734 219854 501000
rect 222294 -1894 222914 501000
rect 222954 465308 223574 501000
rect 226014 465308 226634 501000
rect 229734 465308 230354 501000
rect 232794 465308 233414 501000
rect 233454 465308 234074 501000
rect 236514 465308 237134 501000
rect 240234 465308 240854 501000
rect 243294 465308 243914 501000
rect 243954 465308 244574 501000
rect 247014 465308 247634 501000
rect 250734 465308 251354 501000
rect 253794 465308 254414 501000
rect 254454 465308 255074 501000
rect 257514 465308 258134 501000
rect 261234 465308 261854 501000
rect 264294 465308 264914 501000
rect 264954 465308 265574 501000
rect 268014 465308 268634 501000
rect 271734 465308 272354 501000
rect 274794 465308 275414 501000
rect 275454 465308 276074 501000
rect 278514 465308 279134 501000
rect 282234 465308 282854 501000
rect 285294 465308 285914 501000
rect 285954 465308 286574 501000
rect 289014 465308 289634 501000
rect 292734 465308 293354 501000
rect 295794 465308 296414 501000
rect 296454 465308 297074 501000
rect 299514 465308 300134 501000
rect 303234 465308 303854 501000
rect 306294 465308 306914 501000
rect 306954 465308 307574 501000
rect 310014 465308 310634 501000
rect 313734 465308 314354 501000
rect 316794 465308 317414 501000
rect 317454 465308 318074 501000
rect 320514 465308 321134 501000
rect 324234 465308 324854 501000
rect 327294 465308 327914 501000
rect 327954 465308 328574 501000
rect 331014 465308 331634 501000
rect 334734 465308 335354 709670
rect 337794 465308 338414 705830
rect 338454 465308 339074 711590
rect 341514 465308 342134 707750
rect 345234 465308 345854 709670
rect 348294 465308 348914 705830
rect 348954 465308 349574 711590
rect 352014 465308 352634 707750
rect 355734 465308 356354 709670
rect 358794 465308 359414 705830
rect 359454 465308 360074 711590
rect 362514 465308 363134 707750
rect 222954 355308 223574 378000
rect 226014 355308 226634 378000
rect 229734 355308 230354 378000
rect 232794 355308 233414 378000
rect 233454 355308 234074 378000
rect 236514 355308 237134 378000
rect 240234 355308 240854 378000
rect 243294 355308 243914 378000
rect 243954 355308 244574 378000
rect 247014 355308 247634 378000
rect 250734 355308 251354 378000
rect 253794 355308 254414 378000
rect 254454 355308 255074 378000
rect 257514 355308 258134 378000
rect 261234 355308 261854 378000
rect 264294 355308 264914 378000
rect 264954 355308 265574 378000
rect 268014 355308 268634 378000
rect 271734 355308 272354 378000
rect 274794 355308 275414 378000
rect 275454 355308 276074 378000
rect 278514 355308 279134 378000
rect 282234 355308 282854 378000
rect 285294 355308 285914 378000
rect 285954 355308 286574 378000
rect 289014 355308 289634 378000
rect 292734 355308 293354 378000
rect 295794 355308 296414 378000
rect 296454 355308 297074 378000
rect 299514 355308 300134 378000
rect 303234 355308 303854 378000
rect 306294 355308 306914 378000
rect 306954 355308 307574 378000
rect 310014 355308 310634 378000
rect 313734 355308 314354 378000
rect 316794 355308 317414 378000
rect 317454 355308 318074 378000
rect 320514 355308 321134 378000
rect 324234 355308 324854 378000
rect 327294 355308 327914 378000
rect 327954 355308 328574 378000
rect 331014 355308 331634 378000
rect 334734 355308 335354 378000
rect 337794 355308 338414 378000
rect 338454 355308 339074 378000
rect 341514 355308 342134 378000
rect 345234 355308 345854 378000
rect 348294 355308 348914 378000
rect 348954 355308 349574 378000
rect 352014 355308 352634 378000
rect 355734 355308 356354 378000
rect 358794 355308 359414 378000
rect 359454 355308 360074 378000
rect 362514 355308 363134 378000
rect 222954 245308 223574 268000
rect 226014 245308 226634 268000
rect 229734 245308 230354 268000
rect 232794 245308 233414 268000
rect 233454 245308 234074 268000
rect 236514 245308 237134 268000
rect 240234 245308 240854 268000
rect 243294 245308 243914 268000
rect 243954 245308 244574 268000
rect 247014 245308 247634 268000
rect 250734 245308 251354 268000
rect 253794 245308 254414 268000
rect 254454 245308 255074 268000
rect 257514 245308 258134 268000
rect 261234 245308 261854 268000
rect 264294 245308 264914 268000
rect 264954 245308 265574 268000
rect 268014 245308 268634 268000
rect 271734 245308 272354 268000
rect 274794 245308 275414 268000
rect 275454 245308 276074 268000
rect 278514 245308 279134 268000
rect 282234 245308 282854 268000
rect 285294 245308 285914 268000
rect 285954 245308 286574 268000
rect 289014 245308 289634 268000
rect 292734 245308 293354 268000
rect 295794 245308 296414 268000
rect 296454 245308 297074 268000
rect 299514 245308 300134 268000
rect 303234 245308 303854 268000
rect 306294 245308 306914 268000
rect 306954 245308 307574 268000
rect 310014 245308 310634 268000
rect 313734 245308 314354 268000
rect 316794 245308 317414 268000
rect 317454 245308 318074 268000
rect 320514 245308 321134 268000
rect 324234 245308 324854 268000
rect 327294 245308 327914 268000
rect 327954 245308 328574 268000
rect 331014 245308 331634 268000
rect 334734 245308 335354 268000
rect 337794 245308 338414 268000
rect 338454 245308 339074 268000
rect 341514 245308 342134 268000
rect 345234 245308 345854 268000
rect 348294 245308 348914 268000
rect 348954 245308 349574 268000
rect 352014 245308 352634 268000
rect 355734 245308 356354 268000
rect 358794 245308 359414 268000
rect 359454 245308 360074 268000
rect 362514 245308 363134 268000
rect 222954 135308 223574 158000
rect 226014 135308 226634 158000
rect 229734 135308 230354 158000
rect 232794 135308 233414 158000
rect 233454 135308 234074 158000
rect 236514 135308 237134 158000
rect 240234 135308 240854 158000
rect 243294 135308 243914 158000
rect 243954 135308 244574 158000
rect 247014 135308 247634 158000
rect 250734 135308 251354 158000
rect 253794 135308 254414 158000
rect 254454 135308 255074 158000
rect 257514 135308 258134 158000
rect 261234 135308 261854 158000
rect 264294 135308 264914 158000
rect 264954 135308 265574 158000
rect 268014 135308 268634 158000
rect 271734 135308 272354 158000
rect 274794 135308 275414 158000
rect 275454 135308 276074 158000
rect 278514 135308 279134 158000
rect 282234 135308 282854 158000
rect 285294 135308 285914 158000
rect 285954 135308 286574 158000
rect 289014 135308 289634 158000
rect 292734 135308 293354 158000
rect 295794 135308 296414 158000
rect 296454 135308 297074 158000
rect 299514 135308 300134 158000
rect 303234 135308 303854 158000
rect 306294 135308 306914 158000
rect 306954 135308 307574 158000
rect 310014 135308 310634 158000
rect 313734 135308 314354 158000
rect 316794 135308 317414 158000
rect 317454 135308 318074 158000
rect 320514 135308 321134 158000
rect 324234 135308 324854 158000
rect 327294 135308 327914 158000
rect 327954 135308 328574 158000
rect 331014 135308 331634 158000
rect 334734 135308 335354 158000
rect 337794 135308 338414 158000
rect 338454 135308 339074 158000
rect 341514 135308 342134 158000
rect 345234 135308 345854 158000
rect 348294 135308 348914 158000
rect 348954 135308 349574 158000
rect 352014 135308 352634 158000
rect 355734 135308 356354 158000
rect 358794 135308 359414 158000
rect 359454 135308 360074 158000
rect 362514 135308 363134 158000
rect 222954 -7654 223574 48000
rect 226014 -3814 226634 48000
rect 229734 -5734 230354 48000
rect 232794 -1894 233414 48000
rect 233454 -7654 234074 48000
rect 236514 -3814 237134 48000
rect 240234 -5734 240854 48000
rect 243294 -1894 243914 48000
rect 243954 -7654 244574 48000
rect 247014 -3814 247634 48000
rect 250734 -5734 251354 48000
rect 253794 -1894 254414 48000
rect 254454 -7654 255074 48000
rect 257514 -3814 258134 48000
rect 261234 -5734 261854 48000
rect 264294 -1894 264914 48000
rect 264954 -7654 265574 48000
rect 268014 -3814 268634 48000
rect 271734 -5734 272354 48000
rect 274794 -1894 275414 48000
rect 275454 -7654 276074 48000
rect 278514 -3814 279134 48000
rect 282234 -5734 282854 48000
rect 285294 -1894 285914 48000
rect 285954 -7654 286574 48000
rect 289014 -3814 289634 48000
rect 292734 -5734 293354 48000
rect 295794 -1894 296414 48000
rect 296454 -7654 297074 48000
rect 299514 -3814 300134 48000
rect 303234 -5734 303854 48000
rect 306294 -1894 306914 48000
rect 306954 -7654 307574 48000
rect 310014 -3814 310634 48000
rect 313734 -5734 314354 48000
rect 316794 -1894 317414 48000
rect 317454 -7654 318074 48000
rect 320514 -3814 321134 48000
rect 324234 -5734 324854 48000
rect 327294 -1894 327914 48000
rect 327954 -7654 328574 48000
rect 331014 -3814 331634 48000
rect 334734 -5734 335354 48000
rect 337794 -1894 338414 48000
rect 338454 -7654 339074 48000
rect 341514 -3814 342134 48000
rect 345234 -5734 345854 48000
rect 348294 -1894 348914 48000
rect 348954 -7654 349574 48000
rect 352014 -3814 352634 48000
rect 355734 -5734 356354 48000
rect 358794 -1894 359414 48000
rect 359454 -7654 360074 48000
rect 362514 -3814 363134 48000
rect 366234 -5734 366854 709670
rect 369294 -1894 369914 705830
rect 369954 -7654 370574 711590
rect 373014 -3814 373634 707750
rect 376734 -5734 377354 709670
rect 379794 655099 380414 705830
rect 380454 655099 381074 711590
rect 383514 655099 384134 707750
rect 387234 655099 387854 709670
rect 390294 655099 390914 705830
rect 390954 655099 391574 711590
rect 394014 655099 394634 707750
rect 397734 655099 398354 709670
rect 400794 655099 401414 705830
rect 401454 655099 402074 711590
rect 404514 655099 405134 707750
rect 408234 655099 408854 709670
rect 411294 655099 411914 705830
rect 411954 655099 412574 711590
rect 415014 655099 415634 707750
rect 418734 655099 419354 709670
rect 421794 655099 422414 705830
rect 422454 655099 423074 711590
rect 425514 655099 426134 707750
rect 429234 655099 429854 709670
rect 432294 655099 432914 705830
rect 432954 655099 433574 711590
rect 436014 655099 436634 707750
rect 439734 655099 440354 709670
rect 442794 655099 443414 705830
rect 379794 568099 380414 588000
rect 380454 568099 381074 588000
rect 383514 568099 384134 588000
rect 387234 568099 387854 588000
rect 390294 568099 390914 588000
rect 390954 568099 391574 588000
rect 394014 568099 394634 588000
rect 397734 568099 398354 588000
rect 400794 568099 401414 588000
rect 401454 568099 402074 588000
rect 404514 568099 405134 588000
rect 408234 568099 408854 588000
rect 411294 568099 411914 588000
rect 411954 568099 412574 588000
rect 415014 568099 415634 588000
rect 418734 568099 419354 588000
rect 421794 568099 422414 588000
rect 422454 568099 423074 588000
rect 425514 568099 426134 588000
rect 429234 568099 429854 588000
rect 432294 568099 432914 588000
rect 432954 568099 433574 588000
rect 436014 568099 436634 588000
rect 439734 568099 440354 588000
rect 442794 568099 443414 588000
rect 379794 -1894 380414 501000
rect 380454 -7654 381074 501000
rect 383514 -3814 384134 501000
rect 387234 -5734 387854 501000
rect 390294 -1894 390914 501000
rect 390954 -7654 391574 501000
rect 394014 -3814 394634 501000
rect 397734 465308 398354 501000
rect 400794 465308 401414 501000
rect 401454 465308 402074 501000
rect 404514 465308 405134 501000
rect 408234 465308 408854 501000
rect 411294 465308 411914 501000
rect 411954 465308 412574 501000
rect 415014 465308 415634 501000
rect 418734 465308 419354 501000
rect 421794 465308 422414 501000
rect 422454 465308 423074 501000
rect 425514 465308 426134 501000
rect 429234 465308 429854 501000
rect 432294 465308 432914 501000
rect 432954 465308 433574 501000
rect 436014 465308 436634 501000
rect 439734 465308 440354 501000
rect 442794 465308 443414 501000
rect 443454 465308 444074 711590
rect 446514 465308 447134 707750
rect 450234 465308 450854 709670
rect 453294 465308 453914 705830
rect 453954 465308 454574 711590
rect 457014 465308 457634 707750
rect 460734 465308 461354 709670
rect 463794 465308 464414 705830
rect 464454 465308 465074 711590
rect 467514 465308 468134 707750
rect 471234 465308 471854 709670
rect 474294 655099 474914 705830
rect 474954 655099 475574 711590
rect 478014 655099 478634 707750
rect 481734 655099 482354 709670
rect 484794 655099 485414 705830
rect 485454 655099 486074 711590
rect 488514 655099 489134 707750
rect 492234 655099 492854 709670
rect 495294 655099 495914 705830
rect 495954 655099 496574 711590
rect 499014 655099 499634 707750
rect 502734 655099 503354 709670
rect 505794 655099 506414 705830
rect 506454 655099 507074 711590
rect 509514 655099 510134 707750
rect 513234 655099 513854 709670
rect 516294 655099 516914 705830
rect 516954 655099 517574 711590
rect 520014 655099 520634 707750
rect 523734 655099 524354 709670
rect 526794 655099 527414 705830
rect 527454 655099 528074 711590
rect 530514 655099 531134 707750
rect 534234 655099 534854 709670
rect 537294 655099 537914 705830
rect 537954 655099 538574 711590
rect 474294 568000 474914 588000
rect 474954 568000 475574 588000
rect 478014 568000 478634 588000
rect 481734 568000 482354 588000
rect 484794 568000 485414 588000
rect 485454 568000 486074 588000
rect 488514 568000 489134 588000
rect 492234 568000 492854 588000
rect 495294 568000 495914 588000
rect 495954 568000 496574 588000
rect 499014 568000 499634 588000
rect 502734 568000 503354 588000
rect 505794 568000 506414 588000
rect 506454 568000 507074 588000
rect 509514 568000 510134 588000
rect 513234 568000 513854 588000
rect 516294 568000 516914 588000
rect 516954 568000 517574 588000
rect 520014 568000 520634 588000
rect 523734 568000 524354 588000
rect 526794 568000 527414 588000
rect 474294 465308 474914 514000
rect 474954 465308 475574 514000
rect 478014 465308 478634 514000
rect 481734 465308 482354 514000
rect 484794 465308 485414 514000
rect 485454 465308 486074 514000
rect 488514 465308 489134 514000
rect 492234 465308 492854 514000
rect 495294 465308 495914 514000
rect 495954 465308 496574 514000
rect 499014 465308 499634 514000
rect 502734 465308 503354 514000
rect 505794 465308 506414 514000
rect 506454 465308 507074 514000
rect 509514 465308 510134 514000
rect 513234 465308 513854 514000
rect 516294 465308 516914 514000
rect 516954 465308 517574 514000
rect 520014 465308 520634 514000
rect 523734 465308 524354 514000
rect 526794 465308 527414 514000
rect 527454 465308 528074 588000
rect 530514 465308 531134 588000
rect 534234 465308 534854 588000
rect 537294 465308 537914 588000
rect 537954 465308 538574 588000
rect 397734 355308 398354 378000
rect 400794 355308 401414 378000
rect 401454 355308 402074 378000
rect 404514 355308 405134 378000
rect 408234 355308 408854 378000
rect 411294 355308 411914 378000
rect 411954 355308 412574 378000
rect 415014 355308 415634 378000
rect 418734 355308 419354 378000
rect 421794 355308 422414 378000
rect 422454 355308 423074 378000
rect 425514 355308 426134 378000
rect 429234 355308 429854 378000
rect 432294 355308 432914 378000
rect 432954 355308 433574 378000
rect 436014 355308 436634 378000
rect 439734 355308 440354 378000
rect 442794 355308 443414 378000
rect 443454 355308 444074 378000
rect 446514 355308 447134 378000
rect 450234 355308 450854 378000
rect 453294 355308 453914 378000
rect 453954 355308 454574 378000
rect 457014 355308 457634 378000
rect 460734 355308 461354 378000
rect 463794 355308 464414 378000
rect 464454 355308 465074 378000
rect 467514 355308 468134 378000
rect 471234 355308 471854 378000
rect 474294 355308 474914 378000
rect 474954 355308 475574 378000
rect 478014 355308 478634 378000
rect 481734 355308 482354 378000
rect 484794 355308 485414 378000
rect 485454 355308 486074 378000
rect 488514 355308 489134 378000
rect 492234 355308 492854 378000
rect 495294 355308 495914 378000
rect 495954 355308 496574 378000
rect 499014 355308 499634 378000
rect 502734 355308 503354 378000
rect 505794 355308 506414 378000
rect 506454 355308 507074 378000
rect 509514 355308 510134 378000
rect 513234 355308 513854 378000
rect 516294 355308 516914 378000
rect 516954 355308 517574 378000
rect 520014 355308 520634 378000
rect 523734 355308 524354 378000
rect 526794 355308 527414 378000
rect 527454 355308 528074 378000
rect 530514 355308 531134 378000
rect 534234 355308 534854 378000
rect 537294 355308 537914 378000
rect 537954 355308 538574 378000
rect 397734 245308 398354 268000
rect 400794 245308 401414 268000
rect 401454 245308 402074 268000
rect 404514 245308 405134 268000
rect 408234 245308 408854 268000
rect 411294 245308 411914 268000
rect 411954 245308 412574 268000
rect 415014 245308 415634 268000
rect 418734 245308 419354 268000
rect 421794 245308 422414 268000
rect 422454 245308 423074 268000
rect 425514 245308 426134 268000
rect 429234 245308 429854 268000
rect 432294 245308 432914 268000
rect 432954 245308 433574 268000
rect 436014 245308 436634 268000
rect 439734 245308 440354 268000
rect 442794 245308 443414 268000
rect 443454 245308 444074 268000
rect 446514 245308 447134 268000
rect 450234 245308 450854 268000
rect 453294 245308 453914 268000
rect 453954 245308 454574 268000
rect 457014 245308 457634 268000
rect 460734 245308 461354 268000
rect 463794 245308 464414 268000
rect 464454 245308 465074 268000
rect 467514 245308 468134 268000
rect 471234 245308 471854 268000
rect 474294 245308 474914 268000
rect 474954 245308 475574 268000
rect 478014 245308 478634 268000
rect 481734 245308 482354 268000
rect 484794 245308 485414 268000
rect 485454 245308 486074 268000
rect 488514 245308 489134 268000
rect 492234 245308 492854 268000
rect 495294 245308 495914 268000
rect 495954 245308 496574 268000
rect 499014 245308 499634 268000
rect 502734 245308 503354 268000
rect 505794 245308 506414 268000
rect 506454 245308 507074 268000
rect 509514 245308 510134 268000
rect 513234 245308 513854 268000
rect 516294 245308 516914 268000
rect 516954 245308 517574 268000
rect 520014 245308 520634 268000
rect 523734 245308 524354 268000
rect 526794 245308 527414 268000
rect 527454 245308 528074 268000
rect 530514 245308 531134 268000
rect 534234 245308 534854 268000
rect 537294 245308 537914 268000
rect 537954 245308 538574 268000
rect 397734 135308 398354 158000
rect 400794 135308 401414 158000
rect 401454 135308 402074 158000
rect 404514 135308 405134 158000
rect 408234 135308 408854 158000
rect 411294 135308 411914 158000
rect 411954 135308 412574 158000
rect 415014 135308 415634 158000
rect 418734 135308 419354 158000
rect 421794 135308 422414 158000
rect 422454 135308 423074 158000
rect 425514 135308 426134 158000
rect 429234 135308 429854 158000
rect 432294 135308 432914 158000
rect 432954 135308 433574 158000
rect 436014 135308 436634 158000
rect 439734 135308 440354 158000
rect 442794 135308 443414 158000
rect 443454 135308 444074 158000
rect 446514 135308 447134 158000
rect 450234 135308 450854 158000
rect 453294 135308 453914 158000
rect 453954 135308 454574 158000
rect 457014 135308 457634 158000
rect 460734 135308 461354 158000
rect 463794 135308 464414 158000
rect 464454 135308 465074 158000
rect 467514 135308 468134 158000
rect 471234 135308 471854 158000
rect 474294 135308 474914 158000
rect 474954 135308 475574 158000
rect 478014 135308 478634 158000
rect 481734 135308 482354 158000
rect 484794 135308 485414 158000
rect 485454 135308 486074 158000
rect 488514 135308 489134 158000
rect 492234 135308 492854 158000
rect 495294 135308 495914 158000
rect 495954 135308 496574 158000
rect 499014 135308 499634 158000
rect 502734 135308 503354 158000
rect 505794 135308 506414 158000
rect 506454 135308 507074 158000
rect 509514 135308 510134 158000
rect 513234 135308 513854 158000
rect 516294 135308 516914 158000
rect 516954 135308 517574 158000
rect 520014 135308 520634 158000
rect 523734 135308 524354 158000
rect 526794 135308 527414 158000
rect 527454 135308 528074 158000
rect 530514 135308 531134 158000
rect 534234 135308 534854 158000
rect 537294 135308 537914 158000
rect 537954 135308 538574 158000
rect 397734 -5734 398354 48000
rect 400794 -1894 401414 48000
rect 401454 -7654 402074 48000
rect 404514 -3814 405134 48000
rect 408234 -5734 408854 48000
rect 411294 -1894 411914 48000
rect 411954 -7654 412574 48000
rect 415014 -3814 415634 48000
rect 418734 -5734 419354 48000
rect 421794 -1894 422414 48000
rect 422454 -7654 423074 48000
rect 425514 -3814 426134 48000
rect 429234 -5734 429854 48000
rect 432294 -1894 432914 48000
rect 432954 -7654 433574 48000
rect 436014 -3814 436634 48000
rect 439734 -5734 440354 48000
rect 442794 -1894 443414 48000
rect 443454 -7654 444074 48000
rect 446514 -3814 447134 48000
rect 450234 -5734 450854 48000
rect 453294 -1894 453914 48000
rect 453954 -7654 454574 48000
rect 457014 -3814 457634 48000
rect 460734 -5734 461354 48000
rect 463794 -1894 464414 48000
rect 464454 -7654 465074 48000
rect 467514 -3814 468134 48000
rect 471234 -5734 471854 48000
rect 474294 -1894 474914 48000
rect 474954 -7654 475574 48000
rect 478014 -3814 478634 48000
rect 481734 -5734 482354 48000
rect 484794 -1894 485414 48000
rect 485454 -7654 486074 48000
rect 488514 -3814 489134 48000
rect 492234 -5734 492854 48000
rect 495294 -1894 495914 48000
rect 495954 -7654 496574 48000
rect 499014 -3814 499634 48000
rect 502734 -5734 503354 48000
rect 505794 -1894 506414 48000
rect 506454 -7654 507074 48000
rect 509514 -3814 510134 48000
rect 513234 -5734 513854 48000
rect 516294 -1894 516914 48000
rect 516954 -7654 517574 48000
rect 520014 -3814 520634 48000
rect 523734 -5734 524354 48000
rect 526794 -1894 527414 48000
rect 527454 -7654 528074 48000
rect 530514 -3814 531134 48000
rect 534234 -5734 534854 48000
rect 537294 -1894 537914 48000
rect 537954 -7654 538574 48000
rect 541014 -3814 541634 707750
rect 544734 -5734 545354 709670
rect 547794 -1894 548414 705830
rect 548454 -7654 549074 711590
rect 551514 -3814 552134 707750
rect 555234 -5734 555854 709670
rect 558294 -1894 558914 705830
rect 558954 -7654 559574 711590
rect 562014 -3814 562634 707750
rect 565734 -5734 566354 709670
rect 568794 -1894 569414 705830
rect 569454 -7654 570074 711590
rect 572514 -3814 573134 707750
rect 576234 -5734 576854 709670
rect 579294 -1894 579914 705830
rect 579954 -7654 580574 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 46059 538080 162934 652493
rect 46059 465228 47434 538080
rect 48214 465228 51154 538080
rect 51934 465228 54214 538080
rect 55654 465228 57934 538080
rect 58714 465228 61654 538080
rect 62434 465228 64714 538080
rect 66154 465228 68434 538080
rect 69214 465228 72154 538080
rect 72934 465228 75214 538080
rect 76654 465228 78934 538080
rect 79714 465228 82654 538080
rect 83434 465228 85714 538080
rect 87154 465228 89434 538080
rect 90214 465228 93154 538080
rect 93934 465228 96214 538080
rect 97654 465228 99934 538080
rect 100714 465228 103654 538080
rect 104434 465228 106714 538080
rect 108154 465228 110434 538080
rect 111214 465228 114154 538080
rect 114934 465228 117214 538080
rect 118654 465228 120934 538080
rect 121714 465228 124654 538080
rect 125434 465228 127714 538080
rect 129154 465228 131434 538080
rect 132214 465228 135154 538080
rect 135934 465228 138214 538080
rect 139654 465228 141934 538080
rect 142714 465228 145654 538080
rect 146434 465228 148714 538080
rect 150154 465228 152434 538080
rect 153214 465228 156154 538080
rect 156934 465228 159214 538080
rect 160654 465228 162934 538080
rect 163714 465228 166654 652493
rect 167434 465228 169714 652493
rect 171154 465228 173434 652493
rect 174214 465228 177154 652493
rect 177934 465228 180214 652493
rect 181654 465228 183934 652493
rect 184714 465228 187654 652493
rect 188434 465228 190714 652493
rect 46059 378080 190714 465228
rect 46059 355228 47434 378080
rect 48214 355228 51154 378080
rect 51934 355228 54214 378080
rect 55654 355228 57934 378080
rect 58714 355228 61654 378080
rect 62434 355228 64714 378080
rect 66154 355228 68434 378080
rect 69214 355228 72154 378080
rect 72934 355228 75214 378080
rect 76654 355228 78934 378080
rect 79714 355228 82654 378080
rect 83434 355228 85714 378080
rect 87154 355228 89434 378080
rect 90214 355228 93154 378080
rect 93934 355228 96214 378080
rect 97654 355228 99934 378080
rect 100714 355228 103654 378080
rect 104434 355228 106714 378080
rect 108154 355228 110434 378080
rect 111214 355228 114154 378080
rect 114934 355228 117214 378080
rect 118654 355228 120934 378080
rect 121714 355228 124654 378080
rect 125434 355228 127714 378080
rect 129154 355228 131434 378080
rect 132214 355228 135154 378080
rect 135934 355228 138214 378080
rect 139654 355228 141934 378080
rect 142714 355228 145654 378080
rect 146434 355228 148714 378080
rect 150154 355228 152434 378080
rect 153214 355228 156154 378080
rect 156934 355228 159214 378080
rect 160654 355228 162934 378080
rect 163714 355228 166654 378080
rect 167434 355228 169714 378080
rect 171154 355228 173434 378080
rect 174214 355228 177154 378080
rect 177934 355228 180214 378080
rect 181654 355228 183934 378080
rect 184714 355228 187654 378080
rect 188434 355228 190714 378080
rect 46059 268080 190714 355228
rect 46059 245228 47434 268080
rect 48214 245228 51154 268080
rect 51934 245228 54214 268080
rect 55654 245228 57934 268080
rect 58714 245228 61654 268080
rect 62434 245228 64714 268080
rect 66154 245228 68434 268080
rect 69214 245228 72154 268080
rect 72934 245228 75214 268080
rect 76654 245228 78934 268080
rect 79714 245228 82654 268080
rect 83434 245228 85714 268080
rect 87154 245228 89434 268080
rect 90214 245228 93154 268080
rect 93934 245228 96214 268080
rect 97654 245228 99934 268080
rect 100714 245228 103654 268080
rect 104434 245228 106714 268080
rect 108154 245228 110434 268080
rect 111214 245228 114154 268080
rect 114934 245228 117214 268080
rect 118654 245228 120934 268080
rect 121714 245228 124654 268080
rect 125434 245228 127714 268080
rect 129154 245228 131434 268080
rect 132214 245228 135154 268080
rect 135934 245228 138214 268080
rect 139654 245228 141934 268080
rect 142714 245228 145654 268080
rect 146434 245228 148714 268080
rect 150154 245228 152434 268080
rect 153214 245228 156154 268080
rect 156934 245228 159214 268080
rect 160654 245228 162934 268080
rect 163714 245228 166654 268080
rect 167434 245228 169714 268080
rect 171154 245228 173434 268080
rect 174214 245228 177154 268080
rect 177934 245228 180214 268080
rect 181654 245228 183934 268080
rect 184714 245228 187654 268080
rect 188434 245228 190714 268080
rect 46059 158080 190714 245228
rect 46059 135228 47434 158080
rect 48214 135228 51154 158080
rect 51934 135228 54214 158080
rect 55654 135228 57934 158080
rect 58714 135228 61654 158080
rect 62434 135228 64714 158080
rect 66154 135228 68434 158080
rect 69214 135228 72154 158080
rect 72934 135228 75214 158080
rect 76654 135228 78934 158080
rect 79714 135228 82654 158080
rect 83434 135228 85714 158080
rect 87154 135228 89434 158080
rect 90214 135228 93154 158080
rect 93934 135228 96214 158080
rect 97654 135228 99934 158080
rect 100714 135228 103654 158080
rect 104434 135228 106714 158080
rect 108154 135228 110434 158080
rect 111214 135228 114154 158080
rect 114934 135228 117214 158080
rect 118654 135228 120934 158080
rect 121714 135228 124654 158080
rect 125434 135228 127714 158080
rect 129154 135228 131434 158080
rect 132214 135228 135154 158080
rect 135934 135228 138214 158080
rect 139654 135228 141934 158080
rect 142714 135228 145654 158080
rect 146434 135228 148714 158080
rect 150154 135228 152434 158080
rect 153214 135228 156154 158080
rect 156934 135228 159214 158080
rect 160654 135228 162934 158080
rect 163714 135228 166654 158080
rect 167434 135228 169714 158080
rect 171154 135228 173434 158080
rect 174214 135228 177154 158080
rect 177934 135228 180214 158080
rect 181654 135228 183934 158080
rect 184714 135228 187654 158080
rect 188434 135228 190714 158080
rect 46059 48080 190714 135228
rect 46059 3299 47434 48080
rect 48214 3299 51154 48080
rect 51934 3299 54214 48080
rect 55654 3299 57934 48080
rect 58714 3299 61654 48080
rect 62434 3299 64714 48080
rect 66154 3299 68434 48080
rect 69214 3299 72154 48080
rect 72934 3299 75214 48080
rect 76654 3299 78934 48080
rect 79714 3299 82654 48080
rect 83434 3299 85714 48080
rect 87154 3299 89434 48080
rect 90214 3299 93154 48080
rect 93934 3299 96214 48080
rect 97654 3299 99934 48080
rect 100714 3299 103654 48080
rect 104434 3299 106714 48080
rect 108154 3299 110434 48080
rect 111214 3299 114154 48080
rect 114934 3299 117214 48080
rect 118654 3299 120934 48080
rect 121714 3299 124654 48080
rect 125434 3299 127714 48080
rect 129154 3299 131434 48080
rect 132214 3299 135154 48080
rect 135934 3299 138214 48080
rect 139654 3299 141934 48080
rect 142714 3299 145654 48080
rect 146434 3299 148714 48080
rect 150154 3299 152434 48080
rect 153214 3299 156154 48080
rect 156934 3299 159214 48080
rect 160654 3299 162934 48080
rect 163714 3299 166654 48080
rect 167434 3299 169714 48080
rect 171154 3299 173434 48080
rect 174214 3299 177154 48080
rect 177934 3299 180214 48080
rect 181654 3299 183934 48080
rect 184714 3299 187654 48080
rect 188434 3299 190714 48080
rect 192154 3299 194434 652493
rect 195214 3299 198154 652493
rect 198934 3299 201214 652493
rect 202654 3299 204934 652493
rect 205714 651920 208654 652493
rect 209434 651920 211714 652493
rect 213154 651920 215434 652493
rect 216214 651920 219154 652493
rect 219934 651920 222214 652493
rect 223654 651920 225934 652493
rect 226714 651920 229654 652493
rect 230434 651920 232714 652493
rect 234154 651920 236434 652493
rect 237214 651920 240154 652493
rect 240934 651920 243214 652493
rect 244654 651920 246934 652493
rect 247714 651920 250654 652493
rect 251434 651920 253714 652493
rect 255154 651920 257434 652493
rect 258214 651920 261154 652493
rect 261934 651920 264214 652493
rect 265654 651920 267934 652493
rect 268714 651920 271654 652493
rect 272434 651920 274714 652493
rect 276154 651920 278434 652493
rect 279214 651920 282154 652493
rect 282934 651920 285214 652493
rect 286654 651920 288934 652493
rect 289714 651920 292654 652493
rect 293434 651920 295714 652493
rect 297154 651920 299434 652493
rect 300214 651920 303154 652493
rect 303934 651920 306214 652493
rect 307654 651920 309934 652493
rect 310714 651920 313654 652493
rect 314434 651920 316714 652493
rect 318154 651920 320434 652493
rect 321214 651920 324154 652493
rect 324934 651920 327214 652493
rect 328654 651920 330934 652493
rect 331714 651920 334654 652493
rect 205714 501080 334654 651920
rect 205714 3299 208654 501080
rect 209434 3299 211714 501080
rect 213154 3299 215434 501080
rect 216214 3299 219154 501080
rect 219934 3299 222214 501080
rect 223654 465228 225934 501080
rect 226714 465228 229654 501080
rect 230434 465228 232714 501080
rect 234154 465228 236434 501080
rect 237214 465228 240154 501080
rect 240934 465228 243214 501080
rect 244654 465228 246934 501080
rect 247714 465228 250654 501080
rect 251434 465228 253714 501080
rect 255154 465228 257434 501080
rect 258214 465228 261154 501080
rect 261934 465228 264214 501080
rect 265654 465228 267934 501080
rect 268714 465228 271654 501080
rect 272434 465228 274714 501080
rect 276154 465228 278434 501080
rect 279214 465228 282154 501080
rect 282934 465228 285214 501080
rect 286654 465228 288934 501080
rect 289714 465228 292654 501080
rect 293434 465228 295714 501080
rect 297154 465228 299434 501080
rect 300214 465228 303154 501080
rect 303934 465228 306214 501080
rect 307654 465228 309934 501080
rect 310714 465228 313654 501080
rect 314434 465228 316714 501080
rect 318154 465228 320434 501080
rect 321214 465228 324154 501080
rect 324934 465228 327214 501080
rect 328654 465228 330934 501080
rect 331714 465228 334654 501080
rect 335434 465228 337714 652493
rect 339154 465228 341434 652493
rect 342214 465228 345154 652493
rect 345934 465228 348214 652493
rect 349654 465228 351934 652493
rect 352714 465228 355654 652493
rect 356434 465228 358714 652493
rect 360154 465228 362434 652493
rect 363214 465228 366154 652493
rect 222994 378080 366154 465228
rect 223654 355228 225934 378080
rect 226714 355228 229654 378080
rect 230434 355228 232714 378080
rect 234154 355228 236434 378080
rect 237214 355228 240154 378080
rect 240934 355228 243214 378080
rect 244654 355228 246934 378080
rect 247714 355228 250654 378080
rect 251434 355228 253714 378080
rect 255154 355228 257434 378080
rect 258214 355228 261154 378080
rect 261934 355228 264214 378080
rect 265654 355228 267934 378080
rect 268714 355228 271654 378080
rect 272434 355228 274714 378080
rect 276154 355228 278434 378080
rect 279214 355228 282154 378080
rect 282934 355228 285214 378080
rect 286654 355228 288934 378080
rect 289714 355228 292654 378080
rect 293434 355228 295714 378080
rect 297154 355228 299434 378080
rect 300214 355228 303154 378080
rect 303934 355228 306214 378080
rect 307654 355228 309934 378080
rect 310714 355228 313654 378080
rect 314434 355228 316714 378080
rect 318154 355228 320434 378080
rect 321214 355228 324154 378080
rect 324934 355228 327214 378080
rect 328654 355228 330934 378080
rect 331714 355228 334654 378080
rect 335434 355228 337714 378080
rect 339154 355228 341434 378080
rect 342214 355228 345154 378080
rect 345934 355228 348214 378080
rect 349654 355228 351934 378080
rect 352714 355228 355654 378080
rect 356434 355228 358714 378080
rect 360154 355228 362434 378080
rect 363214 355228 366154 378080
rect 222994 268080 366154 355228
rect 223654 245228 225934 268080
rect 226714 245228 229654 268080
rect 230434 245228 232714 268080
rect 234154 245228 236434 268080
rect 237214 245228 240154 268080
rect 240934 245228 243214 268080
rect 244654 245228 246934 268080
rect 247714 245228 250654 268080
rect 251434 245228 253714 268080
rect 255154 245228 257434 268080
rect 258214 245228 261154 268080
rect 261934 245228 264214 268080
rect 265654 245228 267934 268080
rect 268714 245228 271654 268080
rect 272434 245228 274714 268080
rect 276154 245228 278434 268080
rect 279214 245228 282154 268080
rect 282934 245228 285214 268080
rect 286654 245228 288934 268080
rect 289714 245228 292654 268080
rect 293434 245228 295714 268080
rect 297154 245228 299434 268080
rect 300214 245228 303154 268080
rect 303934 245228 306214 268080
rect 307654 245228 309934 268080
rect 310714 245228 313654 268080
rect 314434 245228 316714 268080
rect 318154 245228 320434 268080
rect 321214 245228 324154 268080
rect 324934 245228 327214 268080
rect 328654 245228 330934 268080
rect 331714 245228 334654 268080
rect 335434 245228 337714 268080
rect 339154 245228 341434 268080
rect 342214 245228 345154 268080
rect 345934 245228 348214 268080
rect 349654 245228 351934 268080
rect 352714 245228 355654 268080
rect 356434 245228 358714 268080
rect 360154 245228 362434 268080
rect 363214 245228 366154 268080
rect 222994 158080 366154 245228
rect 223654 135228 225934 158080
rect 226714 135228 229654 158080
rect 230434 135228 232714 158080
rect 234154 135228 236434 158080
rect 237214 135228 240154 158080
rect 240934 135228 243214 158080
rect 244654 135228 246934 158080
rect 247714 135228 250654 158080
rect 251434 135228 253714 158080
rect 255154 135228 257434 158080
rect 258214 135228 261154 158080
rect 261934 135228 264214 158080
rect 265654 135228 267934 158080
rect 268714 135228 271654 158080
rect 272434 135228 274714 158080
rect 276154 135228 278434 158080
rect 279214 135228 282154 158080
rect 282934 135228 285214 158080
rect 286654 135228 288934 158080
rect 289714 135228 292654 158080
rect 293434 135228 295714 158080
rect 297154 135228 299434 158080
rect 300214 135228 303154 158080
rect 303934 135228 306214 158080
rect 307654 135228 309934 158080
rect 310714 135228 313654 158080
rect 314434 135228 316714 158080
rect 318154 135228 320434 158080
rect 321214 135228 324154 158080
rect 324934 135228 327214 158080
rect 328654 135228 330934 158080
rect 331714 135228 334654 158080
rect 335434 135228 337714 158080
rect 339154 135228 341434 158080
rect 342214 135228 345154 158080
rect 345934 135228 348214 158080
rect 349654 135228 351934 158080
rect 352714 135228 355654 158080
rect 356434 135228 358714 158080
rect 360154 135228 362434 158080
rect 363214 135228 366154 158080
rect 222994 48080 366154 135228
rect 223654 3299 225934 48080
rect 226714 3299 229654 48080
rect 230434 3299 232714 48080
rect 234154 3299 236434 48080
rect 237214 3299 240154 48080
rect 240934 3299 243214 48080
rect 244654 3299 246934 48080
rect 247714 3299 250654 48080
rect 251434 3299 253714 48080
rect 255154 3299 257434 48080
rect 258214 3299 261154 48080
rect 261934 3299 264214 48080
rect 265654 3299 267934 48080
rect 268714 3299 271654 48080
rect 272434 3299 274714 48080
rect 276154 3299 278434 48080
rect 279214 3299 282154 48080
rect 282934 3299 285214 48080
rect 286654 3299 288934 48080
rect 289714 3299 292654 48080
rect 293434 3299 295714 48080
rect 297154 3299 299434 48080
rect 300214 3299 303154 48080
rect 303934 3299 306214 48080
rect 307654 3299 309934 48080
rect 310714 3299 313654 48080
rect 314434 3299 316714 48080
rect 318154 3299 320434 48080
rect 321214 3299 324154 48080
rect 324934 3299 327214 48080
rect 328654 3299 330934 48080
rect 331714 3299 334654 48080
rect 335434 3299 337714 48080
rect 339154 3299 341434 48080
rect 342214 3299 345154 48080
rect 345934 3299 348214 48080
rect 349654 3299 351934 48080
rect 352714 3299 355654 48080
rect 356434 3299 358714 48080
rect 360154 3299 362434 48080
rect 363214 3299 366154 48080
rect 366934 3299 369214 652493
rect 370654 3299 372934 652493
rect 373714 3299 376654 652493
rect 377434 588080 443374 652493
rect 377434 568019 379714 588080
rect 381154 568019 383434 588080
rect 384214 568019 387154 588080
rect 387934 568019 390214 588080
rect 391654 568019 393934 588080
rect 394714 568019 397654 588080
rect 398434 568019 400714 588080
rect 402154 568019 404434 588080
rect 405214 568019 408154 588080
rect 408934 568019 411214 588080
rect 412654 568019 414934 588080
rect 415714 568019 418654 588080
rect 419434 568019 421714 588080
rect 423154 568019 425434 588080
rect 426214 568019 429154 588080
rect 429934 568019 432214 588080
rect 433654 568019 435934 588080
rect 436714 568019 439654 588080
rect 440434 568019 442714 588080
rect 377434 501080 443374 568019
rect 377434 3299 379714 501080
rect 381154 3299 383434 501080
rect 384214 3299 387154 501080
rect 387934 3299 390214 501080
rect 391654 3299 393934 501080
rect 394714 465228 397654 501080
rect 398434 465228 400714 501080
rect 402154 465228 404434 501080
rect 405214 465228 408154 501080
rect 408934 465228 411214 501080
rect 412654 465228 414934 501080
rect 415714 465228 418654 501080
rect 419434 465228 421714 501080
rect 423154 465228 425434 501080
rect 426214 465228 429154 501080
rect 429934 465228 432214 501080
rect 433654 465228 435934 501080
rect 436714 465228 439654 501080
rect 440434 465228 442714 501080
rect 444154 465228 446434 652493
rect 447214 465228 450154 652493
rect 450934 465228 453214 652493
rect 454654 465228 456934 652493
rect 457714 465228 460654 652493
rect 461434 465228 463714 652493
rect 465154 465228 467434 652493
rect 468214 465228 471154 652493
rect 471934 588080 539061 652493
rect 471934 567920 474214 588080
rect 475654 567920 477934 588080
rect 478714 567920 481654 588080
rect 482434 567920 484714 588080
rect 486154 567920 488434 588080
rect 489214 567920 492154 588080
rect 492934 567920 495214 588080
rect 496654 567920 498934 588080
rect 499714 567920 502654 588080
rect 503434 567920 505714 588080
rect 507154 567920 509434 588080
rect 510214 567920 513154 588080
rect 513934 567920 516214 588080
rect 517654 567920 519934 588080
rect 520714 567920 523654 588080
rect 524434 567920 526714 588080
rect 471934 514080 527374 567920
rect 471934 465228 474214 514080
rect 475654 465228 477934 514080
rect 478714 465228 481654 514080
rect 482434 465228 484714 514080
rect 486154 465228 488434 514080
rect 489214 465228 492154 514080
rect 492934 465228 495214 514080
rect 496654 465228 498934 514080
rect 499714 465228 502654 514080
rect 503434 465228 505714 514080
rect 507154 465228 509434 514080
rect 510214 465228 513154 514080
rect 513934 465228 516214 514080
rect 517654 465228 519934 514080
rect 520714 465228 523654 514080
rect 524434 465228 526714 514080
rect 528154 465228 530434 588080
rect 531214 465228 534154 588080
rect 534934 465228 537214 588080
rect 538654 465228 539061 588080
rect 394714 378080 539061 465228
rect 394714 355228 397654 378080
rect 398434 355228 400714 378080
rect 402154 355228 404434 378080
rect 405214 355228 408154 378080
rect 408934 355228 411214 378080
rect 412654 355228 414934 378080
rect 415714 355228 418654 378080
rect 419434 355228 421714 378080
rect 423154 355228 425434 378080
rect 426214 355228 429154 378080
rect 429934 355228 432214 378080
rect 433654 355228 435934 378080
rect 436714 355228 439654 378080
rect 440434 355228 442714 378080
rect 444154 355228 446434 378080
rect 447214 355228 450154 378080
rect 450934 355228 453214 378080
rect 454654 355228 456934 378080
rect 457714 355228 460654 378080
rect 461434 355228 463714 378080
rect 465154 355228 467434 378080
rect 468214 355228 471154 378080
rect 471934 355228 474214 378080
rect 475654 355228 477934 378080
rect 478714 355228 481654 378080
rect 482434 355228 484714 378080
rect 486154 355228 488434 378080
rect 489214 355228 492154 378080
rect 492934 355228 495214 378080
rect 496654 355228 498934 378080
rect 499714 355228 502654 378080
rect 503434 355228 505714 378080
rect 507154 355228 509434 378080
rect 510214 355228 513154 378080
rect 513934 355228 516214 378080
rect 517654 355228 519934 378080
rect 520714 355228 523654 378080
rect 524434 355228 526714 378080
rect 528154 355228 530434 378080
rect 531214 355228 534154 378080
rect 534934 355228 537214 378080
rect 538654 355228 539061 378080
rect 394714 268080 539061 355228
rect 394714 245228 397654 268080
rect 398434 245228 400714 268080
rect 402154 245228 404434 268080
rect 405214 245228 408154 268080
rect 408934 245228 411214 268080
rect 412654 245228 414934 268080
rect 415714 245228 418654 268080
rect 419434 245228 421714 268080
rect 423154 245228 425434 268080
rect 426214 245228 429154 268080
rect 429934 245228 432214 268080
rect 433654 245228 435934 268080
rect 436714 245228 439654 268080
rect 440434 245228 442714 268080
rect 444154 245228 446434 268080
rect 447214 245228 450154 268080
rect 450934 245228 453214 268080
rect 454654 245228 456934 268080
rect 457714 245228 460654 268080
rect 461434 245228 463714 268080
rect 465154 245228 467434 268080
rect 468214 245228 471154 268080
rect 471934 245228 474214 268080
rect 475654 245228 477934 268080
rect 478714 245228 481654 268080
rect 482434 245228 484714 268080
rect 486154 245228 488434 268080
rect 489214 245228 492154 268080
rect 492934 245228 495214 268080
rect 496654 245228 498934 268080
rect 499714 245228 502654 268080
rect 503434 245228 505714 268080
rect 507154 245228 509434 268080
rect 510214 245228 513154 268080
rect 513934 245228 516214 268080
rect 517654 245228 519934 268080
rect 520714 245228 523654 268080
rect 524434 245228 526714 268080
rect 528154 245228 530434 268080
rect 531214 245228 534154 268080
rect 534934 245228 537214 268080
rect 538654 245228 539061 268080
rect 394714 158080 539061 245228
rect 394714 135228 397654 158080
rect 398434 135228 400714 158080
rect 402154 135228 404434 158080
rect 405214 135228 408154 158080
rect 408934 135228 411214 158080
rect 412654 135228 414934 158080
rect 415714 135228 418654 158080
rect 419434 135228 421714 158080
rect 423154 135228 425434 158080
rect 426214 135228 429154 158080
rect 429934 135228 432214 158080
rect 433654 135228 435934 158080
rect 436714 135228 439654 158080
rect 440434 135228 442714 158080
rect 444154 135228 446434 158080
rect 447214 135228 450154 158080
rect 450934 135228 453214 158080
rect 454654 135228 456934 158080
rect 457714 135228 460654 158080
rect 461434 135228 463714 158080
rect 465154 135228 467434 158080
rect 468214 135228 471154 158080
rect 471934 135228 474214 158080
rect 475654 135228 477934 158080
rect 478714 135228 481654 158080
rect 482434 135228 484714 158080
rect 486154 135228 488434 158080
rect 489214 135228 492154 158080
rect 492934 135228 495214 158080
rect 496654 135228 498934 158080
rect 499714 135228 502654 158080
rect 503434 135228 505714 158080
rect 507154 135228 509434 158080
rect 510214 135228 513154 158080
rect 513934 135228 516214 158080
rect 517654 135228 519934 158080
rect 520714 135228 523654 158080
rect 524434 135228 526714 158080
rect 528154 135228 530434 158080
rect 531214 135228 534154 158080
rect 534934 135228 537214 158080
rect 538654 135228 539061 158080
rect 394714 48080 539061 135228
rect 394714 3299 397654 48080
rect 398434 3299 400714 48080
rect 402154 3299 404434 48080
rect 405214 3299 408154 48080
rect 408934 3299 411214 48080
rect 412654 3299 414934 48080
rect 415714 3299 418654 48080
rect 419434 3299 421714 48080
rect 423154 3299 425434 48080
rect 426214 3299 429154 48080
rect 429934 3299 432214 48080
rect 433654 3299 435934 48080
rect 436714 3299 439654 48080
rect 440434 3299 442714 48080
rect 444154 3299 446434 48080
rect 447214 3299 450154 48080
rect 450934 3299 453214 48080
rect 454654 3299 456934 48080
rect 457714 3299 460654 48080
rect 461434 3299 463714 48080
rect 465154 3299 467434 48080
rect 468214 3299 471154 48080
rect 471934 3299 474214 48080
rect 475654 3299 477934 48080
rect 478714 3299 481654 48080
rect 482434 3299 484714 48080
rect 486154 3299 488434 48080
rect 489214 3299 492154 48080
rect 492934 3299 495214 48080
rect 496654 3299 498934 48080
rect 499714 3299 502654 48080
rect 503434 3299 505714 48080
rect 507154 3299 509434 48080
rect 510214 3299 513154 48080
rect 513934 3299 516214 48080
rect 517654 3299 519934 48080
rect 520714 3299 523654 48080
rect 524434 3299 526714 48080
rect 528154 3299 530434 48080
rect 531214 3299 534154 48080
rect 534934 3299 537214 48080
rect 538654 3299 539061 48080
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -4886 699586 588810 700206
rect -8726 696526 592650 697146
rect -2966 695866 586890 696486
rect -6806 692806 590730 693426
rect -4886 689086 588810 689706
rect -8726 686026 592650 686646
rect -2966 685366 586890 685986
rect -6806 682306 590730 682926
rect -4886 678586 588810 679206
rect -8726 675526 592650 676146
rect -2966 674866 586890 675486
rect -6806 671806 590730 672426
rect -4886 668086 588810 668706
rect -8726 665026 592650 665646
rect -2966 664366 586890 664986
rect -6806 661306 590730 661926
rect -4886 657586 588810 658206
rect -8726 654526 592650 655146
rect -2966 653866 586890 654486
rect -6806 650806 590730 651426
rect -4886 647086 588810 647706
rect -8726 644026 592650 644646
rect -2966 643366 586890 643986
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -8726 633526 592650 634146
rect -2966 632866 586890 633486
rect -6806 629806 590730 630426
rect -4886 626086 588810 626706
rect -8726 623026 592650 623646
rect -2966 622366 586890 622986
rect -6806 619306 590730 619926
rect -4886 615586 588810 616206
rect -8726 612526 592650 613146
rect -2966 611866 586890 612486
rect -6806 608806 590730 609426
rect -4886 605086 588810 605706
rect -8726 602026 592650 602646
rect -2966 601366 586890 601986
rect -6806 598306 590730 598926
rect -4886 594586 588810 595206
rect -8726 591526 592650 592146
rect -2966 590866 586890 591486
rect -6806 587806 590730 588426
rect -4886 584086 588810 584706
rect -8726 581026 592650 581646
rect -2966 580366 586890 580986
rect 397734 578246 440354 578866
rect 481734 578246 524354 578866
rect -6806 577306 590730 577926
rect -4886 573586 588810 574206
rect -8726 570526 592650 571146
rect -2966 569866 586890 570486
rect -6806 566806 590730 567426
rect -4886 563086 588810 563706
rect -8726 560026 592650 560646
rect -2966 559366 586890 559986
rect -6806 556306 590730 556926
rect -4886 552586 588810 553206
rect -8726 549526 592650 550146
rect -2966 548866 586890 549486
rect -6806 545806 590730 546426
rect -4886 542086 588810 542706
rect -8726 539026 592650 539646
rect -2966 538366 586890 538986
rect -6806 535306 590730 535926
rect -4886 531586 588810 532206
rect -8726 528526 592650 529146
rect -2966 527866 586890 528486
rect -6806 524806 590730 525426
rect -4886 521086 588810 521706
rect -8726 518026 592650 518646
rect -2966 517366 586890 517986
rect -6806 514306 590730 514926
rect -4886 510586 588810 511206
rect -8726 507526 592650 508146
rect -2966 506866 586890 507486
rect -6806 503806 590730 504426
rect -4886 500086 588810 500706
rect -8726 497026 592650 497646
rect -2966 496366 586890 496986
rect -6806 493306 590730 493926
rect -4886 489586 588810 490206
rect -8726 486526 592650 487146
rect -2966 485866 586890 486486
rect -6806 482806 590730 483426
rect -4886 479086 588810 479706
rect -8726 476026 592650 476646
rect -2966 475366 586890 475986
rect -6806 472306 590730 472926
rect -4886 468586 588810 469206
rect -8726 465526 592650 466146
rect -2966 464866 586890 465486
rect -6806 461806 590730 462426
rect -4886 458086 588810 458706
rect -8726 455026 592650 455646
rect -2966 454366 586890 454986
rect -6806 451306 590730 451926
rect -4886 447586 588810 448206
rect -8726 444526 592650 445146
rect -2966 443866 586890 444486
rect -6806 440806 590730 441426
rect -4886 437086 588810 437706
rect -8726 434026 592650 434646
rect -2966 433366 586890 433986
rect -6806 430306 590730 430926
rect -4886 426586 588810 427206
rect -8726 423526 592650 424146
rect -2966 422866 586890 423486
rect -6806 419806 590730 420426
rect -4886 416086 588810 416706
rect -8726 413026 592650 413646
rect -2966 412366 586890 412986
rect -6806 409306 590730 409926
rect -4886 405586 588810 406206
rect -8726 402526 592650 403146
rect -2966 401866 586890 402486
rect -6806 398806 590730 399426
rect -4886 395086 588810 395706
rect -8726 392026 592650 392646
rect -2966 391366 586890 391986
rect -6806 388306 590730 388926
rect -4886 384586 588810 385206
rect -8726 381526 592650 382146
rect -2966 380866 586890 381486
rect -6806 377806 590730 378426
rect -4886 374086 588810 374706
rect -8726 371026 592650 371646
rect -2966 370366 586890 370986
rect -6806 367306 590730 367926
rect -4886 363586 588810 364206
rect -8726 360526 592650 361146
rect -2966 359866 586890 360486
rect -6806 356806 590730 357426
rect -4886 353086 588810 353706
rect -8726 350026 592650 350646
rect -2966 349366 586890 349986
rect -6806 346306 590730 346926
rect -4886 342586 588810 343206
rect -8726 339526 592650 340146
rect -2966 338866 586890 339486
rect -6806 335806 590730 336426
rect -4886 332086 588810 332706
rect -8726 329026 592650 329646
rect -2966 328366 586890 328986
rect -6806 325306 590730 325926
rect -4886 321586 588810 322206
rect -8726 318526 592650 319146
rect -2966 317866 586890 318486
rect -6806 314806 590730 315426
rect -4886 311086 588810 311706
rect -8726 308026 592650 308646
rect -2966 307366 586890 307986
rect -6806 304306 590730 304926
rect -4886 300586 588810 301206
rect -8726 297526 592650 298146
rect -2966 296866 586890 297486
rect -6806 293806 590730 294426
rect -4886 290086 588810 290706
rect -8726 287026 592650 287646
rect -2966 286366 586890 286986
rect -6806 283306 590730 283926
rect -4886 279586 588810 280206
rect -8726 276526 592650 277146
rect -2966 275866 586890 276486
rect -6806 272806 590730 273426
rect -4886 269086 588810 269706
rect -8726 266026 592650 266646
rect -2966 265366 586890 265986
rect -6806 262306 590730 262926
rect -4886 258586 588810 259206
rect -8726 255526 592650 256146
rect -2966 254866 586890 255486
rect -6806 251806 590730 252426
rect -4886 248086 588810 248706
rect -8726 245026 592650 245646
rect -2966 244366 586890 244986
rect -6806 241306 590730 241926
rect -4886 237586 588810 238206
rect -8726 234526 592650 235146
rect -2966 233866 586890 234486
rect -6806 230806 590730 231426
rect -4886 227086 588810 227706
rect -8726 224026 592650 224646
rect -2966 223366 586890 223986
rect -6806 220306 590730 220926
rect -4886 216586 588810 217206
rect -8726 213526 592650 214146
rect -2966 212866 586890 213486
rect -6806 209806 590730 210426
rect -4886 206086 588810 206706
rect -8726 203026 592650 203646
rect -2966 202366 586890 202986
rect -6806 199306 590730 199926
rect -4886 195586 588810 196206
rect -8726 192526 592650 193146
rect -2966 191866 586890 192486
rect -6806 188806 590730 189426
rect -4886 185086 588810 185706
rect -8726 182026 592650 182646
rect -2966 181366 586890 181986
rect -6806 178306 590730 178926
rect -4886 174586 588810 175206
rect -8726 171526 592650 172146
rect -2966 170866 586890 171486
rect -6806 167806 590730 168426
rect -4886 164086 588810 164706
rect -8726 161026 592650 161646
rect -2966 160366 586890 160986
rect -6806 157306 590730 157926
rect -4886 153586 588810 154206
rect -8726 150526 592650 151146
rect -2966 149866 586890 150486
rect -6806 146806 590730 147426
rect -4886 143086 588810 143706
rect -8726 140026 592650 140646
rect -2966 139366 586890 139986
rect -6806 136306 590730 136926
rect -4886 132586 588810 133206
rect -8726 129526 592650 130146
rect -2966 128866 586890 129486
rect -6806 125806 590730 126426
rect -4886 122086 588810 122706
rect -8726 119026 592650 119646
rect -2966 118366 586890 118986
rect -6806 115306 590730 115926
rect -4886 111586 588810 112206
rect -8726 108526 592650 109146
rect -2966 107866 586890 108486
rect -6806 104806 590730 105426
rect -4886 101086 588810 101706
rect -8726 98026 592650 98646
rect -2966 97366 586890 97986
rect -6806 94306 590730 94926
rect -4886 90586 588810 91206
rect -8726 87526 592650 88146
rect -2966 86866 586890 87486
rect -6806 83806 590730 84426
rect -4886 80086 588810 80706
rect -8726 77026 592650 77646
rect -2966 76366 586890 76986
rect -6806 73306 590730 73926
rect -4886 69586 588810 70206
rect -8726 66526 592650 67146
rect -2966 65866 586890 66486
rect -6806 62806 590730 63426
rect -4886 59086 588810 59706
rect -8726 56026 592650 56646
rect -2966 55366 586890 55986
rect -6806 52306 590730 52926
rect -4886 48586 588810 49206
rect -8726 45526 592650 46146
rect -2966 44866 586890 45486
rect -6806 41806 590730 42426
rect -4886 38086 588810 38706
rect -8726 35026 592650 35646
rect -2966 34366 586890 34986
rect -6806 31306 590730 31926
rect -4886 27586 588810 28206
rect -8726 24526 592650 25146
rect -2966 23866 586890 24486
rect -6806 20806 590730 21426
rect -4886 17086 588810 17706
rect -8726 14026 592650 14646
rect -2966 13366 586890 13986
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 23866 586890 24486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 44866 586890 45486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 65866 586890 66486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 86866 586890 87486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 107866 586890 108486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 128866 586890 129486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 149866 586890 150486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 170866 586890 171486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 191866 586890 192486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 212866 586890 213486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 233866 586890 234486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 275866 586890 276486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 296866 586890 297486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 317866 586890 318486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 338866 586890 339486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 359866 586890 360486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 380866 586890 381486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 401866 586890 402486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 422866 586890 423486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 443866 586890 444486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 464866 586890 465486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 485866 586890 486486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 527866 586890 528486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 548866 586890 549486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 569866 586890 570486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 590866 586890 591486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 611866 586890 612486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 632866 586890 633486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 653866 586890 654486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 674866 586890 675486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 695866 586890 696486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 64794 -1894 65414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 -1894 86414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 106794 -1894 107414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 -1894 128414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 148794 -1894 149414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 -1894 170414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 232794 -1894 233414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 -1894 254414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 274794 -1894 275414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 295794 -1894 296414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 316794 -1894 317414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 -1894 338414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 358794 -1894 359414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 400794 -1894 401414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 -1894 422414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 442794 -1894 443414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 463794 -1894 464414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 484794 -1894 485414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 -1894 506414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 526794 -1894 527414 48000 6 vccd1
port 532 nsew power input
rlabel metal4 s 64794 135308 65414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 135308 86414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 106794 135308 107414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 135308 128414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 148794 135308 149414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 135308 170414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 232794 135308 233414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 135308 254414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 274794 135308 275414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 295794 135308 296414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 316794 135308 317414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 135308 338414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 358794 135308 359414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 400794 135308 401414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 135308 422414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 442794 135308 443414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 463794 135308 464414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 484794 135308 485414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 135308 506414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 526794 135308 527414 158000 6 vccd1
port 532 nsew power input
rlabel metal4 s 64794 245308 65414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 245308 86414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 106794 245308 107414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 245308 128414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 148794 245308 149414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 245308 170414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 232794 245308 233414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 245308 254414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 274794 245308 275414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 295794 245308 296414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 316794 245308 317414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 245308 338414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 358794 245308 359414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 400794 245308 401414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 245308 422414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 442794 245308 443414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 463794 245308 464414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 484794 245308 485414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 245308 506414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 526794 245308 527414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 64794 355308 65414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 355308 86414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 106794 355308 107414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 355308 128414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 148794 355308 149414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 355308 170414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 232794 355308 233414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 355308 254414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 274794 355308 275414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 295794 355308 296414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 316794 355308 317414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 355308 338414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 358794 355308 359414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 400794 355308 401414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 355308 422414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 442794 355308 443414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 463794 355308 464414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 484794 355308 485414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 355308 506414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 526794 355308 527414 378000 6 vccd1
port 532 nsew power input
rlabel metal4 s 211794 -1894 212414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 232794 465308 233414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 465308 254414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 274794 465308 275414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 295794 465308 296414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 316794 465308 317414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 -1894 380414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 400794 465308 401414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 465308 422414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 442794 465308 443414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 484794 465308 485414 514000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 465308 506414 514000 6 vccd1
port 532 nsew power input
rlabel metal4 s 526794 465308 527414 514000 6 vccd1
port 532 nsew power input
rlabel metal4 s 64794 465308 65414 538000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 465308 86414 538000 6 vccd1
port 532 nsew power input
rlabel metal4 s 106794 465308 107414 538000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 465308 128414 538000 6 vccd1
port 532 nsew power input
rlabel metal4 s 148794 465308 149414 538000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 568099 380414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 400794 568099 401414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 568099 422414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 442794 568099 443414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 484794 568000 485414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 568000 506414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 526794 568000 527414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 22794 -1894 23414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 43794 -1894 44414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 64794 653033 65414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 653033 86414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 106794 653033 107414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 653033 128414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 148794 653033 149414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 465308 170414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 190794 -1894 191414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 211794 652000 212414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 232794 652000 233414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 652000 254414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 274794 652000 275414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 295794 652000 296414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 316794 652000 317414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 465308 338414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 358794 465308 359414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 655099 380414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 400794 655099 401414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 655099 422414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 442794 655099 443414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 463794 465308 464414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 484794 655099 485414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 655099 506414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 526794 655099 527414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 547794 -1894 548414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 568794 -1894 569414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 27586 588810 28206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 48586 588810 49206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 69586 588810 70206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 90586 588810 91206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 111586 588810 112206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 132586 588810 133206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 153586 588810 154206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 174586 588810 175206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 195586 588810 196206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 216586 588810 217206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 237586 588810 238206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 279586 588810 280206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 300586 588810 301206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 321586 588810 322206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 342586 588810 343206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 363586 588810 364206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 384586 588810 385206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 405586 588810 406206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 426586 588810 427206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 447586 588810 448206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 468586 588810 469206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 489586 588810 490206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 531586 588810 532206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 552586 588810 553206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 573586 588810 574206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 594586 588810 595206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 615586 588810 616206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 636586 588810 637206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 657586 588810 658206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 678586 588810 679206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 699586 588810 700206 6 vccd2
port 533 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 47514 -3814 48134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 68514 -3814 69134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 -3814 90134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 110514 -3814 111134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 131514 -3814 132134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 152514 -3814 153134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 -3814 174134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 236514 -3814 237134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 -3814 258134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 278514 -3814 279134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 299514 -3814 300134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 320514 -3814 321134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 -3814 342134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 362514 -3814 363134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 404514 -3814 405134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 -3814 426134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 446514 -3814 447134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 467514 -3814 468134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 488514 -3814 489134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 -3814 510134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 530514 -3814 531134 48000 6 vccd2
port 533 nsew power input
rlabel metal4 s 47514 135308 48134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 68514 135308 69134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 135308 90134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 110514 135308 111134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 131514 135308 132134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 152514 135308 153134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 135308 174134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 236514 135308 237134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 135308 258134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 278514 135308 279134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 299514 135308 300134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 320514 135308 321134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 135308 342134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 362514 135308 363134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 404514 135308 405134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 135308 426134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 446514 135308 447134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 467514 135308 468134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 488514 135308 489134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 135308 510134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 530514 135308 531134 158000 6 vccd2
port 533 nsew power input
rlabel metal4 s 47514 245308 48134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 68514 245308 69134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 245308 90134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 110514 245308 111134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 131514 245308 132134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 152514 245308 153134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 245308 174134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 236514 245308 237134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 245308 258134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 278514 245308 279134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 299514 245308 300134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 320514 245308 321134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 245308 342134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 362514 245308 363134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 404514 245308 405134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 245308 426134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 446514 245308 447134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 467514 245308 468134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 488514 245308 489134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 245308 510134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 530514 245308 531134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 47514 355308 48134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 68514 355308 69134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 355308 90134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 110514 355308 111134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 131514 355308 132134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 152514 355308 153134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 355308 174134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 236514 355308 237134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 355308 258134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 278514 355308 279134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 299514 355308 300134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 320514 355308 321134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 355308 342134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 362514 355308 363134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 404514 355308 405134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 355308 426134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 446514 355308 447134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 467514 355308 468134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 488514 355308 489134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 355308 510134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 530514 355308 531134 378000 6 vccd2
port 533 nsew power input
rlabel metal4 s 215514 -3814 216134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 236514 465308 237134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 465308 258134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 278514 465308 279134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 299514 465308 300134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 320514 465308 321134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 383514 -3814 384134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 404514 465308 405134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 465308 426134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 488514 465308 489134 514000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 465308 510134 514000 6 vccd2
port 533 nsew power input
rlabel metal4 s 47514 465308 48134 538000 6 vccd2
port 533 nsew power input
rlabel metal4 s 68514 465308 69134 538000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 465308 90134 538000 6 vccd2
port 533 nsew power input
rlabel metal4 s 110514 465308 111134 538000 6 vccd2
port 533 nsew power input
rlabel metal4 s 131514 465308 132134 538000 6 vccd2
port 533 nsew power input
rlabel metal4 s 152514 465308 153134 538000 6 vccd2
port 533 nsew power input
rlabel metal4 s 383514 568099 384134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 404514 568099 405134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 568099 426134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 488514 568000 489134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 568000 510134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 530514 465308 531134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 26514 -3814 27134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 47514 653033 48134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 68514 653033 69134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 653033 90134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 110514 653033 111134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 131514 653033 132134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 152514 653033 153134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 465308 174134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 194514 -3814 195134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 215514 652000 216134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 236514 652000 237134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 652000 258134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 278514 652000 279134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 299514 652000 300134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 320514 652000 321134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 465308 342134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 362514 465308 363134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 383514 655099 384134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 404514 655099 405134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 655099 426134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 446514 465308 447134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 467514 465308 468134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 488514 655099 489134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 655099 510134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 530514 655099 531134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 551514 -3814 552134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 572514 -3814 573134 707750 6 vccd2
port 533 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 31306 590730 31926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 52306 590730 52926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 73306 590730 73926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 94306 590730 94926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 115306 590730 115926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 136306 590730 136926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 157306 590730 157926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 178306 590730 178926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 199306 590730 199926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 220306 590730 220926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 241306 590730 241926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 283306 590730 283926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 304306 590730 304926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 325306 590730 325926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 346306 590730 346926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 367306 590730 367926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 388306 590730 388926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 409306 590730 409926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 430306 590730 430926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 451306 590730 451926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 472306 590730 472926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 493306 590730 493926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 535306 590730 535926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 556306 590730 556926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 577306 590730 577926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 598306 590730 598926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 619306 590730 619926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 640306 590730 640926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 661306 590730 661926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 682306 590730 682926 6 vdda1
port 534 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 51234 -5734 51854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 72234 -5734 72854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 -5734 93854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 114234 -5734 114854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 135234 -5734 135854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 156234 -5734 156854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 -5734 177854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 240234 -5734 240854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 -5734 261854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 282234 -5734 282854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 303234 -5734 303854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 324234 -5734 324854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 -5734 345854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 408234 -5734 408854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 -5734 429854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 450234 -5734 450854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 471234 -5734 471854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 492234 -5734 492854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 -5734 513854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 534234 -5734 534854 48000 6 vdda1
port 534 nsew power input
rlabel metal4 s 51234 135308 51854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 72234 135308 72854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 135308 93854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 114234 135308 114854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 135234 135308 135854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 156234 135308 156854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 135308 177854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 240234 135308 240854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 135308 261854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 282234 135308 282854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 303234 135308 303854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 324234 135308 324854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 135308 345854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 408234 135308 408854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 135308 429854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 450234 135308 450854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 471234 135308 471854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 492234 135308 492854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 135308 513854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 534234 135308 534854 158000 6 vdda1
port 534 nsew power input
rlabel metal4 s 51234 245308 51854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 72234 245308 72854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 245308 93854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 114234 245308 114854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 135234 245308 135854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 156234 245308 156854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 245308 177854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 240234 245308 240854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 245308 261854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 282234 245308 282854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 303234 245308 303854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 324234 245308 324854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 245308 345854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 408234 245308 408854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 245308 429854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 450234 245308 450854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 471234 245308 471854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 492234 245308 492854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 245308 513854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 534234 245308 534854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 51234 355308 51854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 72234 355308 72854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 355308 93854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 114234 355308 114854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 135234 355308 135854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 156234 355308 156854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 355308 177854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 240234 355308 240854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 355308 261854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 282234 355308 282854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 303234 355308 303854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 324234 355308 324854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 355308 345854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 408234 355308 408854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 355308 429854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 450234 355308 450854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 471234 355308 471854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 492234 355308 492854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 355308 513854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 534234 355308 534854 378000 6 vdda1
port 534 nsew power input
rlabel metal4 s 219234 -5734 219854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 240234 465308 240854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 465308 261854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 282234 465308 282854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 303234 465308 303854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 324234 465308 324854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 387234 -5734 387854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 408234 465308 408854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 465308 429854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 492234 465308 492854 514000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 465308 513854 514000 6 vdda1
port 534 nsew power input
rlabel metal4 s 51234 465308 51854 538000 6 vdda1
port 534 nsew power input
rlabel metal4 s 72234 465308 72854 538000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 465308 93854 538000 6 vdda1
port 534 nsew power input
rlabel metal4 s 114234 465308 114854 538000 6 vdda1
port 534 nsew power input
rlabel metal4 s 135234 465308 135854 538000 6 vdda1
port 534 nsew power input
rlabel metal4 s 156234 465308 156854 538000 6 vdda1
port 534 nsew power input
rlabel metal4 s 387234 568099 387854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 408234 568099 408854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 568099 429854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 492234 568000 492854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 568000 513854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 534234 465308 534854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 30234 -5734 30854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 51234 653033 51854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 72234 653033 72854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 653033 93854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 114234 653033 114854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 135234 653033 135854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 156234 653033 156854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 465308 177854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 198234 -5734 198854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 219234 652000 219854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 240234 652000 240854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 652000 261854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 282234 652000 282854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 303234 652000 303854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 324234 652000 324854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 465308 345854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 366234 -5734 366854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 387234 655099 387854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 408234 655099 408854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 655099 429854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 450234 465308 450854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 471234 465308 471854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 492234 655099 492854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 655099 513854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 534234 655099 534854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 555234 -5734 555854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 576234 -5734 576854 709670 6 vdda1
port 534 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 35026 592650 35646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 56026 592650 56646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 77026 592650 77646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 98026 592650 98646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 119026 592650 119646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 140026 592650 140646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 161026 592650 161646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 182026 592650 182646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 203026 592650 203646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 224026 592650 224646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 245026 592650 245646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 287026 592650 287646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 308026 592650 308646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 329026 592650 329646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 350026 592650 350646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 371026 592650 371646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 392026 592650 392646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 413026 592650 413646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 434026 592650 434646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 455026 592650 455646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 476026 592650 476646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 497026 592650 497646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 539026 592650 539646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 560026 592650 560646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 581026 592650 581646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 602026 592650 602646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 623026 592650 623646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 644026 592650 644646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 665026 592650 665646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 686026 592650 686646 6 vdda2
port 535 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 54954 -7654 55574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 75954 -7654 76574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 -7654 97574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 117954 -7654 118574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 138954 -7654 139574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 159954 -7654 160574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 -7654 181574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 222954 -7654 223574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 243954 -7654 244574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 -7654 265574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 285954 -7654 286574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 306954 -7654 307574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 327954 -7654 328574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 -7654 349574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 411954 -7654 412574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 -7654 433574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 453954 -7654 454574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 474954 -7654 475574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 495954 -7654 496574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 -7654 517574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 537954 -7654 538574 48000 6 vdda2
port 535 nsew power input
rlabel metal4 s 54954 135308 55574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 75954 135308 76574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 135308 97574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 117954 135308 118574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 138954 135308 139574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 159954 135308 160574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 135308 181574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 222954 135308 223574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 243954 135308 244574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 135308 265574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 285954 135308 286574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 306954 135308 307574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 327954 135308 328574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 135308 349574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 411954 135308 412574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 135308 433574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 453954 135308 454574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 474954 135308 475574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 495954 135308 496574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 135308 517574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 537954 135308 538574 158000 6 vdda2
port 535 nsew power input
rlabel metal4 s 54954 245308 55574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 75954 245308 76574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 245308 97574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 117954 245308 118574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 138954 245308 139574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 159954 245308 160574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 245308 181574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 222954 245308 223574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 243954 245308 244574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 245308 265574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 285954 245308 286574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 306954 245308 307574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 327954 245308 328574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 245308 349574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 411954 245308 412574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 245308 433574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 453954 245308 454574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 474954 245308 475574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 495954 245308 496574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 245308 517574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 537954 245308 538574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 54954 355308 55574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 75954 355308 76574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 355308 97574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 117954 355308 118574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 138954 355308 139574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 159954 355308 160574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 355308 181574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 222954 355308 223574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 243954 355308 244574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 355308 265574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 285954 355308 286574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 306954 355308 307574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 327954 355308 328574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 355308 349574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 411954 355308 412574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 355308 433574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 453954 355308 454574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 474954 355308 475574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 495954 355308 496574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 355308 517574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 537954 355308 538574 378000 6 vdda2
port 535 nsew power input
rlabel metal4 s 222954 465308 223574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 243954 465308 244574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 465308 265574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 285954 465308 286574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 306954 465308 307574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 327954 465308 328574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 390954 -7654 391574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 411954 465308 412574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 465308 433574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 474954 465308 475574 514000 6 vdda2
port 535 nsew power input
rlabel metal4 s 495954 465308 496574 514000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 465308 517574 514000 6 vdda2
port 535 nsew power input
rlabel metal4 s 54954 465308 55574 538000 6 vdda2
port 535 nsew power input
rlabel metal4 s 75954 465308 76574 538000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 465308 97574 538000 6 vdda2
port 535 nsew power input
rlabel metal4 s 117954 465308 118574 538000 6 vdda2
port 535 nsew power input
rlabel metal4 s 138954 465308 139574 538000 6 vdda2
port 535 nsew power input
rlabel metal4 s 159954 465308 160574 538000 6 vdda2
port 535 nsew power input
rlabel metal4 s 390954 568099 391574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 411954 568099 412574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 568099 433574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 474954 568000 475574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 495954 568000 496574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 568000 517574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 537954 465308 538574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 33954 -7654 34574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 54954 653033 55574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 75954 653033 76574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 653033 97574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 117954 653033 118574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 138954 653033 139574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 159954 653033 160574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 465308 181574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 201954 -7654 202574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 222954 652000 223574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 243954 652000 244574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 652000 265574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 285954 652000 286574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 306954 652000 307574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 327954 652000 328574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 465308 349574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 369954 -7654 370574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 390954 655099 391574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 411954 655099 412574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 655099 433574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 453954 465308 454574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 474954 655099 475574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 495954 655099 496574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 655099 517574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 537954 655099 538574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 558954 -7654 559574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 579954 -7654 580574 711590 6 vdda2
port 535 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 20806 590730 21426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 41806 590730 42426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 62806 590730 63426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 83806 590730 84426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 104806 590730 105426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 125806 590730 126426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 146806 590730 147426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 167806 590730 168426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 188806 590730 189426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 209806 590730 210426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 230806 590730 231426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 251806 590730 252426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 272806 590730 273426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 293806 590730 294426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 314806 590730 315426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 335806 590730 336426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 356806 590730 357426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 377806 590730 378426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 398806 590730 399426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 419806 590730 420426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 440806 590730 441426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 461806 590730 462426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 482806 590730 483426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 503806 590730 504426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 524806 590730 525426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 545806 590730 546426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 566806 590730 567426 6 vssa1
port 536 nsew ground input
rlabel metal5 s 397734 578246 440354 578866 6 vssa1
port 536 nsew ground input
rlabel metal5 s 481734 578246 524354 578866 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 587806 590730 588426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 608806 590730 609426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 629806 590730 630426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 650806 590730 651426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 671806 590730 672426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 692806 590730 693426 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 61734 -5734 62354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 82734 -5734 83354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 103734 -5734 104354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 124734 -5734 125354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 145734 -5734 146354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 166734 -5734 167354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 187734 -5734 188354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229734 -5734 230354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 250734 -5734 251354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 271734 -5734 272354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 292734 -5734 293354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 313734 -5734 314354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 334734 -5734 335354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 355734 -5734 356354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 397734 -5734 398354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 418734 -5734 419354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439734 -5734 440354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 460734 -5734 461354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 481734 -5734 482354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 502734 -5734 503354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 523734 -5734 524354 48000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 61734 135308 62354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 82734 135308 83354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 103734 135308 104354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 124734 135308 125354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 145734 135308 146354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 166734 135308 167354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 187734 135308 188354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229734 135308 230354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 250734 135308 251354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 271734 135308 272354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 292734 135308 293354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 313734 135308 314354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 334734 135308 335354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 355734 135308 356354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 397734 135308 398354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 418734 135308 419354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439734 135308 440354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 460734 135308 461354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 481734 135308 482354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 502734 135308 503354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 523734 135308 524354 158000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 61734 245308 62354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 82734 245308 83354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 103734 245308 104354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 124734 245308 125354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 145734 245308 146354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 166734 245308 167354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 187734 245308 188354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229734 245308 230354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 250734 245308 251354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 271734 245308 272354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 292734 245308 293354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 313734 245308 314354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 334734 245308 335354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 355734 245308 356354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 397734 245308 398354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 418734 245308 419354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439734 245308 440354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 460734 245308 461354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 481734 245308 482354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 502734 245308 503354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 523734 245308 524354 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 61734 355308 62354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 82734 355308 83354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 103734 355308 104354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 124734 355308 125354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 145734 355308 146354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 166734 355308 167354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 187734 355308 188354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229734 355308 230354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 250734 355308 251354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 271734 355308 272354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 292734 355308 293354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 313734 355308 314354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 334734 355308 335354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 355734 355308 356354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 397734 355308 398354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 418734 355308 419354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439734 355308 440354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 460734 355308 461354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 481734 355308 482354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 502734 355308 503354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 523734 355308 524354 378000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 208734 -5734 209354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229734 465308 230354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 250734 465308 251354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 271734 465308 272354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 292734 465308 293354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 313734 465308 314354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 397734 465308 398354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 418734 465308 419354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439734 465308 440354 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 481734 465308 482354 514000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 502734 465308 503354 514000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 523734 465308 524354 514000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 61734 465308 62354 538000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 82734 465308 83354 538000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 103734 465308 104354 538000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 124734 465308 125354 538000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 145734 465308 146354 538000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 397734 568099 398354 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 418734 568099 419354 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439734 568099 440354 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 481734 568000 482354 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 502734 568000 503354 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 523734 568000 524354 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground input
rlabel metal4 s 19734 -5734 20354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 40734 -5734 41354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 61734 653033 62354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 82734 653033 83354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 103734 653033 104354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 124734 653033 125354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 145734 653033 146354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 166734 465308 167354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 187734 465308 188354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 208734 652000 209354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229734 652000 230354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 250734 652000 251354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 271734 652000 272354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 292734 652000 293354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 313734 652000 314354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 334734 465308 335354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 355734 465308 356354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 376734 -5734 377354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 397734 655099 398354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 418734 655099 419354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439734 655099 440354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 460734 465308 461354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 481734 655099 482354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 502734 655099 503354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 523734 655099 524354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 544734 -5734 545354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 565734 -5734 566354 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 24526 592650 25146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 45526 592650 46146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 66526 592650 67146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 87526 592650 88146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 108526 592650 109146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 129526 592650 130146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 150526 592650 151146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 171526 592650 172146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 192526 592650 193146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 213526 592650 214146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 234526 592650 235146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 255526 592650 256146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 276526 592650 277146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 297526 592650 298146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 318526 592650 319146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 339526 592650 340146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 360526 592650 361146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 381526 592650 382146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 402526 592650 403146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 423526 592650 424146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 444526 592650 445146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 465526 592650 466146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 486526 592650 487146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 507526 592650 508146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 528526 592650 529146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 549526 592650 550146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 570526 592650 571146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 591526 592650 592146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 612526 592650 613146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 633526 592650 634146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 654526 592650 655146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 675526 592650 676146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 696526 592650 697146 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 65454 -7654 66074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 86454 -7654 87074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 107454 -7654 108074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 128454 -7654 129074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 149454 -7654 150074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 170454 -7654 171074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 233454 -7654 234074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 254454 -7654 255074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 275454 -7654 276074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 296454 -7654 297074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 317454 -7654 318074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 338454 -7654 339074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 359454 -7654 360074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 401454 -7654 402074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422454 -7654 423074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 443454 -7654 444074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 464454 -7654 465074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 485454 -7654 486074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 506454 -7654 507074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 527454 -7654 528074 48000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 65454 135308 66074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 86454 135308 87074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 107454 135308 108074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 128454 135308 129074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 149454 135308 150074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 170454 135308 171074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 233454 135308 234074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 254454 135308 255074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 275454 135308 276074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 296454 135308 297074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 317454 135308 318074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 338454 135308 339074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 359454 135308 360074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 401454 135308 402074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422454 135308 423074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 443454 135308 444074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 464454 135308 465074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 485454 135308 486074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 506454 135308 507074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 527454 135308 528074 158000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 65454 245308 66074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 86454 245308 87074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 107454 245308 108074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 128454 245308 129074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 149454 245308 150074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 170454 245308 171074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 233454 245308 234074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 254454 245308 255074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 275454 245308 276074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 296454 245308 297074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 317454 245308 318074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 338454 245308 339074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 359454 245308 360074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 401454 245308 402074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422454 245308 423074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 443454 245308 444074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 464454 245308 465074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 485454 245308 486074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 506454 245308 507074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 527454 245308 528074 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 65454 355308 66074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 86454 355308 87074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 107454 355308 108074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 128454 355308 129074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 149454 355308 150074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 170454 355308 171074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 233454 355308 234074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 254454 355308 255074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 275454 355308 276074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 296454 355308 297074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 317454 355308 318074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 338454 355308 339074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 359454 355308 360074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 401454 355308 402074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422454 355308 423074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 443454 355308 444074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 464454 355308 465074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 485454 355308 486074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 506454 355308 507074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 527454 355308 528074 378000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 212454 -7654 213074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 233454 465308 234074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 254454 465308 255074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 275454 465308 276074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 296454 465308 297074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 317454 465308 318074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 380454 -7654 381074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 401454 465308 402074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422454 465308 423074 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 485454 465308 486074 514000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 506454 465308 507074 514000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 65454 465308 66074 538000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 86454 465308 87074 538000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 107454 465308 108074 538000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 128454 465308 129074 538000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 149454 465308 150074 538000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 380454 568099 381074 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 401454 568099 402074 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422454 568099 423074 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 485454 568000 486074 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 506454 568000 507074 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 527454 465308 528074 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground input
rlabel metal4 s 23454 -7654 24074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 44454 -7654 45074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 65454 653033 66074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 86454 653033 87074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 107454 653033 108074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 128454 653033 129074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 149454 653033 150074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 170454 465308 171074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 191454 -7654 192074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 212454 652000 213074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 233454 652000 234074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 254454 652000 255074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 275454 652000 276074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 296454 652000 297074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 317454 652000 318074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 338454 465308 339074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 359454 465308 360074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 380454 655099 381074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 401454 655099 402074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422454 655099 423074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 443454 465308 444074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 464454 465308 465074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 485454 655099 486074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 506454 655099 507074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 527454 655099 528074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 548454 -7654 549074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 569454 -7654 570074 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 13366 586890 13986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 34366 586890 34986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 55366 586890 55986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 76366 586890 76986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 97366 586890 97986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 118366 586890 118986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 139366 586890 139986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 160366 586890 160986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 181366 586890 181986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 202366 586890 202986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 223366 586890 223986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 244366 586890 244986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 265366 586890 265986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 286366 586890 286986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 307366 586890 307986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 328366 586890 328986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 349366 586890 349986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 370366 586890 370986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 391366 586890 391986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 412366 586890 412986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 433366 586890 433986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 454366 586890 454986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 475366 586890 475986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 496366 586890 496986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 517366 586890 517986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 538366 586890 538986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 559366 586890 559986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 580366 586890 580986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 601366 586890 601986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 622366 586890 622986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 643366 586890 643986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 664366 586890 664986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 685366 586890 685986 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 54294 -1894 54914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 75294 -1894 75914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 96294 -1894 96914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 117294 -1894 117914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 138294 -1894 138914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 159294 -1894 159914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 180294 -1894 180914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 243294 -1894 243914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 264294 -1894 264914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 285294 -1894 285914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 306294 -1894 306914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 327294 -1894 327914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 348294 -1894 348914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411294 -1894 411914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 432294 -1894 432914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 453294 -1894 453914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 474294 -1894 474914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 495294 -1894 495914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 516294 -1894 516914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 537294 -1894 537914 48000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 54294 135308 54914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 75294 135308 75914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 96294 135308 96914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 117294 135308 117914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 138294 135308 138914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 159294 135308 159914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 180294 135308 180914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 243294 135308 243914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 264294 135308 264914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 285294 135308 285914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 306294 135308 306914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 327294 135308 327914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 348294 135308 348914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411294 135308 411914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 432294 135308 432914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 453294 135308 453914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 474294 135308 474914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 495294 135308 495914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 516294 135308 516914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 537294 135308 537914 158000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 54294 245308 54914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 75294 245308 75914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 96294 245308 96914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 117294 245308 117914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 138294 245308 138914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 159294 245308 159914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 180294 245308 180914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 243294 245308 243914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 264294 245308 264914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 285294 245308 285914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 306294 245308 306914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 327294 245308 327914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 348294 245308 348914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411294 245308 411914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 432294 245308 432914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 453294 245308 453914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 474294 245308 474914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 495294 245308 495914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 516294 245308 516914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 537294 245308 537914 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 54294 355308 54914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 75294 355308 75914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 96294 355308 96914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 117294 355308 117914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 138294 355308 138914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 159294 355308 159914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 180294 355308 180914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 243294 355308 243914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 264294 355308 264914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 285294 355308 285914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 306294 355308 306914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 327294 355308 327914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 348294 355308 348914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411294 355308 411914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 432294 355308 432914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 453294 355308 453914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 474294 355308 474914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 495294 355308 495914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 516294 355308 516914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 537294 355308 537914 378000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 222294 -1894 222914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 243294 465308 243914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 264294 465308 264914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 285294 465308 285914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 306294 465308 306914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 327294 465308 327914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 390294 -1894 390914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411294 465308 411914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 432294 465308 432914 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 474294 465308 474914 514000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 495294 465308 495914 514000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 516294 465308 516914 514000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 54294 465308 54914 538000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 75294 465308 75914 538000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 96294 465308 96914 538000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 117294 465308 117914 538000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 138294 465308 138914 538000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 159294 465308 159914 538000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 390294 568099 390914 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411294 568099 411914 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 432294 568099 432914 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 474294 568000 474914 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 495294 568000 495914 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 516294 568000 516914 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 537294 465308 537914 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground input
rlabel metal4 s 12294 -1894 12914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 33294 -1894 33914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 54294 653033 54914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 75294 653033 75914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 96294 653033 96914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 117294 653033 117914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 138294 653033 138914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 159294 653033 159914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 180294 465308 180914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 201294 -1894 201914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 222294 652000 222914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 243294 652000 243914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 264294 652000 264914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 285294 652000 285914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 306294 652000 306914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 327294 652000 327914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 348294 465308 348914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 369294 -1894 369914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 390294 655099 390914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411294 655099 411914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 432294 655099 432914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 453294 465308 453914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 474294 655099 474914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 495294 655099 495914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 516294 655099 516914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 537294 655099 537914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 558294 -1894 558914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 579294 -1894 579914 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 17086 588810 17706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 38086 588810 38706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 59086 588810 59706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 80086 588810 80706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 101086 588810 101706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 122086 588810 122706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 143086 588810 143706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 164086 588810 164706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 185086 588810 185706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 206086 588810 206706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 227086 588810 227706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 248086 588810 248706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 269086 588810 269706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 290086 588810 290706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 311086 588810 311706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 332086 588810 332706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 353086 588810 353706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 374086 588810 374706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 395086 588810 395706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 416086 588810 416706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 437086 588810 437706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 458086 588810 458706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 479086 588810 479706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 500086 588810 500706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 521086 588810 521706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 542086 588810 542706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 563086 588810 563706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 584086 588810 584706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 605086 588810 605706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 626086 588810 626706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 647086 588810 647706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 668086 588810 668706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 689086 588810 689706 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 58014 -3814 58634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 79014 -3814 79634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 100014 -3814 100634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 121014 -3814 121634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 142014 -3814 142634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 163014 -3814 163634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 184014 -3814 184634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 226014 -3814 226634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 247014 -3814 247634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 268014 -3814 268634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 289014 -3814 289634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 310014 -3814 310634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 331014 -3814 331634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 352014 -3814 352634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415014 -3814 415634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 436014 -3814 436634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 457014 -3814 457634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 478014 -3814 478634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 499014 -3814 499634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 520014 -3814 520634 48000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 58014 135308 58634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 79014 135308 79634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 100014 135308 100634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 121014 135308 121634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 142014 135308 142634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 163014 135308 163634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 184014 135308 184634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 226014 135308 226634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 247014 135308 247634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 268014 135308 268634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 289014 135308 289634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 310014 135308 310634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 331014 135308 331634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 352014 135308 352634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415014 135308 415634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 436014 135308 436634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 457014 135308 457634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 478014 135308 478634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 499014 135308 499634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 520014 135308 520634 158000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 58014 245308 58634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 79014 245308 79634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 100014 245308 100634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 121014 245308 121634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 142014 245308 142634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 163014 245308 163634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 184014 245308 184634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 226014 245308 226634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 247014 245308 247634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 268014 245308 268634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 289014 245308 289634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 310014 245308 310634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 331014 245308 331634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 352014 245308 352634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415014 245308 415634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 436014 245308 436634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 457014 245308 457634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 478014 245308 478634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 499014 245308 499634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 520014 245308 520634 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 58014 355308 58634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 79014 355308 79634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 100014 355308 100634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 121014 355308 121634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 142014 355308 142634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 163014 355308 163634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 184014 355308 184634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 226014 355308 226634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 247014 355308 247634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 268014 355308 268634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 289014 355308 289634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 310014 355308 310634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 331014 355308 331634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 352014 355308 352634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415014 355308 415634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 436014 355308 436634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 457014 355308 457634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 478014 355308 478634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 499014 355308 499634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 520014 355308 520634 378000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 226014 465308 226634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 247014 465308 247634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 268014 465308 268634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 289014 465308 289634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 310014 465308 310634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 331014 465308 331634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 394014 -3814 394634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415014 465308 415634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 436014 465308 436634 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 478014 465308 478634 514000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 499014 465308 499634 514000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 520014 465308 520634 514000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 58014 465308 58634 538000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 79014 465308 79634 538000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 100014 465308 100634 538000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 121014 465308 121634 538000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 142014 465308 142634 538000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 394014 568099 394634 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415014 568099 415634 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 436014 568099 436634 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 478014 568000 478634 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 499014 568000 499634 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 520014 568000 520634 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground input
rlabel metal4 s 16014 -3814 16634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 37014 -3814 37634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 58014 653033 58634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 79014 653033 79634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 100014 653033 100634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 121014 653033 121634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 142014 653033 142634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 163014 465308 163634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 184014 465308 184634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 205014 -3814 205634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 226014 652000 226634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 247014 652000 247634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 268014 652000 268634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 289014 652000 289634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 310014 652000 310634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 331014 652000 331634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 352014 465308 352634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 373014 -3814 373634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 394014 655099 394634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415014 655099 415634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 436014 655099 436634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 457014 465308 457634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 478014 655099 478634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 499014 655099 499634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 520014 655099 520634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 541014 -3814 541634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 562014 -3814 562634 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 95132510
string GDS_FILE /home/burak/asic_tools/caravel_vscpu3x/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 90644312
<< end >>

