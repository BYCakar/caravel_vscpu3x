VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO main_controller
  CLASS BLOCK ;
  FOREIGN main_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 735.000 ;
  PIN agent_1_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 445.440 600.000 446.040 ;
    END
  END agent_1_mem_ctrl_addr[0]
  PIN agent_1_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 472.640 600.000 473.240 ;
    END
  END agent_1_mem_ctrl_addr[10]
  PIN agent_1_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 475.360 600.000 475.960 ;
    END
  END agent_1_mem_ctrl_addr[11]
  PIN agent_1_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 478.080 600.000 478.680 ;
    END
  END agent_1_mem_ctrl_addr[12]
  PIN agent_1_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 480.800 600.000 481.400 ;
    END
  END agent_1_mem_ctrl_addr[13]
  PIN agent_1_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 448.160 600.000 448.760 ;
    END
  END agent_1_mem_ctrl_addr[1]
  PIN agent_1_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 450.880 600.000 451.480 ;
    END
  END agent_1_mem_ctrl_addr[2]
  PIN agent_1_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 453.600 600.000 454.200 ;
    END
  END agent_1_mem_ctrl_addr[3]
  PIN agent_1_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 456.320 600.000 456.920 ;
    END
  END agent_1_mem_ctrl_addr[4]
  PIN agent_1_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 459.040 600.000 459.640 ;
    END
  END agent_1_mem_ctrl_addr[5]
  PIN agent_1_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 461.760 600.000 462.360 ;
    END
  END agent_1_mem_ctrl_addr[6]
  PIN agent_1_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 464.480 600.000 465.080 ;
    END
  END agent_1_mem_ctrl_addr[7]
  PIN agent_1_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 467.200 600.000 467.800 ;
    END
  END agent_1_mem_ctrl_addr[8]
  PIN agent_1_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 469.920 600.000 470.520 ;
    END
  END agent_1_mem_ctrl_addr[9]
  PIN agent_1_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 483.520 600.000 484.120 ;
    END
  END agent_1_mem_ctrl_in[0]
  PIN agent_1_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 511.400 600.000 512.000 ;
    END
  END agent_1_mem_ctrl_in[10]
  PIN agent_1_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 514.120 600.000 514.720 ;
    END
  END agent_1_mem_ctrl_in[11]
  PIN agent_1_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 516.840 600.000 517.440 ;
    END
  END agent_1_mem_ctrl_in[12]
  PIN agent_1_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 519.560 600.000 520.160 ;
    END
  END agent_1_mem_ctrl_in[13]
  PIN agent_1_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 522.280 600.000 522.880 ;
    END
  END agent_1_mem_ctrl_in[14]
  PIN agent_1_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 525.000 600.000 525.600 ;
    END
  END agent_1_mem_ctrl_in[15]
  PIN agent_1_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 527.720 600.000 528.320 ;
    END
  END agent_1_mem_ctrl_in[16]
  PIN agent_1_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 530.440 600.000 531.040 ;
    END
  END agent_1_mem_ctrl_in[17]
  PIN agent_1_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 533.160 600.000 533.760 ;
    END
  END agent_1_mem_ctrl_in[18]
  PIN agent_1_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 535.880 600.000 536.480 ;
    END
  END agent_1_mem_ctrl_in[19]
  PIN agent_1_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 486.240 600.000 486.840 ;
    END
  END agent_1_mem_ctrl_in[1]
  PIN agent_1_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 538.600 600.000 539.200 ;
    END
  END agent_1_mem_ctrl_in[20]
  PIN agent_1_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 541.320 600.000 541.920 ;
    END
  END agent_1_mem_ctrl_in[21]
  PIN agent_1_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 544.040 600.000 544.640 ;
    END
  END agent_1_mem_ctrl_in[22]
  PIN agent_1_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 546.760 600.000 547.360 ;
    END
  END agent_1_mem_ctrl_in[23]
  PIN agent_1_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 549.480 600.000 550.080 ;
    END
  END agent_1_mem_ctrl_in[24]
  PIN agent_1_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 552.200 600.000 552.800 ;
    END
  END agent_1_mem_ctrl_in[25]
  PIN agent_1_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 554.920 600.000 555.520 ;
    END
  END agent_1_mem_ctrl_in[26]
  PIN agent_1_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 557.640 600.000 558.240 ;
    END
  END agent_1_mem_ctrl_in[27]
  PIN agent_1_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 560.360 600.000 560.960 ;
    END
  END agent_1_mem_ctrl_in[28]
  PIN agent_1_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 563.080 600.000 563.680 ;
    END
  END agent_1_mem_ctrl_in[29]
  PIN agent_1_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 488.960 600.000 489.560 ;
    END
  END agent_1_mem_ctrl_in[2]
  PIN agent_1_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 565.800 600.000 566.400 ;
    END
  END agent_1_mem_ctrl_in[30]
  PIN agent_1_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 568.520 600.000 569.120 ;
    END
  END agent_1_mem_ctrl_in[31]
  PIN agent_1_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 492.360 600.000 492.960 ;
    END
  END agent_1_mem_ctrl_in[3]
  PIN agent_1_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 495.080 600.000 495.680 ;
    END
  END agent_1_mem_ctrl_in[4]
  PIN agent_1_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 497.800 600.000 498.400 ;
    END
  END agent_1_mem_ctrl_in[5]
  PIN agent_1_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 500.520 600.000 501.120 ;
    END
  END agent_1_mem_ctrl_in[6]
  PIN agent_1_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 503.240 600.000 503.840 ;
    END
  END agent_1_mem_ctrl_in[7]
  PIN agent_1_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 505.960 600.000 506.560 ;
    END
  END agent_1_mem_ctrl_in[8]
  PIN agent_1_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 508.680 600.000 509.280 ;
    END
  END agent_1_mem_ctrl_in[9]
  PIN agent_1_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 571.240 600.000 571.840 ;
    END
  END agent_1_mem_ctrl_out[0]
  PIN agent_1_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 599.120 600.000 599.720 ;
    END
  END agent_1_mem_ctrl_out[10]
  PIN agent_1_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 601.840 600.000 602.440 ;
    END
  END agent_1_mem_ctrl_out[11]
  PIN agent_1_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 604.560 600.000 605.160 ;
    END
  END agent_1_mem_ctrl_out[12]
  PIN agent_1_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 607.280 600.000 607.880 ;
    END
  END agent_1_mem_ctrl_out[13]
  PIN agent_1_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 610.000 600.000 610.600 ;
    END
  END agent_1_mem_ctrl_out[14]
  PIN agent_1_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 612.720 600.000 613.320 ;
    END
  END agent_1_mem_ctrl_out[15]
  PIN agent_1_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 615.440 600.000 616.040 ;
    END
  END agent_1_mem_ctrl_out[16]
  PIN agent_1_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 618.160 600.000 618.760 ;
    END
  END agent_1_mem_ctrl_out[17]
  PIN agent_1_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 620.880 600.000 621.480 ;
    END
  END agent_1_mem_ctrl_out[18]
  PIN agent_1_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 623.600 600.000 624.200 ;
    END
  END agent_1_mem_ctrl_out[19]
  PIN agent_1_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 574.640 600.000 575.240 ;
    END
  END agent_1_mem_ctrl_out[1]
  PIN agent_1_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 626.320 600.000 626.920 ;
    END
  END agent_1_mem_ctrl_out[20]
  PIN agent_1_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 629.040 600.000 629.640 ;
    END
  END agent_1_mem_ctrl_out[21]
  PIN agent_1_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 631.760 600.000 632.360 ;
    END
  END agent_1_mem_ctrl_out[22]
  PIN agent_1_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 634.480 600.000 635.080 ;
    END
  END agent_1_mem_ctrl_out[23]
  PIN agent_1_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 637.200 600.000 637.800 ;
    END
  END agent_1_mem_ctrl_out[24]
  PIN agent_1_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 639.920 600.000 640.520 ;
    END
  END agent_1_mem_ctrl_out[25]
  PIN agent_1_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 642.640 600.000 643.240 ;
    END
  END agent_1_mem_ctrl_out[26]
  PIN agent_1_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 645.360 600.000 645.960 ;
    END
  END agent_1_mem_ctrl_out[27]
  PIN agent_1_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 648.080 600.000 648.680 ;
    END
  END agent_1_mem_ctrl_out[28]
  PIN agent_1_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 650.800 600.000 651.400 ;
    END
  END agent_1_mem_ctrl_out[29]
  PIN agent_1_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 577.360 600.000 577.960 ;
    END
  END agent_1_mem_ctrl_out[2]
  PIN agent_1_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 653.520 600.000 654.120 ;
    END
  END agent_1_mem_ctrl_out[30]
  PIN agent_1_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 656.920 600.000 657.520 ;
    END
  END agent_1_mem_ctrl_out[31]
  PIN agent_1_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 580.080 600.000 580.680 ;
    END
  END agent_1_mem_ctrl_out[3]
  PIN agent_1_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 582.800 600.000 583.400 ;
    END
  END agent_1_mem_ctrl_out[4]
  PIN agent_1_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 585.520 600.000 586.120 ;
    END
  END agent_1_mem_ctrl_out[5]
  PIN agent_1_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 588.240 600.000 588.840 ;
    END
  END agent_1_mem_ctrl_out[6]
  PIN agent_1_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 590.960 600.000 591.560 ;
    END
  END agent_1_mem_ctrl_out[7]
  PIN agent_1_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 593.680 600.000 594.280 ;
    END
  END agent_1_mem_ctrl_out[8]
  PIN agent_1_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 596.400 600.000 597.000 ;
    END
  END agent_1_mem_ctrl_out[9]
  PIN agent_1_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 659.640 600.000 660.240 ;
    END
  END agent_1_mem_ctrl_req
  PIN agent_1_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 662.360 600.000 662.960 ;
    END
  END agent_1_mem_ctrl_vld
  PIN agent_1_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 665.080 600.000 665.680 ;
    END
  END agent_1_mem_ctrl_we
  PIN agent_1_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END agent_1_sram0_csb0
  PIN agent_1_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END agent_1_sram0_dout0[0]
  PIN agent_1_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END agent_1_sram0_dout0[10]
  PIN agent_1_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END agent_1_sram0_dout0[11]
  PIN agent_1_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END agent_1_sram0_dout0[12]
  PIN agent_1_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END agent_1_sram0_dout0[13]
  PIN agent_1_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END agent_1_sram0_dout0[14]
  PIN agent_1_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END agent_1_sram0_dout0[15]
  PIN agent_1_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END agent_1_sram0_dout0[16]
  PIN agent_1_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END agent_1_sram0_dout0[17]
  PIN agent_1_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END agent_1_sram0_dout0[18]
  PIN agent_1_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END agent_1_sram0_dout0[19]
  PIN agent_1_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END agent_1_sram0_dout0[1]
  PIN agent_1_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END agent_1_sram0_dout0[20]
  PIN agent_1_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END agent_1_sram0_dout0[21]
  PIN agent_1_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END agent_1_sram0_dout0[22]
  PIN agent_1_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END agent_1_sram0_dout0[23]
  PIN agent_1_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END agent_1_sram0_dout0[24]
  PIN agent_1_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END agent_1_sram0_dout0[25]
  PIN agent_1_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END agent_1_sram0_dout0[26]
  PIN agent_1_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END agent_1_sram0_dout0[27]
  PIN agent_1_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END agent_1_sram0_dout0[28]
  PIN agent_1_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END agent_1_sram0_dout0[29]
  PIN agent_1_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END agent_1_sram0_dout0[2]
  PIN agent_1_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END agent_1_sram0_dout0[30]
  PIN agent_1_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END agent_1_sram0_dout0[31]
  PIN agent_1_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END agent_1_sram0_dout0[3]
  PIN agent_1_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END agent_1_sram0_dout0[4]
  PIN agent_1_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END agent_1_sram0_dout0[5]
  PIN agent_1_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END agent_1_sram0_dout0[6]
  PIN agent_1_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END agent_1_sram0_dout0[7]
  PIN agent_1_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END agent_1_sram0_dout0[8]
  PIN agent_1_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END agent_1_sram0_dout0[9]
  PIN agent_1_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END agent_1_sram0_web0
  PIN agent_1_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END agent_1_sram1_csb0
  PIN agent_1_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END agent_1_sram1_dout0[0]
  PIN agent_1_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END agent_1_sram1_dout0[10]
  PIN agent_1_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END agent_1_sram1_dout0[11]
  PIN agent_1_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END agent_1_sram1_dout0[12]
  PIN agent_1_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END agent_1_sram1_dout0[13]
  PIN agent_1_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END agent_1_sram1_dout0[14]
  PIN agent_1_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END agent_1_sram1_dout0[15]
  PIN agent_1_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END agent_1_sram1_dout0[16]
  PIN agent_1_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END agent_1_sram1_dout0[17]
  PIN agent_1_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END agent_1_sram1_dout0[18]
  PIN agent_1_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END agent_1_sram1_dout0[19]
  PIN agent_1_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END agent_1_sram1_dout0[1]
  PIN agent_1_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END agent_1_sram1_dout0[20]
  PIN agent_1_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END agent_1_sram1_dout0[21]
  PIN agent_1_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END agent_1_sram1_dout0[22]
  PIN agent_1_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END agent_1_sram1_dout0[23]
  PIN agent_1_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END agent_1_sram1_dout0[24]
  PIN agent_1_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END agent_1_sram1_dout0[25]
  PIN agent_1_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END agent_1_sram1_dout0[26]
  PIN agent_1_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END agent_1_sram1_dout0[27]
  PIN agent_1_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END agent_1_sram1_dout0[28]
  PIN agent_1_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END agent_1_sram1_dout0[29]
  PIN agent_1_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END agent_1_sram1_dout0[2]
  PIN agent_1_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END agent_1_sram1_dout0[30]
  PIN agent_1_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END agent_1_sram1_dout0[31]
  PIN agent_1_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END agent_1_sram1_dout0[3]
  PIN agent_1_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END agent_1_sram1_dout0[4]
  PIN agent_1_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END agent_1_sram1_dout0[5]
  PIN agent_1_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END agent_1_sram1_dout0[6]
  PIN agent_1_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END agent_1_sram1_dout0[7]
  PIN agent_1_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END agent_1_sram1_dout0[8]
  PIN agent_1_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END agent_1_sram1_dout0[9]
  PIN agent_1_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END agent_1_sram1_web0
  PIN agent_1_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END agent_1_sram2_csb0
  PIN agent_1_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END agent_1_sram2_dout0[0]
  PIN agent_1_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END agent_1_sram2_dout0[10]
  PIN agent_1_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END agent_1_sram2_dout0[11]
  PIN agent_1_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END agent_1_sram2_dout0[12]
  PIN agent_1_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END agent_1_sram2_dout0[13]
  PIN agent_1_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END agent_1_sram2_dout0[14]
  PIN agent_1_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END agent_1_sram2_dout0[15]
  PIN agent_1_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END agent_1_sram2_dout0[16]
  PIN agent_1_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END agent_1_sram2_dout0[17]
  PIN agent_1_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END agent_1_sram2_dout0[18]
  PIN agent_1_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END agent_1_sram2_dout0[19]
  PIN agent_1_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END agent_1_sram2_dout0[1]
  PIN agent_1_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 551.520 4.000 552.120 ;
    END
  END agent_1_sram2_dout0[20]
  PIN agent_1_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END agent_1_sram2_dout0[21]
  PIN agent_1_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END agent_1_sram2_dout0[22]
  PIN agent_1_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END agent_1_sram2_dout0[23]
  PIN agent_1_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.120 4.000 565.720 ;
    END
  END agent_1_sram2_dout0[24]
  PIN agent_1_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END agent_1_sram2_dout0[25]
  PIN agent_1_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END agent_1_sram2_dout0[26]
  PIN agent_1_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END agent_1_sram2_dout0[27]
  PIN agent_1_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END agent_1_sram2_dout0[28]
  PIN agent_1_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END agent_1_sram2_dout0[29]
  PIN agent_1_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END agent_1_sram2_dout0[2]
  PIN agent_1_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END agent_1_sram2_dout0[30]
  PIN agent_1_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END agent_1_sram2_dout0[31]
  PIN agent_1_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END agent_1_sram2_dout0[3]
  PIN agent_1_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END agent_1_sram2_dout0[4]
  PIN agent_1_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END agent_1_sram2_dout0[5]
  PIN agent_1_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END agent_1_sram2_dout0[6]
  PIN agent_1_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END agent_1_sram2_dout0[7]
  PIN agent_1_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.720 4.000 511.320 ;
    END
  END agent_1_sram2_dout0[8]
  PIN agent_1_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END agent_1_sram2_dout0[9]
  PIN agent_1_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END agent_1_sram2_web0
  PIN agent_1_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END agent_1_sram_comm_addr0[0]
  PIN agent_1_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END agent_1_sram_comm_addr0[1]
  PIN agent_1_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END agent_1_sram_comm_addr0[2]
  PIN agent_1_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END agent_1_sram_comm_addr0[3]
  PIN agent_1_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END agent_1_sram_comm_addr0[4]
  PIN agent_1_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END agent_1_sram_comm_addr0[5]
  PIN agent_1_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END agent_1_sram_comm_addr0[6]
  PIN agent_1_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END agent_1_sram_comm_addr0[7]
  PIN agent_1_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END agent_1_sram_comm_addr0[8]
  PIN agent_1_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END agent_1_sram_comm_din0[0]
  PIN agent_1_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END agent_1_sram_comm_din0[10]
  PIN agent_1_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END agent_1_sram_comm_din0[11]
  PIN agent_1_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END agent_1_sram_comm_din0[12]
  PIN agent_1_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.200 4.000 671.800 ;
    END
  END agent_1_sram_comm_din0[13]
  PIN agent_1_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END agent_1_sram_comm_din0[14]
  PIN agent_1_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END agent_1_sram_comm_din0[15]
  PIN agent_1_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END agent_1_sram_comm_din0[16]
  PIN agent_1_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END agent_1_sram_comm_din0[17]
  PIN agent_1_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END agent_1_sram_comm_din0[18]
  PIN agent_1_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END agent_1_sram_comm_din0[19]
  PIN agent_1_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END agent_1_sram_comm_din0[1]
  PIN agent_1_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END agent_1_sram_comm_din0[20]
  PIN agent_1_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 698.400 4.000 699.000 ;
    END
  END agent_1_sram_comm_din0[21]
  PIN agent_1_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END agent_1_sram_comm_din0[22]
  PIN agent_1_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END agent_1_sram_comm_din0[23]
  PIN agent_1_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END agent_1_sram_comm_din0[24]
  PIN agent_1_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END agent_1_sram_comm_din0[25]
  PIN agent_1_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END agent_1_sram_comm_din0[26]
  PIN agent_1_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.800 4.000 719.400 ;
    END
  END agent_1_sram_comm_din0[27]
  PIN agent_1_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END agent_1_sram_comm_din0[28]
  PIN agent_1_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END agent_1_sram_comm_din0[29]
  PIN agent_1_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END agent_1_sram_comm_din0[2]
  PIN agent_1_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 4.000 729.600 ;
    END
  END agent_1_sram_comm_din0[30]
  PIN agent_1_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 732.400 4.000 733.000 ;
    END
  END agent_1_sram_comm_din0[31]
  PIN agent_1_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.200 4.000 637.800 ;
    END
  END agent_1_sram_comm_din0[3]
  PIN agent_1_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END agent_1_sram_comm_din0[4]
  PIN agent_1_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.000 4.000 644.600 ;
    END
  END agent_1_sram_comm_din0[5]
  PIN agent_1_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END agent_1_sram_comm_din0[6]
  PIN agent_1_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END agent_1_sram_comm_din0[7]
  PIN agent_1_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END agent_1_sram_comm_din0[8]
  PIN agent_1_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END agent_1_sram_comm_din0[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END clk
  PIN cm_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 1.400 600.000 2.000 ;
    END
  END cm_mem_ctrl_addr[0]
  PIN cm_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 28.600 600.000 29.200 ;
    END
  END cm_mem_ctrl_addr[10]
  PIN cm_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 31.320 600.000 31.920 ;
    END
  END cm_mem_ctrl_addr[11]
  PIN cm_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 34.040 600.000 34.640 ;
    END
  END cm_mem_ctrl_addr[12]
  PIN cm_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 36.760 600.000 37.360 ;
    END
  END cm_mem_ctrl_addr[13]
  PIN cm_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 4.120 600.000 4.720 ;
    END
  END cm_mem_ctrl_addr[1]
  PIN cm_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 6.840 600.000 7.440 ;
    END
  END cm_mem_ctrl_addr[2]
  PIN cm_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 9.560 600.000 10.160 ;
    END
  END cm_mem_ctrl_addr[3]
  PIN cm_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 12.280 600.000 12.880 ;
    END
  END cm_mem_ctrl_addr[4]
  PIN cm_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 15.000 600.000 15.600 ;
    END
  END cm_mem_ctrl_addr[5]
  PIN cm_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 17.720 600.000 18.320 ;
    END
  END cm_mem_ctrl_addr[6]
  PIN cm_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 20.440 600.000 21.040 ;
    END
  END cm_mem_ctrl_addr[7]
  PIN cm_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 23.160 600.000 23.760 ;
    END
  END cm_mem_ctrl_addr[8]
  PIN cm_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 25.880 600.000 26.480 ;
    END
  END cm_mem_ctrl_addr[9]
  PIN cm_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 39.480 600.000 40.080 ;
    END
  END cm_mem_ctrl_in[0]
  PIN cm_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 66.680 600.000 67.280 ;
    END
  END cm_mem_ctrl_in[10]
  PIN cm_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 69.400 600.000 70.000 ;
    END
  END cm_mem_ctrl_in[11]
  PIN cm_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 72.120 600.000 72.720 ;
    END
  END cm_mem_ctrl_in[12]
  PIN cm_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 74.840 600.000 75.440 ;
    END
  END cm_mem_ctrl_in[13]
  PIN cm_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 77.560 600.000 78.160 ;
    END
  END cm_mem_ctrl_in[14]
  PIN cm_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 80.280 600.000 80.880 ;
    END
  END cm_mem_ctrl_in[15]
  PIN cm_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 83.680 600.000 84.280 ;
    END
  END cm_mem_ctrl_in[16]
  PIN cm_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 86.400 600.000 87.000 ;
    END
  END cm_mem_ctrl_in[17]
  PIN cm_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 89.120 600.000 89.720 ;
    END
  END cm_mem_ctrl_in[18]
  PIN cm_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 91.840 600.000 92.440 ;
    END
  END cm_mem_ctrl_in[19]
  PIN cm_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 42.200 600.000 42.800 ;
    END
  END cm_mem_ctrl_in[1]
  PIN cm_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 94.560 600.000 95.160 ;
    END
  END cm_mem_ctrl_in[20]
  PIN cm_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 97.280 600.000 97.880 ;
    END
  END cm_mem_ctrl_in[21]
  PIN cm_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 100.000 600.000 100.600 ;
    END
  END cm_mem_ctrl_in[22]
  PIN cm_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 102.720 600.000 103.320 ;
    END
  END cm_mem_ctrl_in[23]
  PIN cm_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 105.440 600.000 106.040 ;
    END
  END cm_mem_ctrl_in[24]
  PIN cm_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 108.160 600.000 108.760 ;
    END
  END cm_mem_ctrl_in[25]
  PIN cm_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 110.880 600.000 111.480 ;
    END
  END cm_mem_ctrl_in[26]
  PIN cm_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 113.600 600.000 114.200 ;
    END
  END cm_mem_ctrl_in[27]
  PIN cm_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 116.320 600.000 116.920 ;
    END
  END cm_mem_ctrl_in[28]
  PIN cm_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 119.040 600.000 119.640 ;
    END
  END cm_mem_ctrl_in[29]
  PIN cm_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 44.920 600.000 45.520 ;
    END
  END cm_mem_ctrl_in[2]
  PIN cm_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 121.760 600.000 122.360 ;
    END
  END cm_mem_ctrl_in[30]
  PIN cm_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 124.480 600.000 125.080 ;
    END
  END cm_mem_ctrl_in[31]
  PIN cm_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 47.640 600.000 48.240 ;
    END
  END cm_mem_ctrl_in[3]
  PIN cm_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 50.360 600.000 50.960 ;
    END
  END cm_mem_ctrl_in[4]
  PIN cm_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 53.080 600.000 53.680 ;
    END
  END cm_mem_ctrl_in[5]
  PIN cm_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 55.800 600.000 56.400 ;
    END
  END cm_mem_ctrl_in[6]
  PIN cm_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 58.520 600.000 59.120 ;
    END
  END cm_mem_ctrl_in[7]
  PIN cm_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 61.240 600.000 61.840 ;
    END
  END cm_mem_ctrl_in[8]
  PIN cm_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 63.960 600.000 64.560 ;
    END
  END cm_mem_ctrl_in[9]
  PIN cm_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 127.200 600.000 127.800 ;
    END
  END cm_mem_ctrl_out[0]
  PIN cm_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 154.400 600.000 155.000 ;
    END
  END cm_mem_ctrl_out[10]
  PIN cm_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 157.120 600.000 157.720 ;
    END
  END cm_mem_ctrl_out[11]
  PIN cm_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 159.840 600.000 160.440 ;
    END
  END cm_mem_ctrl_out[12]
  PIN cm_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 162.560 600.000 163.160 ;
    END
  END cm_mem_ctrl_out[13]
  PIN cm_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 165.960 600.000 166.560 ;
    END
  END cm_mem_ctrl_out[14]
  PIN cm_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 168.680 600.000 169.280 ;
    END
  END cm_mem_ctrl_out[15]
  PIN cm_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 171.400 600.000 172.000 ;
    END
  END cm_mem_ctrl_out[16]
  PIN cm_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 174.120 600.000 174.720 ;
    END
  END cm_mem_ctrl_out[17]
  PIN cm_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 176.840 600.000 177.440 ;
    END
  END cm_mem_ctrl_out[18]
  PIN cm_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 179.560 600.000 180.160 ;
    END
  END cm_mem_ctrl_out[19]
  PIN cm_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 129.920 600.000 130.520 ;
    END
  END cm_mem_ctrl_out[1]
  PIN cm_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 182.280 600.000 182.880 ;
    END
  END cm_mem_ctrl_out[20]
  PIN cm_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 185.000 600.000 185.600 ;
    END
  END cm_mem_ctrl_out[21]
  PIN cm_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 187.720 600.000 188.320 ;
    END
  END cm_mem_ctrl_out[22]
  PIN cm_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 190.440 600.000 191.040 ;
    END
  END cm_mem_ctrl_out[23]
  PIN cm_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 193.160 600.000 193.760 ;
    END
  END cm_mem_ctrl_out[24]
  PIN cm_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 195.880 600.000 196.480 ;
    END
  END cm_mem_ctrl_out[25]
  PIN cm_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 198.600 600.000 199.200 ;
    END
  END cm_mem_ctrl_out[26]
  PIN cm_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 201.320 600.000 201.920 ;
    END
  END cm_mem_ctrl_out[27]
  PIN cm_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 204.040 600.000 204.640 ;
    END
  END cm_mem_ctrl_out[28]
  PIN cm_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 206.760 600.000 207.360 ;
    END
  END cm_mem_ctrl_out[29]
  PIN cm_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 132.640 600.000 133.240 ;
    END
  END cm_mem_ctrl_out[2]
  PIN cm_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 209.480 600.000 210.080 ;
    END
  END cm_mem_ctrl_out[30]
  PIN cm_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 212.200 600.000 212.800 ;
    END
  END cm_mem_ctrl_out[31]
  PIN cm_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 135.360 600.000 135.960 ;
    END
  END cm_mem_ctrl_out[3]
  PIN cm_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 138.080 600.000 138.680 ;
    END
  END cm_mem_ctrl_out[4]
  PIN cm_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 140.800 600.000 141.400 ;
    END
  END cm_mem_ctrl_out[5]
  PIN cm_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 143.520 600.000 144.120 ;
    END
  END cm_mem_ctrl_out[6]
  PIN cm_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 146.240 600.000 146.840 ;
    END
  END cm_mem_ctrl_out[7]
  PIN cm_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 148.960 600.000 149.560 ;
    END
  END cm_mem_ctrl_out[8]
  PIN cm_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 151.680 600.000 152.280 ;
    END
  END cm_mem_ctrl_out[9]
  PIN cm_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 214.920 600.000 215.520 ;
    END
  END cm_mem_ctrl_req
  PIN cm_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 217.640 600.000 218.240 ;
    END
  END cm_mem_ctrl_vld
  PIN cm_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 220.360 600.000 220.960 ;
    END
  END cm_mem_ctrl_we
  PIN cm_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END cm_sram0_csb0
  PIN cm_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END cm_sram0_dout0[0]
  PIN cm_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END cm_sram0_dout0[10]
  PIN cm_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END cm_sram0_dout0[11]
  PIN cm_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END cm_sram0_dout0[12]
  PIN cm_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END cm_sram0_dout0[13]
  PIN cm_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END cm_sram0_dout0[14]
  PIN cm_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END cm_sram0_dout0[15]
  PIN cm_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END cm_sram0_dout0[16]
  PIN cm_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END cm_sram0_dout0[17]
  PIN cm_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END cm_sram0_dout0[18]
  PIN cm_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END cm_sram0_dout0[19]
  PIN cm_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END cm_sram0_dout0[1]
  PIN cm_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END cm_sram0_dout0[20]
  PIN cm_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END cm_sram0_dout0[21]
  PIN cm_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END cm_sram0_dout0[22]
  PIN cm_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END cm_sram0_dout0[23]
  PIN cm_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END cm_sram0_dout0[24]
  PIN cm_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END cm_sram0_dout0[25]
  PIN cm_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END cm_sram0_dout0[26]
  PIN cm_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END cm_sram0_dout0[27]
  PIN cm_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END cm_sram0_dout0[28]
  PIN cm_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END cm_sram0_dout0[29]
  PIN cm_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END cm_sram0_dout0[2]
  PIN cm_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END cm_sram0_dout0[30]
  PIN cm_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END cm_sram0_dout0[31]
  PIN cm_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END cm_sram0_dout0[3]
  PIN cm_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END cm_sram0_dout0[4]
  PIN cm_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END cm_sram0_dout0[5]
  PIN cm_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END cm_sram0_dout0[6]
  PIN cm_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END cm_sram0_dout0[7]
  PIN cm_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END cm_sram0_dout0[8]
  PIN cm_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END cm_sram0_dout0[9]
  PIN cm_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END cm_sram0_web0
  PIN cm_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END cm_sram1_csb0
  PIN cm_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END cm_sram1_dout0[0]
  PIN cm_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END cm_sram1_dout0[10]
  PIN cm_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END cm_sram1_dout0[11]
  PIN cm_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END cm_sram1_dout0[12]
  PIN cm_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END cm_sram1_dout0[13]
  PIN cm_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END cm_sram1_dout0[14]
  PIN cm_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END cm_sram1_dout0[15]
  PIN cm_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END cm_sram1_dout0[16]
  PIN cm_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END cm_sram1_dout0[17]
  PIN cm_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END cm_sram1_dout0[18]
  PIN cm_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END cm_sram1_dout0[19]
  PIN cm_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END cm_sram1_dout0[1]
  PIN cm_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END cm_sram1_dout0[20]
  PIN cm_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END cm_sram1_dout0[21]
  PIN cm_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END cm_sram1_dout0[22]
  PIN cm_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END cm_sram1_dout0[23]
  PIN cm_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END cm_sram1_dout0[24]
  PIN cm_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END cm_sram1_dout0[25]
  PIN cm_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END cm_sram1_dout0[26]
  PIN cm_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END cm_sram1_dout0[27]
  PIN cm_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END cm_sram1_dout0[28]
  PIN cm_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END cm_sram1_dout0[29]
  PIN cm_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END cm_sram1_dout0[2]
  PIN cm_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END cm_sram1_dout0[30]
  PIN cm_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END cm_sram1_dout0[31]
  PIN cm_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END cm_sram1_dout0[3]
  PIN cm_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END cm_sram1_dout0[4]
  PIN cm_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END cm_sram1_dout0[5]
  PIN cm_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END cm_sram1_dout0[6]
  PIN cm_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END cm_sram1_dout0[7]
  PIN cm_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END cm_sram1_dout0[8]
  PIN cm_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END cm_sram1_dout0[9]
  PIN cm_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END cm_sram1_web0
  PIN cm_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END cm_sram2_csb0
  PIN cm_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END cm_sram2_dout0[0]
  PIN cm_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END cm_sram2_dout0[10]
  PIN cm_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END cm_sram2_dout0[11]
  PIN cm_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END cm_sram2_dout0[12]
  PIN cm_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END cm_sram2_dout0[13]
  PIN cm_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END cm_sram2_dout0[14]
  PIN cm_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END cm_sram2_dout0[15]
  PIN cm_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END cm_sram2_dout0[16]
  PIN cm_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END cm_sram2_dout0[17]
  PIN cm_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END cm_sram2_dout0[18]
  PIN cm_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END cm_sram2_dout0[19]
  PIN cm_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END cm_sram2_dout0[1]
  PIN cm_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END cm_sram2_dout0[20]
  PIN cm_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END cm_sram2_dout0[21]
  PIN cm_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END cm_sram2_dout0[22]
  PIN cm_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END cm_sram2_dout0[23]
  PIN cm_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END cm_sram2_dout0[24]
  PIN cm_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END cm_sram2_dout0[25]
  PIN cm_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END cm_sram2_dout0[26]
  PIN cm_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END cm_sram2_dout0[27]
  PIN cm_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END cm_sram2_dout0[28]
  PIN cm_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END cm_sram2_dout0[29]
  PIN cm_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END cm_sram2_dout0[2]
  PIN cm_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END cm_sram2_dout0[30]
  PIN cm_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END cm_sram2_dout0[31]
  PIN cm_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END cm_sram2_dout0[3]
  PIN cm_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END cm_sram2_dout0[4]
  PIN cm_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END cm_sram2_dout0[5]
  PIN cm_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END cm_sram2_dout0[6]
  PIN cm_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END cm_sram2_dout0[7]
  PIN cm_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END cm_sram2_dout0[8]
  PIN cm_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END cm_sram2_dout0[9]
  PIN cm_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END cm_sram2_web0
  PIN cm_sram3_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END cm_sram3_csb0
  PIN cm_sram3_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END cm_sram3_dout0[0]
  PIN cm_sram3_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END cm_sram3_dout0[10]
  PIN cm_sram3_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END cm_sram3_dout0[11]
  PIN cm_sram3_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END cm_sram3_dout0[12]
  PIN cm_sram3_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END cm_sram3_dout0[13]
  PIN cm_sram3_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END cm_sram3_dout0[14]
  PIN cm_sram3_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END cm_sram3_dout0[15]
  PIN cm_sram3_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END cm_sram3_dout0[16]
  PIN cm_sram3_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END cm_sram3_dout0[17]
  PIN cm_sram3_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END cm_sram3_dout0[18]
  PIN cm_sram3_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END cm_sram3_dout0[19]
  PIN cm_sram3_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END cm_sram3_dout0[1]
  PIN cm_sram3_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END cm_sram3_dout0[20]
  PIN cm_sram3_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END cm_sram3_dout0[21]
  PIN cm_sram3_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END cm_sram3_dout0[22]
  PIN cm_sram3_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END cm_sram3_dout0[23]
  PIN cm_sram3_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END cm_sram3_dout0[24]
  PIN cm_sram3_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END cm_sram3_dout0[25]
  PIN cm_sram3_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END cm_sram3_dout0[26]
  PIN cm_sram3_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END cm_sram3_dout0[27]
  PIN cm_sram3_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END cm_sram3_dout0[28]
  PIN cm_sram3_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END cm_sram3_dout0[29]
  PIN cm_sram3_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END cm_sram3_dout0[2]
  PIN cm_sram3_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END cm_sram3_dout0[30]
  PIN cm_sram3_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END cm_sram3_dout0[31]
  PIN cm_sram3_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END cm_sram3_dout0[3]
  PIN cm_sram3_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END cm_sram3_dout0[4]
  PIN cm_sram3_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END cm_sram3_dout0[5]
  PIN cm_sram3_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END cm_sram3_dout0[6]
  PIN cm_sram3_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END cm_sram3_dout0[7]
  PIN cm_sram3_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END cm_sram3_dout0[8]
  PIN cm_sram3_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END cm_sram3_dout0[9]
  PIN cm_sram3_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END cm_sram3_web0
  PIN cm_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END cm_sram_comm_addr0[0]
  PIN cm_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END cm_sram_comm_addr0[1]
  PIN cm_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END cm_sram_comm_addr0[2]
  PIN cm_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END cm_sram_comm_addr0[3]
  PIN cm_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END cm_sram_comm_addr0[4]
  PIN cm_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END cm_sram_comm_addr0[5]
  PIN cm_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END cm_sram_comm_addr0[6]
  PIN cm_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END cm_sram_comm_addr0[7]
  PIN cm_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END cm_sram_comm_addr0[8]
  PIN cm_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END cm_sram_comm_din0[0]
  PIN cm_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END cm_sram_comm_din0[10]
  PIN cm_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END cm_sram_comm_din0[11]
  PIN cm_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END cm_sram_comm_din0[12]
  PIN cm_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END cm_sram_comm_din0[13]
  PIN cm_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END cm_sram_comm_din0[14]
  PIN cm_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END cm_sram_comm_din0[15]
  PIN cm_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END cm_sram_comm_din0[16]
  PIN cm_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END cm_sram_comm_din0[17]
  PIN cm_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END cm_sram_comm_din0[18]
  PIN cm_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END cm_sram_comm_din0[19]
  PIN cm_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END cm_sram_comm_din0[1]
  PIN cm_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END cm_sram_comm_din0[20]
  PIN cm_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END cm_sram_comm_din0[21]
  PIN cm_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END cm_sram_comm_din0[22]
  PIN cm_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END cm_sram_comm_din0[23]
  PIN cm_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END cm_sram_comm_din0[24]
  PIN cm_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END cm_sram_comm_din0[25]
  PIN cm_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END cm_sram_comm_din0[26]
  PIN cm_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END cm_sram_comm_din0[27]
  PIN cm_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END cm_sram_comm_din0[28]
  PIN cm_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END cm_sram_comm_din0[29]
  PIN cm_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END cm_sram_comm_din0[2]
  PIN cm_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END cm_sram_comm_din0[30]
  PIN cm_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END cm_sram_comm_din0[31]
  PIN cm_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END cm_sram_comm_din0[3]
  PIN cm_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END cm_sram_comm_din0[4]
  PIN cm_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END cm_sram_comm_din0[5]
  PIN cm_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END cm_sram_comm_din0[6]
  PIN cm_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END cm_sram_comm_din0[7]
  PIN cm_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END cm_sram_comm_din0[8]
  PIN cm_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END cm_sram_comm_din0[9]
  PIN ct_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 223.080 600.000 223.680 ;
    END
  END ct_mem_ctrl_addr[0]
  PIN ct_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 250.960 600.000 251.560 ;
    END
  END ct_mem_ctrl_addr[10]
  PIN ct_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 253.680 600.000 254.280 ;
    END
  END ct_mem_ctrl_addr[11]
  PIN ct_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 256.400 600.000 257.000 ;
    END
  END ct_mem_ctrl_addr[12]
  PIN ct_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 259.120 600.000 259.720 ;
    END
  END ct_mem_ctrl_addr[13]
  PIN ct_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 225.800 600.000 226.400 ;
    END
  END ct_mem_ctrl_addr[1]
  PIN ct_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 228.520 600.000 229.120 ;
    END
  END ct_mem_ctrl_addr[2]
  PIN ct_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 231.240 600.000 231.840 ;
    END
  END ct_mem_ctrl_addr[3]
  PIN ct_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 233.960 600.000 234.560 ;
    END
  END ct_mem_ctrl_addr[4]
  PIN ct_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 236.680 600.000 237.280 ;
    END
  END ct_mem_ctrl_addr[5]
  PIN ct_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 239.400 600.000 240.000 ;
    END
  END ct_mem_ctrl_addr[6]
  PIN ct_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 242.120 600.000 242.720 ;
    END
  END ct_mem_ctrl_addr[7]
  PIN ct_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 244.840 600.000 245.440 ;
    END
  END ct_mem_ctrl_addr[8]
  PIN ct_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 248.240 600.000 248.840 ;
    END
  END ct_mem_ctrl_addr[9]
  PIN ct_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 261.840 600.000 262.440 ;
    END
  END ct_mem_ctrl_in[0]
  PIN ct_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 289.040 600.000 289.640 ;
    END
  END ct_mem_ctrl_in[10]
  PIN ct_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 291.760 600.000 292.360 ;
    END
  END ct_mem_ctrl_in[11]
  PIN ct_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 294.480 600.000 295.080 ;
    END
  END ct_mem_ctrl_in[12]
  PIN ct_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 297.200 600.000 297.800 ;
    END
  END ct_mem_ctrl_in[13]
  PIN ct_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 299.920 600.000 300.520 ;
    END
  END ct_mem_ctrl_in[14]
  PIN ct_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 302.640 600.000 303.240 ;
    END
  END ct_mem_ctrl_in[15]
  PIN ct_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 305.360 600.000 305.960 ;
    END
  END ct_mem_ctrl_in[16]
  PIN ct_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 308.080 600.000 308.680 ;
    END
  END ct_mem_ctrl_in[17]
  PIN ct_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 310.800 600.000 311.400 ;
    END
  END ct_mem_ctrl_in[18]
  PIN ct_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 313.520 600.000 314.120 ;
    END
  END ct_mem_ctrl_in[19]
  PIN ct_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 264.560 600.000 265.160 ;
    END
  END ct_mem_ctrl_in[1]
  PIN ct_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 316.240 600.000 316.840 ;
    END
  END ct_mem_ctrl_in[20]
  PIN ct_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 318.960 600.000 319.560 ;
    END
  END ct_mem_ctrl_in[21]
  PIN ct_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 321.680 600.000 322.280 ;
    END
  END ct_mem_ctrl_in[22]
  PIN ct_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 324.400 600.000 325.000 ;
    END
  END ct_mem_ctrl_in[23]
  PIN ct_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 327.120 600.000 327.720 ;
    END
  END ct_mem_ctrl_in[24]
  PIN ct_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 330.520 600.000 331.120 ;
    END
  END ct_mem_ctrl_in[25]
  PIN ct_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 333.240 600.000 333.840 ;
    END
  END ct_mem_ctrl_in[26]
  PIN ct_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 335.960 600.000 336.560 ;
    END
  END ct_mem_ctrl_in[27]
  PIN ct_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 338.680 600.000 339.280 ;
    END
  END ct_mem_ctrl_in[28]
  PIN ct_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 341.400 600.000 342.000 ;
    END
  END ct_mem_ctrl_in[29]
  PIN ct_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 267.280 600.000 267.880 ;
    END
  END ct_mem_ctrl_in[2]
  PIN ct_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 344.120 600.000 344.720 ;
    END
  END ct_mem_ctrl_in[30]
  PIN ct_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 346.840 600.000 347.440 ;
    END
  END ct_mem_ctrl_in[31]
  PIN ct_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 270.000 600.000 270.600 ;
    END
  END ct_mem_ctrl_in[3]
  PIN ct_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 272.720 600.000 273.320 ;
    END
  END ct_mem_ctrl_in[4]
  PIN ct_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 275.440 600.000 276.040 ;
    END
  END ct_mem_ctrl_in[5]
  PIN ct_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 278.160 600.000 278.760 ;
    END
  END ct_mem_ctrl_in[6]
  PIN ct_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 280.880 600.000 281.480 ;
    END
  END ct_mem_ctrl_in[7]
  PIN ct_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 283.600 600.000 284.200 ;
    END
  END ct_mem_ctrl_in[8]
  PIN ct_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 286.320 600.000 286.920 ;
    END
  END ct_mem_ctrl_in[9]
  PIN ct_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 349.560 600.000 350.160 ;
    END
  END ct_mem_ctrl_out[0]
  PIN ct_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 376.760 600.000 377.360 ;
    END
  END ct_mem_ctrl_out[10]
  PIN ct_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 379.480 600.000 380.080 ;
    END
  END ct_mem_ctrl_out[11]
  PIN ct_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 382.200 600.000 382.800 ;
    END
  END ct_mem_ctrl_out[12]
  PIN ct_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 384.920 600.000 385.520 ;
    END
  END ct_mem_ctrl_out[13]
  PIN ct_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 387.640 600.000 388.240 ;
    END
  END ct_mem_ctrl_out[14]
  PIN ct_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 390.360 600.000 390.960 ;
    END
  END ct_mem_ctrl_out[15]
  PIN ct_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 393.080 600.000 393.680 ;
    END
  END ct_mem_ctrl_out[16]
  PIN ct_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 395.800 600.000 396.400 ;
    END
  END ct_mem_ctrl_out[17]
  PIN ct_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 398.520 600.000 399.120 ;
    END
  END ct_mem_ctrl_out[18]
  PIN ct_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 401.240 600.000 401.840 ;
    END
  END ct_mem_ctrl_out[19]
  PIN ct_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 352.280 600.000 352.880 ;
    END
  END ct_mem_ctrl_out[1]
  PIN ct_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 403.960 600.000 404.560 ;
    END
  END ct_mem_ctrl_out[20]
  PIN ct_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 406.680 600.000 407.280 ;
    END
  END ct_mem_ctrl_out[21]
  PIN ct_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 410.080 600.000 410.680 ;
    END
  END ct_mem_ctrl_out[22]
  PIN ct_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 412.800 600.000 413.400 ;
    END
  END ct_mem_ctrl_out[23]
  PIN ct_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 415.520 600.000 416.120 ;
    END
  END ct_mem_ctrl_out[24]
  PIN ct_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 418.240 600.000 418.840 ;
    END
  END ct_mem_ctrl_out[25]
  PIN ct_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 420.960 600.000 421.560 ;
    END
  END ct_mem_ctrl_out[26]
  PIN ct_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 423.680 600.000 424.280 ;
    END
  END ct_mem_ctrl_out[27]
  PIN ct_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 426.400 600.000 427.000 ;
    END
  END ct_mem_ctrl_out[28]
  PIN ct_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 429.120 600.000 429.720 ;
    END
  END ct_mem_ctrl_out[29]
  PIN ct_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 355.000 600.000 355.600 ;
    END
  END ct_mem_ctrl_out[2]
  PIN ct_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 431.840 600.000 432.440 ;
    END
  END ct_mem_ctrl_out[30]
  PIN ct_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 434.560 600.000 435.160 ;
    END
  END ct_mem_ctrl_out[31]
  PIN ct_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 357.720 600.000 358.320 ;
    END
  END ct_mem_ctrl_out[3]
  PIN ct_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 360.440 600.000 361.040 ;
    END
  END ct_mem_ctrl_out[4]
  PIN ct_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 363.160 600.000 363.760 ;
    END
  END ct_mem_ctrl_out[5]
  PIN ct_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 365.880 600.000 366.480 ;
    END
  END ct_mem_ctrl_out[6]
  PIN ct_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 368.600 600.000 369.200 ;
    END
  END ct_mem_ctrl_out[7]
  PIN ct_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 371.320 600.000 371.920 ;
    END
  END ct_mem_ctrl_out[8]
  PIN ct_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 374.040 600.000 374.640 ;
    END
  END ct_mem_ctrl_out[9]
  PIN ct_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 437.280 600.000 437.880 ;
    END
  END ct_mem_ctrl_req
  PIN ct_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 440.000 600.000 440.600 ;
    END
  END ct_mem_ctrl_vld
  PIN ct_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 442.720 600.000 443.320 ;
    END
  END ct_mem_ctrl_we
  PIN ct_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END ct_sram0_csb0
  PIN ct_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END ct_sram0_dout0[0]
  PIN ct_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END ct_sram0_dout0[10]
  PIN ct_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END ct_sram0_dout0[11]
  PIN ct_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END ct_sram0_dout0[12]
  PIN ct_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END ct_sram0_dout0[13]
  PIN ct_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END ct_sram0_dout0[14]
  PIN ct_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END ct_sram0_dout0[15]
  PIN ct_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END ct_sram0_dout0[16]
  PIN ct_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END ct_sram0_dout0[17]
  PIN ct_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END ct_sram0_dout0[18]
  PIN ct_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END ct_sram0_dout0[19]
  PIN ct_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END ct_sram0_dout0[1]
  PIN ct_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END ct_sram0_dout0[20]
  PIN ct_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END ct_sram0_dout0[21]
  PIN ct_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END ct_sram0_dout0[22]
  PIN ct_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END ct_sram0_dout0[23]
  PIN ct_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END ct_sram0_dout0[24]
  PIN ct_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END ct_sram0_dout0[25]
  PIN ct_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END ct_sram0_dout0[26]
  PIN ct_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END ct_sram0_dout0[27]
  PIN ct_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END ct_sram0_dout0[28]
  PIN ct_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END ct_sram0_dout0[29]
  PIN ct_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END ct_sram0_dout0[2]
  PIN ct_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END ct_sram0_dout0[30]
  PIN ct_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END ct_sram0_dout0[31]
  PIN ct_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END ct_sram0_dout0[3]
  PIN ct_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END ct_sram0_dout0[4]
  PIN ct_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END ct_sram0_dout0[5]
  PIN ct_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END ct_sram0_dout0[6]
  PIN ct_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END ct_sram0_dout0[7]
  PIN ct_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END ct_sram0_dout0[8]
  PIN ct_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END ct_sram0_dout0[9]
  PIN ct_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END ct_sram0_web0
  PIN ct_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END ct_sram1_csb0
  PIN ct_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END ct_sram1_dout0[0]
  PIN ct_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END ct_sram1_dout0[10]
  PIN ct_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END ct_sram1_dout0[11]
  PIN ct_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END ct_sram1_dout0[12]
  PIN ct_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END ct_sram1_dout0[13]
  PIN ct_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END ct_sram1_dout0[14]
  PIN ct_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END ct_sram1_dout0[15]
  PIN ct_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END ct_sram1_dout0[16]
  PIN ct_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END ct_sram1_dout0[17]
  PIN ct_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END ct_sram1_dout0[18]
  PIN ct_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END ct_sram1_dout0[19]
  PIN ct_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END ct_sram1_dout0[1]
  PIN ct_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END ct_sram1_dout0[20]
  PIN ct_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END ct_sram1_dout0[21]
  PIN ct_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END ct_sram1_dout0[22]
  PIN ct_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END ct_sram1_dout0[23]
  PIN ct_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END ct_sram1_dout0[24]
  PIN ct_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END ct_sram1_dout0[25]
  PIN ct_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END ct_sram1_dout0[26]
  PIN ct_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END ct_sram1_dout0[27]
  PIN ct_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END ct_sram1_dout0[28]
  PIN ct_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END ct_sram1_dout0[29]
  PIN ct_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END ct_sram1_dout0[2]
  PIN ct_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END ct_sram1_dout0[30]
  PIN ct_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END ct_sram1_dout0[31]
  PIN ct_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END ct_sram1_dout0[3]
  PIN ct_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END ct_sram1_dout0[4]
  PIN ct_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END ct_sram1_dout0[5]
  PIN ct_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END ct_sram1_dout0[6]
  PIN ct_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END ct_sram1_dout0[7]
  PIN ct_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END ct_sram1_dout0[8]
  PIN ct_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END ct_sram1_dout0[9]
  PIN ct_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END ct_sram1_web0
  PIN ct_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END ct_sram2_csb0
  PIN ct_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END ct_sram2_dout0[0]
  PIN ct_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END ct_sram2_dout0[10]
  PIN ct_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END ct_sram2_dout0[11]
  PIN ct_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END ct_sram2_dout0[12]
  PIN ct_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END ct_sram2_dout0[13]
  PIN ct_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END ct_sram2_dout0[14]
  PIN ct_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END ct_sram2_dout0[15]
  PIN ct_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END ct_sram2_dout0[16]
  PIN ct_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END ct_sram2_dout0[17]
  PIN ct_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END ct_sram2_dout0[18]
  PIN ct_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END ct_sram2_dout0[19]
  PIN ct_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END ct_sram2_dout0[1]
  PIN ct_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END ct_sram2_dout0[20]
  PIN ct_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END ct_sram2_dout0[21]
  PIN ct_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END ct_sram2_dout0[22]
  PIN ct_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END ct_sram2_dout0[23]
  PIN ct_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END ct_sram2_dout0[24]
  PIN ct_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END ct_sram2_dout0[25]
  PIN ct_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END ct_sram2_dout0[26]
  PIN ct_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END ct_sram2_dout0[27]
  PIN ct_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END ct_sram2_dout0[28]
  PIN ct_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END ct_sram2_dout0[29]
  PIN ct_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END ct_sram2_dout0[2]
  PIN ct_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END ct_sram2_dout0[30]
  PIN ct_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END ct_sram2_dout0[31]
  PIN ct_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END ct_sram2_dout0[3]
  PIN ct_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END ct_sram2_dout0[4]
  PIN ct_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END ct_sram2_dout0[5]
  PIN ct_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END ct_sram2_dout0[6]
  PIN ct_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END ct_sram2_dout0[7]
  PIN ct_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END ct_sram2_dout0[8]
  PIN ct_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END ct_sram2_dout0[9]
  PIN ct_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END ct_sram2_web0
  PIN ct_sram3_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END ct_sram3_csb0
  PIN ct_sram3_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END ct_sram3_dout0[0]
  PIN ct_sram3_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END ct_sram3_dout0[10]
  PIN ct_sram3_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END ct_sram3_dout0[11]
  PIN ct_sram3_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END ct_sram3_dout0[12]
  PIN ct_sram3_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END ct_sram3_dout0[13]
  PIN ct_sram3_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END ct_sram3_dout0[14]
  PIN ct_sram3_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END ct_sram3_dout0[15]
  PIN ct_sram3_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END ct_sram3_dout0[16]
  PIN ct_sram3_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END ct_sram3_dout0[17]
  PIN ct_sram3_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END ct_sram3_dout0[18]
  PIN ct_sram3_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END ct_sram3_dout0[19]
  PIN ct_sram3_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END ct_sram3_dout0[1]
  PIN ct_sram3_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END ct_sram3_dout0[20]
  PIN ct_sram3_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END ct_sram3_dout0[21]
  PIN ct_sram3_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END ct_sram3_dout0[22]
  PIN ct_sram3_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END ct_sram3_dout0[23]
  PIN ct_sram3_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END ct_sram3_dout0[24]
  PIN ct_sram3_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END ct_sram3_dout0[25]
  PIN ct_sram3_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END ct_sram3_dout0[26]
  PIN ct_sram3_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END ct_sram3_dout0[27]
  PIN ct_sram3_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END ct_sram3_dout0[28]
  PIN ct_sram3_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END ct_sram3_dout0[29]
  PIN ct_sram3_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END ct_sram3_dout0[2]
  PIN ct_sram3_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END ct_sram3_dout0[30]
  PIN ct_sram3_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END ct_sram3_dout0[31]
  PIN ct_sram3_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END ct_sram3_dout0[3]
  PIN ct_sram3_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END ct_sram3_dout0[4]
  PIN ct_sram3_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END ct_sram3_dout0[5]
  PIN ct_sram3_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END ct_sram3_dout0[6]
  PIN ct_sram3_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END ct_sram3_dout0[7]
  PIN ct_sram3_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END ct_sram3_dout0[8]
  PIN ct_sram3_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END ct_sram3_dout0[9]
  PIN ct_sram3_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END ct_sram3_web0
  PIN ct_sram4_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END ct_sram4_csb0
  PIN ct_sram4_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END ct_sram4_dout0[0]
  PIN ct_sram4_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END ct_sram4_dout0[10]
  PIN ct_sram4_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END ct_sram4_dout0[11]
  PIN ct_sram4_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END ct_sram4_dout0[12]
  PIN ct_sram4_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END ct_sram4_dout0[13]
  PIN ct_sram4_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END ct_sram4_dout0[14]
  PIN ct_sram4_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END ct_sram4_dout0[15]
  PIN ct_sram4_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END ct_sram4_dout0[16]
  PIN ct_sram4_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END ct_sram4_dout0[17]
  PIN ct_sram4_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 0.000 516.950 4.000 ;
    END
  END ct_sram4_dout0[18]
  PIN ct_sram4_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END ct_sram4_dout0[19]
  PIN ct_sram4_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END ct_sram4_dout0[1]
  PIN ct_sram4_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END ct_sram4_dout0[20]
  PIN ct_sram4_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END ct_sram4_dout0[21]
  PIN ct_sram4_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END ct_sram4_dout0[22]
  PIN ct_sram4_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END ct_sram4_dout0[23]
  PIN ct_sram4_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END ct_sram4_dout0[24]
  PIN ct_sram4_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END ct_sram4_dout0[25]
  PIN ct_sram4_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END ct_sram4_dout0[26]
  PIN ct_sram4_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END ct_sram4_dout0[27]
  PIN ct_sram4_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END ct_sram4_dout0[28]
  PIN ct_sram4_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END ct_sram4_dout0[29]
  PIN ct_sram4_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END ct_sram4_dout0[2]
  PIN ct_sram4_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END ct_sram4_dout0[30]
  PIN ct_sram4_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END ct_sram4_dout0[31]
  PIN ct_sram4_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END ct_sram4_dout0[3]
  PIN ct_sram4_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END ct_sram4_dout0[4]
  PIN ct_sram4_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END ct_sram4_dout0[5]
  PIN ct_sram4_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END ct_sram4_dout0[6]
  PIN ct_sram4_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END ct_sram4_dout0[7]
  PIN ct_sram4_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END ct_sram4_dout0[8]
  PIN ct_sram4_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END ct_sram4_dout0[9]
  PIN ct_sram4_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END ct_sram4_web0
  PIN ct_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END ct_sram_comm_addr0[0]
  PIN ct_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END ct_sram_comm_addr0[1]
  PIN ct_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END ct_sram_comm_addr0[2]
  PIN ct_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END ct_sram_comm_addr0[3]
  PIN ct_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END ct_sram_comm_addr0[4]
  PIN ct_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END ct_sram_comm_addr0[5]
  PIN ct_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END ct_sram_comm_addr0[6]
  PIN ct_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END ct_sram_comm_addr0[7]
  PIN ct_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END ct_sram_comm_addr0[8]
  PIN ct_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END ct_sram_comm_din0[0]
  PIN ct_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END ct_sram_comm_din0[10]
  PIN ct_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END ct_sram_comm_din0[11]
  PIN ct_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END ct_sram_comm_din0[12]
  PIN ct_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END ct_sram_comm_din0[13]
  PIN ct_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END ct_sram_comm_din0[14]
  PIN ct_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END ct_sram_comm_din0[15]
  PIN ct_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END ct_sram_comm_din0[16]
  PIN ct_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END ct_sram_comm_din0[17]
  PIN ct_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END ct_sram_comm_din0[18]
  PIN ct_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END ct_sram_comm_din0[19]
  PIN ct_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END ct_sram_comm_din0[1]
  PIN ct_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END ct_sram_comm_din0[20]
  PIN ct_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END ct_sram_comm_din0[21]
  PIN ct_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END ct_sram_comm_din0[22]
  PIN ct_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END ct_sram_comm_din0[23]
  PIN ct_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END ct_sram_comm_din0[24]
  PIN ct_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END ct_sram_comm_din0[25]
  PIN ct_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END ct_sram_comm_din0[26]
  PIN ct_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END ct_sram_comm_din0[27]
  PIN ct_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END ct_sram_comm_din0[28]
  PIN ct_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END ct_sram_comm_din0[29]
  PIN ct_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END ct_sram_comm_din0[2]
  PIN ct_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 0.000 597.450 4.000 ;
    END
  END ct_sram_comm_din0[30]
  PIN ct_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END ct_sram_comm_din0[31]
  PIN ct_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END ct_sram_comm_din0[3]
  PIN ct_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END ct_sram_comm_din0[4]
  PIN ct_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END ct_sram_comm_din0[5]
  PIN ct_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END ct_sram_comm_din0[6]
  PIN ct_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END ct_sram_comm_din0[7]
  PIN ct_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END ct_sram_comm_din0[8]
  PIN ct_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END ct_sram_comm_din0[9]
  PIN main_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END main_mem_addr[0]
  PIN main_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END main_mem_addr[1]
  PIN main_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END main_mem_addr[2]
  PIN main_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END main_mem_addr[3]
  PIN main_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END main_mem_addr[4]
  PIN main_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END main_mem_addr[5]
  PIN main_mem_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END main_mem_in[0]
  PIN main_mem_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END main_mem_in[10]
  PIN main_mem_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END main_mem_in[11]
  PIN main_mem_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END main_mem_in[12]
  PIN main_mem_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END main_mem_in[13]
  PIN main_mem_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END main_mem_in[14]
  PIN main_mem_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END main_mem_in[15]
  PIN main_mem_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END main_mem_in[16]
  PIN main_mem_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END main_mem_in[17]
  PIN main_mem_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END main_mem_in[18]
  PIN main_mem_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END main_mem_in[19]
  PIN main_mem_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END main_mem_in[1]
  PIN main_mem_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END main_mem_in[20]
  PIN main_mem_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END main_mem_in[21]
  PIN main_mem_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END main_mem_in[22]
  PIN main_mem_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END main_mem_in[23]
  PIN main_mem_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END main_mem_in[24]
  PIN main_mem_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END main_mem_in[25]
  PIN main_mem_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END main_mem_in[26]
  PIN main_mem_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END main_mem_in[27]
  PIN main_mem_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END main_mem_in[28]
  PIN main_mem_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END main_mem_in[29]
  PIN main_mem_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END main_mem_in[2]
  PIN main_mem_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END main_mem_in[30]
  PIN main_mem_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END main_mem_in[31]
  PIN main_mem_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END main_mem_in[3]
  PIN main_mem_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END main_mem_in[4]
  PIN main_mem_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END main_mem_in[5]
  PIN main_mem_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END main_mem_in[6]
  PIN main_mem_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END main_mem_in[7]
  PIN main_mem_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END main_mem_in[8]
  PIN main_mem_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END main_mem_in[9]
  PIN main_mem_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END main_mem_out[0]
  PIN main_mem_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END main_mem_out[10]
  PIN main_mem_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END main_mem_out[11]
  PIN main_mem_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END main_mem_out[12]
  PIN main_mem_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END main_mem_out[13]
  PIN main_mem_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END main_mem_out[14]
  PIN main_mem_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END main_mem_out[15]
  PIN main_mem_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END main_mem_out[16]
  PIN main_mem_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END main_mem_out[17]
  PIN main_mem_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END main_mem_out[18]
  PIN main_mem_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END main_mem_out[19]
  PIN main_mem_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END main_mem_out[1]
  PIN main_mem_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END main_mem_out[20]
  PIN main_mem_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END main_mem_out[21]
  PIN main_mem_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END main_mem_out[22]
  PIN main_mem_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END main_mem_out[23]
  PIN main_mem_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END main_mem_out[24]
  PIN main_mem_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END main_mem_out[25]
  PIN main_mem_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END main_mem_out[26]
  PIN main_mem_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END main_mem_out[27]
  PIN main_mem_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END main_mem_out[28]
  PIN main_mem_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END main_mem_out[29]
  PIN main_mem_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END main_mem_out[2]
  PIN main_mem_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END main_mem_out[30]
  PIN main_mem_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END main_mem_out[31]
  PIN main_mem_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END main_mem_out[3]
  PIN main_mem_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END main_mem_out[4]
  PIN main_mem_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END main_mem_out[5]
  PIN main_mem_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END main_mem_out[6]
  PIN main_mem_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END main_mem_out[7]
  PIN main_mem_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END main_mem_out[8]
  PIN main_mem_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END main_mem_out[9]
  PIN main_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END main_mem_we
  PIN program_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 673.240 600.000 673.840 ;
    END
  END program_sel[0]
  PIN program_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 675.960 600.000 676.560 ;
    END
  END program_sel[1]
  PIN r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 714.040 600.000 714.640 ;
    END
  END r_data[0]
  PIN r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 716.760 600.000 717.360 ;
    END
  END r_data[1]
  PIN r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 719.480 600.000 720.080 ;
    END
  END r_data[2]
  PIN r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 722.200 600.000 722.800 ;
    END
  END r_data[3]
  PIN r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 724.920 600.000 725.520 ;
    END
  END r_data[4]
  PIN r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 727.640 600.000 728.240 ;
    END
  END r_data[5]
  PIN r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 730.360 600.000 730.960 ;
    END
  END r_data[6]
  PIN r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 733.080 600.000 733.680 ;
    END
  END r_data[7]
  PIN rd_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 681.400 600.000 682.000 ;
    END
  END rd_uart
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 667.800 600.000 668.400 ;
    END
  END rst
  PIN rst_asserted
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 670.520 600.000 671.120 ;
    END
  END rst_asserted
  PIN rx_empty
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 711.320 600.000 711.920 ;
    END
  END rx_empty
  PIN rx_fifo_flush_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 678.680 600.000 679.280 ;
    END
  END rx_fifo_flush_enable
  PIN sram_const_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END sram_const_addr1[0]
  PIN sram_const_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END sram_const_addr1[1]
  PIN sram_const_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END sram_const_addr1[2]
  PIN sram_const_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END sram_const_addr1[3]
  PIN sram_const_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END sram_const_addr1[4]
  PIN sram_const_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END sram_const_addr1[5]
  PIN sram_const_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END sram_const_addr1[6]
  PIN sram_const_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END sram_const_addr1[7]
  PIN sram_const_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END sram_const_addr1[8]
  PIN sram_const_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END sram_const_csb1
  PIN sram_const_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END sram_const_wmask0[0]
  PIN sram_const_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END sram_const_wmask0[1]
  PIN sram_const_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END sram_const_wmask0[2]
  PIN sram_const_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END sram_const_wmask0[3]
  PIN tx_full
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 708.600 600.000 709.200 ;
    END
  END tx_full
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 723.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 723.760 ;
    END
  END vssd1
  PIN w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 686.840 600.000 687.440 ;
    END
  END w_data[0]
  PIN w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 689.560 600.000 690.160 ;
    END
  END w_data[1]
  PIN w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 692.280 600.000 692.880 ;
    END
  END w_data[2]
  PIN w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 695.000 600.000 695.600 ;
    END
  END w_data[3]
  PIN w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 697.720 600.000 698.320 ;
    END
  END w_data[4]
  PIN w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 700.440 600.000 701.040 ;
    END
  END w_data[5]
  PIN w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 703.160 600.000 703.760 ;
    END
  END w_data[6]
  PIN w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 705.880 600.000 706.480 ;
    END
  END w_data[7]
  PIN wr_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 684.120 600.000 684.720 ;
    END
  END wr_uart
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 723.605 ;
      LAYER met1 ;
        RECT 0.530 1.740 599.770 723.760 ;
      LAYER met2 ;
        RECT 0.560 4.280 599.740 733.565 ;
        RECT 1.110 1.515 1.650 4.280 ;
        RECT 2.490 1.515 3.030 4.280 ;
        RECT 3.870 1.515 4.410 4.280 ;
        RECT 5.250 1.515 5.790 4.280 ;
        RECT 6.630 1.515 7.630 4.280 ;
        RECT 8.470 1.515 9.010 4.280 ;
        RECT 9.850 1.515 10.390 4.280 ;
        RECT 11.230 1.515 11.770 4.280 ;
        RECT 12.610 1.515 13.610 4.280 ;
        RECT 14.450 1.515 14.990 4.280 ;
        RECT 15.830 1.515 16.370 4.280 ;
        RECT 17.210 1.515 17.750 4.280 ;
        RECT 18.590 1.515 19.590 4.280 ;
        RECT 20.430 1.515 20.970 4.280 ;
        RECT 21.810 1.515 22.350 4.280 ;
        RECT 23.190 1.515 23.730 4.280 ;
        RECT 24.570 1.515 25.570 4.280 ;
        RECT 26.410 1.515 26.950 4.280 ;
        RECT 27.790 1.515 28.330 4.280 ;
        RECT 29.170 1.515 29.710 4.280 ;
        RECT 30.550 1.515 31.550 4.280 ;
        RECT 32.390 1.515 32.930 4.280 ;
        RECT 33.770 1.515 34.310 4.280 ;
        RECT 35.150 1.515 35.690 4.280 ;
        RECT 36.530 1.515 37.530 4.280 ;
        RECT 38.370 1.515 38.910 4.280 ;
        RECT 39.750 1.515 40.290 4.280 ;
        RECT 41.130 1.515 41.670 4.280 ;
        RECT 42.510 1.515 43.510 4.280 ;
        RECT 44.350 1.515 44.890 4.280 ;
        RECT 45.730 1.515 46.270 4.280 ;
        RECT 47.110 1.515 47.650 4.280 ;
        RECT 48.490 1.515 49.490 4.280 ;
        RECT 50.330 1.515 50.870 4.280 ;
        RECT 51.710 1.515 52.250 4.280 ;
        RECT 53.090 1.515 53.630 4.280 ;
        RECT 54.470 1.515 55.470 4.280 ;
        RECT 56.310 1.515 56.850 4.280 ;
        RECT 57.690 1.515 58.230 4.280 ;
        RECT 59.070 1.515 59.610 4.280 ;
        RECT 60.450 1.515 60.990 4.280 ;
        RECT 61.830 1.515 62.830 4.280 ;
        RECT 63.670 1.515 64.210 4.280 ;
        RECT 65.050 1.515 65.590 4.280 ;
        RECT 66.430 1.515 66.970 4.280 ;
        RECT 67.810 1.515 68.810 4.280 ;
        RECT 69.650 1.515 70.190 4.280 ;
        RECT 71.030 1.515 71.570 4.280 ;
        RECT 72.410 1.515 72.950 4.280 ;
        RECT 73.790 1.515 74.790 4.280 ;
        RECT 75.630 1.515 76.170 4.280 ;
        RECT 77.010 1.515 77.550 4.280 ;
        RECT 78.390 1.515 78.930 4.280 ;
        RECT 79.770 1.515 80.770 4.280 ;
        RECT 81.610 1.515 82.150 4.280 ;
        RECT 82.990 1.515 83.530 4.280 ;
        RECT 84.370 1.515 84.910 4.280 ;
        RECT 85.750 1.515 86.750 4.280 ;
        RECT 87.590 1.515 88.130 4.280 ;
        RECT 88.970 1.515 89.510 4.280 ;
        RECT 90.350 1.515 90.890 4.280 ;
        RECT 91.730 1.515 92.730 4.280 ;
        RECT 93.570 1.515 94.110 4.280 ;
        RECT 94.950 1.515 95.490 4.280 ;
        RECT 96.330 1.515 96.870 4.280 ;
        RECT 97.710 1.515 98.710 4.280 ;
        RECT 99.550 1.515 100.090 4.280 ;
        RECT 100.930 1.515 101.470 4.280 ;
        RECT 102.310 1.515 102.850 4.280 ;
        RECT 103.690 1.515 104.690 4.280 ;
        RECT 105.530 1.515 106.070 4.280 ;
        RECT 106.910 1.515 107.450 4.280 ;
        RECT 108.290 1.515 108.830 4.280 ;
        RECT 109.670 1.515 110.670 4.280 ;
        RECT 111.510 1.515 112.050 4.280 ;
        RECT 112.890 1.515 113.430 4.280 ;
        RECT 114.270 1.515 114.810 4.280 ;
        RECT 115.650 1.515 116.650 4.280 ;
        RECT 117.490 1.515 118.030 4.280 ;
        RECT 118.870 1.515 119.410 4.280 ;
        RECT 120.250 1.515 120.790 4.280 ;
        RECT 121.630 1.515 122.170 4.280 ;
        RECT 123.010 1.515 124.010 4.280 ;
        RECT 124.850 1.515 125.390 4.280 ;
        RECT 126.230 1.515 126.770 4.280 ;
        RECT 127.610 1.515 128.150 4.280 ;
        RECT 128.990 1.515 129.990 4.280 ;
        RECT 130.830 1.515 131.370 4.280 ;
        RECT 132.210 1.515 132.750 4.280 ;
        RECT 133.590 1.515 134.130 4.280 ;
        RECT 134.970 1.515 135.970 4.280 ;
        RECT 136.810 1.515 137.350 4.280 ;
        RECT 138.190 1.515 138.730 4.280 ;
        RECT 139.570 1.515 140.110 4.280 ;
        RECT 140.950 1.515 141.950 4.280 ;
        RECT 142.790 1.515 143.330 4.280 ;
        RECT 144.170 1.515 144.710 4.280 ;
        RECT 145.550 1.515 146.090 4.280 ;
        RECT 146.930 1.515 147.930 4.280 ;
        RECT 148.770 1.515 149.310 4.280 ;
        RECT 150.150 1.515 150.690 4.280 ;
        RECT 151.530 1.515 152.070 4.280 ;
        RECT 152.910 1.515 153.910 4.280 ;
        RECT 154.750 1.515 155.290 4.280 ;
        RECT 156.130 1.515 156.670 4.280 ;
        RECT 157.510 1.515 158.050 4.280 ;
        RECT 158.890 1.515 159.890 4.280 ;
        RECT 160.730 1.515 161.270 4.280 ;
        RECT 162.110 1.515 162.650 4.280 ;
        RECT 163.490 1.515 164.030 4.280 ;
        RECT 164.870 1.515 165.870 4.280 ;
        RECT 166.710 1.515 167.250 4.280 ;
        RECT 168.090 1.515 168.630 4.280 ;
        RECT 169.470 1.515 170.010 4.280 ;
        RECT 170.850 1.515 171.850 4.280 ;
        RECT 172.690 1.515 173.230 4.280 ;
        RECT 174.070 1.515 174.610 4.280 ;
        RECT 175.450 1.515 175.990 4.280 ;
        RECT 176.830 1.515 177.830 4.280 ;
        RECT 178.670 1.515 179.210 4.280 ;
        RECT 180.050 1.515 180.590 4.280 ;
        RECT 181.430 1.515 181.970 4.280 ;
        RECT 182.810 1.515 183.350 4.280 ;
        RECT 184.190 1.515 185.190 4.280 ;
        RECT 186.030 1.515 186.570 4.280 ;
        RECT 187.410 1.515 187.950 4.280 ;
        RECT 188.790 1.515 189.330 4.280 ;
        RECT 190.170 1.515 191.170 4.280 ;
        RECT 192.010 1.515 192.550 4.280 ;
        RECT 193.390 1.515 193.930 4.280 ;
        RECT 194.770 1.515 195.310 4.280 ;
        RECT 196.150 1.515 197.150 4.280 ;
        RECT 197.990 1.515 198.530 4.280 ;
        RECT 199.370 1.515 199.910 4.280 ;
        RECT 200.750 1.515 201.290 4.280 ;
        RECT 202.130 1.515 203.130 4.280 ;
        RECT 203.970 1.515 204.510 4.280 ;
        RECT 205.350 1.515 205.890 4.280 ;
        RECT 206.730 1.515 207.270 4.280 ;
        RECT 208.110 1.515 209.110 4.280 ;
        RECT 209.950 1.515 210.490 4.280 ;
        RECT 211.330 1.515 211.870 4.280 ;
        RECT 212.710 1.515 213.250 4.280 ;
        RECT 214.090 1.515 215.090 4.280 ;
        RECT 215.930 1.515 216.470 4.280 ;
        RECT 217.310 1.515 217.850 4.280 ;
        RECT 218.690 1.515 219.230 4.280 ;
        RECT 220.070 1.515 221.070 4.280 ;
        RECT 221.910 1.515 222.450 4.280 ;
        RECT 223.290 1.515 223.830 4.280 ;
        RECT 224.670 1.515 225.210 4.280 ;
        RECT 226.050 1.515 227.050 4.280 ;
        RECT 227.890 1.515 228.430 4.280 ;
        RECT 229.270 1.515 229.810 4.280 ;
        RECT 230.650 1.515 231.190 4.280 ;
        RECT 232.030 1.515 233.030 4.280 ;
        RECT 233.870 1.515 234.410 4.280 ;
        RECT 235.250 1.515 235.790 4.280 ;
        RECT 236.630 1.515 237.170 4.280 ;
        RECT 238.010 1.515 239.010 4.280 ;
        RECT 239.850 1.515 240.390 4.280 ;
        RECT 241.230 1.515 241.770 4.280 ;
        RECT 242.610 1.515 243.150 4.280 ;
        RECT 243.990 1.515 244.530 4.280 ;
        RECT 245.370 1.515 246.370 4.280 ;
        RECT 247.210 1.515 247.750 4.280 ;
        RECT 248.590 1.515 249.130 4.280 ;
        RECT 249.970 1.515 250.510 4.280 ;
        RECT 251.350 1.515 252.350 4.280 ;
        RECT 253.190 1.515 253.730 4.280 ;
        RECT 254.570 1.515 255.110 4.280 ;
        RECT 255.950 1.515 256.490 4.280 ;
        RECT 257.330 1.515 258.330 4.280 ;
        RECT 259.170 1.515 259.710 4.280 ;
        RECT 260.550 1.515 261.090 4.280 ;
        RECT 261.930 1.515 262.470 4.280 ;
        RECT 263.310 1.515 264.310 4.280 ;
        RECT 265.150 1.515 265.690 4.280 ;
        RECT 266.530 1.515 267.070 4.280 ;
        RECT 267.910 1.515 268.450 4.280 ;
        RECT 269.290 1.515 270.290 4.280 ;
        RECT 271.130 1.515 271.670 4.280 ;
        RECT 272.510 1.515 273.050 4.280 ;
        RECT 273.890 1.515 274.430 4.280 ;
        RECT 275.270 1.515 276.270 4.280 ;
        RECT 277.110 1.515 277.650 4.280 ;
        RECT 278.490 1.515 279.030 4.280 ;
        RECT 279.870 1.515 280.410 4.280 ;
        RECT 281.250 1.515 282.250 4.280 ;
        RECT 283.090 1.515 283.630 4.280 ;
        RECT 284.470 1.515 285.010 4.280 ;
        RECT 285.850 1.515 286.390 4.280 ;
        RECT 287.230 1.515 288.230 4.280 ;
        RECT 289.070 1.515 289.610 4.280 ;
        RECT 290.450 1.515 290.990 4.280 ;
        RECT 291.830 1.515 292.370 4.280 ;
        RECT 293.210 1.515 294.210 4.280 ;
        RECT 295.050 1.515 295.590 4.280 ;
        RECT 296.430 1.515 296.970 4.280 ;
        RECT 297.810 1.515 298.350 4.280 ;
        RECT 299.190 1.515 300.190 4.280 ;
        RECT 301.030 1.515 301.570 4.280 ;
        RECT 302.410 1.515 302.950 4.280 ;
        RECT 303.790 1.515 304.330 4.280 ;
        RECT 305.170 1.515 305.710 4.280 ;
        RECT 306.550 1.515 307.550 4.280 ;
        RECT 308.390 1.515 308.930 4.280 ;
        RECT 309.770 1.515 310.310 4.280 ;
        RECT 311.150 1.515 311.690 4.280 ;
        RECT 312.530 1.515 313.530 4.280 ;
        RECT 314.370 1.515 314.910 4.280 ;
        RECT 315.750 1.515 316.290 4.280 ;
        RECT 317.130 1.515 317.670 4.280 ;
        RECT 318.510 1.515 319.510 4.280 ;
        RECT 320.350 1.515 320.890 4.280 ;
        RECT 321.730 1.515 322.270 4.280 ;
        RECT 323.110 1.515 323.650 4.280 ;
        RECT 324.490 1.515 325.490 4.280 ;
        RECT 326.330 1.515 326.870 4.280 ;
        RECT 327.710 1.515 328.250 4.280 ;
        RECT 329.090 1.515 329.630 4.280 ;
        RECT 330.470 1.515 331.470 4.280 ;
        RECT 332.310 1.515 332.850 4.280 ;
        RECT 333.690 1.515 334.230 4.280 ;
        RECT 335.070 1.515 335.610 4.280 ;
        RECT 336.450 1.515 337.450 4.280 ;
        RECT 338.290 1.515 338.830 4.280 ;
        RECT 339.670 1.515 340.210 4.280 ;
        RECT 341.050 1.515 341.590 4.280 ;
        RECT 342.430 1.515 343.430 4.280 ;
        RECT 344.270 1.515 344.810 4.280 ;
        RECT 345.650 1.515 346.190 4.280 ;
        RECT 347.030 1.515 347.570 4.280 ;
        RECT 348.410 1.515 349.410 4.280 ;
        RECT 350.250 1.515 350.790 4.280 ;
        RECT 351.630 1.515 352.170 4.280 ;
        RECT 353.010 1.515 353.550 4.280 ;
        RECT 354.390 1.515 355.390 4.280 ;
        RECT 356.230 1.515 356.770 4.280 ;
        RECT 357.610 1.515 358.150 4.280 ;
        RECT 358.990 1.515 359.530 4.280 ;
        RECT 360.370 1.515 360.910 4.280 ;
        RECT 361.750 1.515 362.750 4.280 ;
        RECT 363.590 1.515 364.130 4.280 ;
        RECT 364.970 1.515 365.510 4.280 ;
        RECT 366.350 1.515 366.890 4.280 ;
        RECT 367.730 1.515 368.730 4.280 ;
        RECT 369.570 1.515 370.110 4.280 ;
        RECT 370.950 1.515 371.490 4.280 ;
        RECT 372.330 1.515 372.870 4.280 ;
        RECT 373.710 1.515 374.710 4.280 ;
        RECT 375.550 1.515 376.090 4.280 ;
        RECT 376.930 1.515 377.470 4.280 ;
        RECT 378.310 1.515 378.850 4.280 ;
        RECT 379.690 1.515 380.690 4.280 ;
        RECT 381.530 1.515 382.070 4.280 ;
        RECT 382.910 1.515 383.450 4.280 ;
        RECT 384.290 1.515 384.830 4.280 ;
        RECT 385.670 1.515 386.670 4.280 ;
        RECT 387.510 1.515 388.050 4.280 ;
        RECT 388.890 1.515 389.430 4.280 ;
        RECT 390.270 1.515 390.810 4.280 ;
        RECT 391.650 1.515 392.650 4.280 ;
        RECT 393.490 1.515 394.030 4.280 ;
        RECT 394.870 1.515 395.410 4.280 ;
        RECT 396.250 1.515 396.790 4.280 ;
        RECT 397.630 1.515 398.630 4.280 ;
        RECT 399.470 1.515 400.010 4.280 ;
        RECT 400.850 1.515 401.390 4.280 ;
        RECT 402.230 1.515 402.770 4.280 ;
        RECT 403.610 1.515 404.610 4.280 ;
        RECT 405.450 1.515 405.990 4.280 ;
        RECT 406.830 1.515 407.370 4.280 ;
        RECT 408.210 1.515 408.750 4.280 ;
        RECT 409.590 1.515 410.590 4.280 ;
        RECT 411.430 1.515 411.970 4.280 ;
        RECT 412.810 1.515 413.350 4.280 ;
        RECT 414.190 1.515 414.730 4.280 ;
        RECT 415.570 1.515 416.570 4.280 ;
        RECT 417.410 1.515 417.950 4.280 ;
        RECT 418.790 1.515 419.330 4.280 ;
        RECT 420.170 1.515 420.710 4.280 ;
        RECT 421.550 1.515 422.090 4.280 ;
        RECT 422.930 1.515 423.930 4.280 ;
        RECT 424.770 1.515 425.310 4.280 ;
        RECT 426.150 1.515 426.690 4.280 ;
        RECT 427.530 1.515 428.070 4.280 ;
        RECT 428.910 1.515 429.910 4.280 ;
        RECT 430.750 1.515 431.290 4.280 ;
        RECT 432.130 1.515 432.670 4.280 ;
        RECT 433.510 1.515 434.050 4.280 ;
        RECT 434.890 1.515 435.890 4.280 ;
        RECT 436.730 1.515 437.270 4.280 ;
        RECT 438.110 1.515 438.650 4.280 ;
        RECT 439.490 1.515 440.030 4.280 ;
        RECT 440.870 1.515 441.870 4.280 ;
        RECT 442.710 1.515 443.250 4.280 ;
        RECT 444.090 1.515 444.630 4.280 ;
        RECT 445.470 1.515 446.010 4.280 ;
        RECT 446.850 1.515 447.850 4.280 ;
        RECT 448.690 1.515 449.230 4.280 ;
        RECT 450.070 1.515 450.610 4.280 ;
        RECT 451.450 1.515 451.990 4.280 ;
        RECT 452.830 1.515 453.830 4.280 ;
        RECT 454.670 1.515 455.210 4.280 ;
        RECT 456.050 1.515 456.590 4.280 ;
        RECT 457.430 1.515 457.970 4.280 ;
        RECT 458.810 1.515 459.810 4.280 ;
        RECT 460.650 1.515 461.190 4.280 ;
        RECT 462.030 1.515 462.570 4.280 ;
        RECT 463.410 1.515 463.950 4.280 ;
        RECT 464.790 1.515 465.790 4.280 ;
        RECT 466.630 1.515 467.170 4.280 ;
        RECT 468.010 1.515 468.550 4.280 ;
        RECT 469.390 1.515 469.930 4.280 ;
        RECT 470.770 1.515 471.770 4.280 ;
        RECT 472.610 1.515 473.150 4.280 ;
        RECT 473.990 1.515 474.530 4.280 ;
        RECT 475.370 1.515 475.910 4.280 ;
        RECT 476.750 1.515 477.750 4.280 ;
        RECT 478.590 1.515 479.130 4.280 ;
        RECT 479.970 1.515 480.510 4.280 ;
        RECT 481.350 1.515 481.890 4.280 ;
        RECT 482.730 1.515 483.270 4.280 ;
        RECT 484.110 1.515 485.110 4.280 ;
        RECT 485.950 1.515 486.490 4.280 ;
        RECT 487.330 1.515 487.870 4.280 ;
        RECT 488.710 1.515 489.250 4.280 ;
        RECT 490.090 1.515 491.090 4.280 ;
        RECT 491.930 1.515 492.470 4.280 ;
        RECT 493.310 1.515 493.850 4.280 ;
        RECT 494.690 1.515 495.230 4.280 ;
        RECT 496.070 1.515 497.070 4.280 ;
        RECT 497.910 1.515 498.450 4.280 ;
        RECT 499.290 1.515 499.830 4.280 ;
        RECT 500.670 1.515 501.210 4.280 ;
        RECT 502.050 1.515 503.050 4.280 ;
        RECT 503.890 1.515 504.430 4.280 ;
        RECT 505.270 1.515 505.810 4.280 ;
        RECT 506.650 1.515 507.190 4.280 ;
        RECT 508.030 1.515 509.030 4.280 ;
        RECT 509.870 1.515 510.410 4.280 ;
        RECT 511.250 1.515 511.790 4.280 ;
        RECT 512.630 1.515 513.170 4.280 ;
        RECT 514.010 1.515 515.010 4.280 ;
        RECT 515.850 1.515 516.390 4.280 ;
        RECT 517.230 1.515 517.770 4.280 ;
        RECT 518.610 1.515 519.150 4.280 ;
        RECT 519.990 1.515 520.990 4.280 ;
        RECT 521.830 1.515 522.370 4.280 ;
        RECT 523.210 1.515 523.750 4.280 ;
        RECT 524.590 1.515 525.130 4.280 ;
        RECT 525.970 1.515 526.970 4.280 ;
        RECT 527.810 1.515 528.350 4.280 ;
        RECT 529.190 1.515 529.730 4.280 ;
        RECT 530.570 1.515 531.110 4.280 ;
        RECT 531.950 1.515 532.950 4.280 ;
        RECT 533.790 1.515 534.330 4.280 ;
        RECT 535.170 1.515 535.710 4.280 ;
        RECT 536.550 1.515 537.090 4.280 ;
        RECT 537.930 1.515 538.930 4.280 ;
        RECT 539.770 1.515 540.310 4.280 ;
        RECT 541.150 1.515 541.690 4.280 ;
        RECT 542.530 1.515 543.070 4.280 ;
        RECT 543.910 1.515 544.450 4.280 ;
        RECT 545.290 1.515 546.290 4.280 ;
        RECT 547.130 1.515 547.670 4.280 ;
        RECT 548.510 1.515 549.050 4.280 ;
        RECT 549.890 1.515 550.430 4.280 ;
        RECT 551.270 1.515 552.270 4.280 ;
        RECT 553.110 1.515 553.650 4.280 ;
        RECT 554.490 1.515 555.030 4.280 ;
        RECT 555.870 1.515 556.410 4.280 ;
        RECT 557.250 1.515 558.250 4.280 ;
        RECT 559.090 1.515 559.630 4.280 ;
        RECT 560.470 1.515 561.010 4.280 ;
        RECT 561.850 1.515 562.390 4.280 ;
        RECT 563.230 1.515 564.230 4.280 ;
        RECT 565.070 1.515 565.610 4.280 ;
        RECT 566.450 1.515 566.990 4.280 ;
        RECT 567.830 1.515 568.370 4.280 ;
        RECT 569.210 1.515 570.210 4.280 ;
        RECT 571.050 1.515 571.590 4.280 ;
        RECT 572.430 1.515 572.970 4.280 ;
        RECT 573.810 1.515 574.350 4.280 ;
        RECT 575.190 1.515 576.190 4.280 ;
        RECT 577.030 1.515 577.570 4.280 ;
        RECT 578.410 1.515 578.950 4.280 ;
        RECT 579.790 1.515 580.330 4.280 ;
        RECT 581.170 1.515 582.170 4.280 ;
        RECT 583.010 1.515 583.550 4.280 ;
        RECT 584.390 1.515 584.930 4.280 ;
        RECT 585.770 1.515 586.310 4.280 ;
        RECT 587.150 1.515 588.150 4.280 ;
        RECT 588.990 1.515 589.530 4.280 ;
        RECT 590.370 1.515 590.910 4.280 ;
        RECT 591.750 1.515 592.290 4.280 ;
        RECT 593.130 1.515 594.130 4.280 ;
        RECT 594.970 1.515 595.510 4.280 ;
        RECT 596.350 1.515 596.890 4.280 ;
        RECT 597.730 1.515 598.270 4.280 ;
        RECT 599.110 1.515 599.740 4.280 ;
      LAYER met3 ;
        RECT 3.285 733.400 595.600 733.545 ;
        RECT 4.400 732.680 595.600 733.400 ;
        RECT 4.400 732.000 597.015 732.680 ;
        RECT 3.285 731.360 597.015 732.000 ;
        RECT 3.285 730.000 595.600 731.360 ;
        RECT 4.400 729.960 595.600 730.000 ;
        RECT 4.400 728.640 597.015 729.960 ;
        RECT 4.400 728.600 595.600 728.640 ;
        RECT 3.285 727.240 595.600 728.600 ;
        RECT 3.285 726.600 597.015 727.240 ;
        RECT 4.400 725.920 597.015 726.600 ;
        RECT 4.400 725.200 595.600 725.920 ;
        RECT 3.285 724.520 595.600 725.200 ;
        RECT 3.285 723.200 597.015 724.520 ;
        RECT 4.400 721.800 595.600 723.200 ;
        RECT 3.285 720.480 597.015 721.800 ;
        RECT 3.285 719.800 595.600 720.480 ;
        RECT 4.400 719.080 595.600 719.800 ;
        RECT 4.400 718.400 597.015 719.080 ;
        RECT 3.285 717.760 597.015 718.400 ;
        RECT 3.285 716.400 595.600 717.760 ;
        RECT 4.400 716.360 595.600 716.400 ;
        RECT 4.400 715.040 597.015 716.360 ;
        RECT 4.400 715.000 595.600 715.040 ;
        RECT 3.285 713.640 595.600 715.000 ;
        RECT 3.285 713.000 597.015 713.640 ;
        RECT 4.400 712.320 597.015 713.000 ;
        RECT 4.400 711.600 595.600 712.320 ;
        RECT 3.285 710.920 595.600 711.600 ;
        RECT 3.285 709.600 597.015 710.920 ;
        RECT 4.400 708.200 595.600 709.600 ;
        RECT 3.285 706.880 597.015 708.200 ;
        RECT 3.285 706.200 595.600 706.880 ;
        RECT 4.400 705.480 595.600 706.200 ;
        RECT 4.400 704.800 597.015 705.480 ;
        RECT 3.285 704.160 597.015 704.800 ;
        RECT 3.285 702.800 595.600 704.160 ;
        RECT 4.400 702.760 595.600 702.800 ;
        RECT 4.400 701.440 597.015 702.760 ;
        RECT 4.400 701.400 595.600 701.440 ;
        RECT 3.285 700.040 595.600 701.400 ;
        RECT 3.285 699.400 597.015 700.040 ;
        RECT 4.400 698.720 597.015 699.400 ;
        RECT 4.400 698.000 595.600 698.720 ;
        RECT 3.285 697.320 595.600 698.000 ;
        RECT 3.285 696.000 597.015 697.320 ;
        RECT 4.400 694.600 595.600 696.000 ;
        RECT 3.285 693.280 597.015 694.600 ;
        RECT 3.285 692.600 595.600 693.280 ;
        RECT 4.400 691.880 595.600 692.600 ;
        RECT 4.400 691.200 597.015 691.880 ;
        RECT 3.285 690.560 597.015 691.200 ;
        RECT 3.285 689.200 595.600 690.560 ;
        RECT 4.400 689.160 595.600 689.200 ;
        RECT 4.400 687.840 597.015 689.160 ;
        RECT 4.400 687.800 595.600 687.840 ;
        RECT 3.285 686.440 595.600 687.800 ;
        RECT 3.285 685.800 597.015 686.440 ;
        RECT 4.400 685.120 597.015 685.800 ;
        RECT 4.400 684.400 595.600 685.120 ;
        RECT 3.285 683.720 595.600 684.400 ;
        RECT 3.285 682.400 597.015 683.720 ;
        RECT 4.400 681.000 595.600 682.400 ;
        RECT 3.285 679.680 597.015 681.000 ;
        RECT 3.285 679.000 595.600 679.680 ;
        RECT 4.400 678.280 595.600 679.000 ;
        RECT 4.400 677.600 597.015 678.280 ;
        RECT 3.285 676.960 597.015 677.600 ;
        RECT 3.285 675.600 595.600 676.960 ;
        RECT 4.400 675.560 595.600 675.600 ;
        RECT 4.400 674.240 597.015 675.560 ;
        RECT 4.400 674.200 595.600 674.240 ;
        RECT 3.285 672.840 595.600 674.200 ;
        RECT 3.285 672.200 597.015 672.840 ;
        RECT 4.400 671.520 597.015 672.200 ;
        RECT 4.400 670.800 595.600 671.520 ;
        RECT 3.285 670.120 595.600 670.800 ;
        RECT 3.285 668.800 597.015 670.120 ;
        RECT 4.400 667.400 595.600 668.800 ;
        RECT 3.285 666.080 597.015 667.400 ;
        RECT 3.285 665.400 595.600 666.080 ;
        RECT 4.400 664.680 595.600 665.400 ;
        RECT 4.400 664.000 597.015 664.680 ;
        RECT 3.285 663.360 597.015 664.000 ;
        RECT 3.285 662.000 595.600 663.360 ;
        RECT 4.400 661.960 595.600 662.000 ;
        RECT 4.400 660.640 597.015 661.960 ;
        RECT 4.400 660.600 595.600 660.640 ;
        RECT 3.285 659.240 595.600 660.600 ;
        RECT 3.285 658.600 597.015 659.240 ;
        RECT 4.400 657.920 597.015 658.600 ;
        RECT 4.400 657.200 595.600 657.920 ;
        RECT 3.285 656.520 595.600 657.200 ;
        RECT 3.285 655.200 597.015 656.520 ;
        RECT 4.400 654.520 597.015 655.200 ;
        RECT 4.400 653.800 595.600 654.520 ;
        RECT 3.285 653.120 595.600 653.800 ;
        RECT 3.285 651.800 597.015 653.120 ;
        RECT 4.400 650.400 595.600 651.800 ;
        RECT 3.285 649.080 597.015 650.400 ;
        RECT 3.285 648.400 595.600 649.080 ;
        RECT 4.400 647.680 595.600 648.400 ;
        RECT 4.400 647.000 597.015 647.680 ;
        RECT 3.285 646.360 597.015 647.000 ;
        RECT 3.285 645.000 595.600 646.360 ;
        RECT 4.400 644.960 595.600 645.000 ;
        RECT 4.400 643.640 597.015 644.960 ;
        RECT 4.400 643.600 595.600 643.640 ;
        RECT 3.285 642.240 595.600 643.600 ;
        RECT 3.285 641.600 597.015 642.240 ;
        RECT 4.400 640.920 597.015 641.600 ;
        RECT 4.400 640.200 595.600 640.920 ;
        RECT 3.285 639.520 595.600 640.200 ;
        RECT 3.285 638.200 597.015 639.520 ;
        RECT 4.400 636.800 595.600 638.200 ;
        RECT 3.285 635.480 597.015 636.800 ;
        RECT 3.285 634.800 595.600 635.480 ;
        RECT 4.400 634.080 595.600 634.800 ;
        RECT 4.400 633.400 597.015 634.080 ;
        RECT 3.285 632.760 597.015 633.400 ;
        RECT 3.285 631.400 595.600 632.760 ;
        RECT 4.400 631.360 595.600 631.400 ;
        RECT 4.400 630.040 597.015 631.360 ;
        RECT 4.400 630.000 595.600 630.040 ;
        RECT 3.285 628.640 595.600 630.000 ;
        RECT 3.285 628.000 597.015 628.640 ;
        RECT 4.400 627.320 597.015 628.000 ;
        RECT 4.400 626.600 595.600 627.320 ;
        RECT 3.285 625.920 595.600 626.600 ;
        RECT 3.285 624.600 597.015 625.920 ;
        RECT 4.400 623.200 595.600 624.600 ;
        RECT 3.285 621.880 597.015 623.200 ;
        RECT 3.285 621.200 595.600 621.880 ;
        RECT 4.400 620.480 595.600 621.200 ;
        RECT 4.400 619.800 597.015 620.480 ;
        RECT 3.285 619.160 597.015 619.800 ;
        RECT 3.285 617.800 595.600 619.160 ;
        RECT 4.400 617.760 595.600 617.800 ;
        RECT 4.400 616.440 597.015 617.760 ;
        RECT 4.400 616.400 595.600 616.440 ;
        RECT 3.285 615.040 595.600 616.400 ;
        RECT 3.285 613.720 597.015 615.040 ;
        RECT 4.400 612.320 595.600 613.720 ;
        RECT 3.285 611.000 597.015 612.320 ;
        RECT 3.285 610.320 595.600 611.000 ;
        RECT 4.400 609.600 595.600 610.320 ;
        RECT 4.400 608.920 597.015 609.600 ;
        RECT 3.285 608.280 597.015 608.920 ;
        RECT 3.285 606.920 595.600 608.280 ;
        RECT 4.400 606.880 595.600 606.920 ;
        RECT 4.400 605.560 597.015 606.880 ;
        RECT 4.400 605.520 595.600 605.560 ;
        RECT 3.285 604.160 595.600 605.520 ;
        RECT 3.285 603.520 597.015 604.160 ;
        RECT 4.400 602.840 597.015 603.520 ;
        RECT 4.400 602.120 595.600 602.840 ;
        RECT 3.285 601.440 595.600 602.120 ;
        RECT 3.285 600.120 597.015 601.440 ;
        RECT 4.400 598.720 595.600 600.120 ;
        RECT 3.285 597.400 597.015 598.720 ;
        RECT 3.285 596.720 595.600 597.400 ;
        RECT 4.400 596.000 595.600 596.720 ;
        RECT 4.400 595.320 597.015 596.000 ;
        RECT 3.285 594.680 597.015 595.320 ;
        RECT 3.285 593.320 595.600 594.680 ;
        RECT 4.400 593.280 595.600 593.320 ;
        RECT 4.400 591.960 597.015 593.280 ;
        RECT 4.400 591.920 595.600 591.960 ;
        RECT 3.285 590.560 595.600 591.920 ;
        RECT 3.285 589.920 597.015 590.560 ;
        RECT 4.400 589.240 597.015 589.920 ;
        RECT 4.400 588.520 595.600 589.240 ;
        RECT 3.285 587.840 595.600 588.520 ;
        RECT 3.285 586.520 597.015 587.840 ;
        RECT 4.400 585.120 595.600 586.520 ;
        RECT 3.285 583.800 597.015 585.120 ;
        RECT 3.285 583.120 595.600 583.800 ;
        RECT 4.400 582.400 595.600 583.120 ;
        RECT 4.400 581.720 597.015 582.400 ;
        RECT 3.285 581.080 597.015 581.720 ;
        RECT 3.285 579.720 595.600 581.080 ;
        RECT 4.400 579.680 595.600 579.720 ;
        RECT 4.400 578.360 597.015 579.680 ;
        RECT 4.400 578.320 595.600 578.360 ;
        RECT 3.285 576.960 595.600 578.320 ;
        RECT 3.285 576.320 597.015 576.960 ;
        RECT 4.400 575.640 597.015 576.320 ;
        RECT 4.400 574.920 595.600 575.640 ;
        RECT 3.285 574.240 595.600 574.920 ;
        RECT 3.285 572.920 597.015 574.240 ;
        RECT 4.400 572.240 597.015 572.920 ;
        RECT 4.400 571.520 595.600 572.240 ;
        RECT 3.285 570.840 595.600 571.520 ;
        RECT 3.285 569.520 597.015 570.840 ;
        RECT 4.400 568.120 595.600 569.520 ;
        RECT 3.285 566.800 597.015 568.120 ;
        RECT 3.285 566.120 595.600 566.800 ;
        RECT 4.400 565.400 595.600 566.120 ;
        RECT 4.400 564.720 597.015 565.400 ;
        RECT 3.285 564.080 597.015 564.720 ;
        RECT 3.285 562.720 595.600 564.080 ;
        RECT 4.400 562.680 595.600 562.720 ;
        RECT 4.400 561.360 597.015 562.680 ;
        RECT 4.400 561.320 595.600 561.360 ;
        RECT 3.285 559.960 595.600 561.320 ;
        RECT 3.285 559.320 597.015 559.960 ;
        RECT 4.400 558.640 597.015 559.320 ;
        RECT 4.400 557.920 595.600 558.640 ;
        RECT 3.285 557.240 595.600 557.920 ;
        RECT 3.285 555.920 597.015 557.240 ;
        RECT 4.400 554.520 595.600 555.920 ;
        RECT 3.285 553.200 597.015 554.520 ;
        RECT 3.285 552.520 595.600 553.200 ;
        RECT 4.400 551.800 595.600 552.520 ;
        RECT 4.400 551.120 597.015 551.800 ;
        RECT 3.285 550.480 597.015 551.120 ;
        RECT 3.285 549.120 595.600 550.480 ;
        RECT 4.400 549.080 595.600 549.120 ;
        RECT 4.400 547.760 597.015 549.080 ;
        RECT 4.400 547.720 595.600 547.760 ;
        RECT 3.285 546.360 595.600 547.720 ;
        RECT 3.285 545.720 597.015 546.360 ;
        RECT 4.400 545.040 597.015 545.720 ;
        RECT 4.400 544.320 595.600 545.040 ;
        RECT 3.285 543.640 595.600 544.320 ;
        RECT 3.285 542.320 597.015 543.640 ;
        RECT 4.400 540.920 595.600 542.320 ;
        RECT 3.285 539.600 597.015 540.920 ;
        RECT 3.285 538.920 595.600 539.600 ;
        RECT 4.400 538.200 595.600 538.920 ;
        RECT 4.400 537.520 597.015 538.200 ;
        RECT 3.285 536.880 597.015 537.520 ;
        RECT 3.285 535.520 595.600 536.880 ;
        RECT 4.400 535.480 595.600 535.520 ;
        RECT 4.400 534.160 597.015 535.480 ;
        RECT 4.400 534.120 595.600 534.160 ;
        RECT 3.285 532.760 595.600 534.120 ;
        RECT 3.285 532.120 597.015 532.760 ;
        RECT 4.400 531.440 597.015 532.120 ;
        RECT 4.400 530.720 595.600 531.440 ;
        RECT 3.285 530.040 595.600 530.720 ;
        RECT 3.285 528.720 597.015 530.040 ;
        RECT 4.400 527.320 595.600 528.720 ;
        RECT 3.285 526.000 597.015 527.320 ;
        RECT 3.285 525.320 595.600 526.000 ;
        RECT 4.400 524.600 595.600 525.320 ;
        RECT 4.400 523.920 597.015 524.600 ;
        RECT 3.285 523.280 597.015 523.920 ;
        RECT 3.285 521.920 595.600 523.280 ;
        RECT 4.400 521.880 595.600 521.920 ;
        RECT 4.400 520.560 597.015 521.880 ;
        RECT 4.400 520.520 595.600 520.560 ;
        RECT 3.285 519.160 595.600 520.520 ;
        RECT 3.285 518.520 597.015 519.160 ;
        RECT 4.400 517.840 597.015 518.520 ;
        RECT 4.400 517.120 595.600 517.840 ;
        RECT 3.285 516.440 595.600 517.120 ;
        RECT 3.285 515.120 597.015 516.440 ;
        RECT 4.400 513.720 595.600 515.120 ;
        RECT 3.285 512.400 597.015 513.720 ;
        RECT 3.285 511.720 595.600 512.400 ;
        RECT 4.400 511.000 595.600 511.720 ;
        RECT 4.400 510.320 597.015 511.000 ;
        RECT 3.285 509.680 597.015 510.320 ;
        RECT 3.285 508.320 595.600 509.680 ;
        RECT 4.400 508.280 595.600 508.320 ;
        RECT 4.400 506.960 597.015 508.280 ;
        RECT 4.400 506.920 595.600 506.960 ;
        RECT 3.285 505.560 595.600 506.920 ;
        RECT 3.285 504.920 597.015 505.560 ;
        RECT 4.400 504.240 597.015 504.920 ;
        RECT 4.400 503.520 595.600 504.240 ;
        RECT 3.285 502.840 595.600 503.520 ;
        RECT 3.285 501.520 597.015 502.840 ;
        RECT 4.400 500.120 595.600 501.520 ;
        RECT 3.285 498.800 597.015 500.120 ;
        RECT 3.285 498.120 595.600 498.800 ;
        RECT 4.400 497.400 595.600 498.120 ;
        RECT 4.400 496.720 597.015 497.400 ;
        RECT 3.285 496.080 597.015 496.720 ;
        RECT 3.285 494.720 595.600 496.080 ;
        RECT 4.400 494.680 595.600 494.720 ;
        RECT 4.400 493.360 597.015 494.680 ;
        RECT 4.400 493.320 595.600 493.360 ;
        RECT 3.285 491.960 595.600 493.320 ;
        RECT 3.285 490.640 597.015 491.960 ;
        RECT 4.400 489.960 597.015 490.640 ;
        RECT 4.400 489.240 595.600 489.960 ;
        RECT 3.285 488.560 595.600 489.240 ;
        RECT 3.285 487.240 597.015 488.560 ;
        RECT 4.400 485.840 595.600 487.240 ;
        RECT 3.285 484.520 597.015 485.840 ;
        RECT 3.285 483.840 595.600 484.520 ;
        RECT 4.400 483.120 595.600 483.840 ;
        RECT 4.400 482.440 597.015 483.120 ;
        RECT 3.285 481.800 597.015 482.440 ;
        RECT 3.285 480.440 595.600 481.800 ;
        RECT 4.400 480.400 595.600 480.440 ;
        RECT 4.400 479.080 597.015 480.400 ;
        RECT 4.400 479.040 595.600 479.080 ;
        RECT 3.285 477.680 595.600 479.040 ;
        RECT 3.285 477.040 597.015 477.680 ;
        RECT 4.400 476.360 597.015 477.040 ;
        RECT 4.400 475.640 595.600 476.360 ;
        RECT 3.285 474.960 595.600 475.640 ;
        RECT 3.285 473.640 597.015 474.960 ;
        RECT 4.400 472.240 595.600 473.640 ;
        RECT 3.285 470.920 597.015 472.240 ;
        RECT 3.285 470.240 595.600 470.920 ;
        RECT 4.400 469.520 595.600 470.240 ;
        RECT 4.400 468.840 597.015 469.520 ;
        RECT 3.285 468.200 597.015 468.840 ;
        RECT 3.285 466.840 595.600 468.200 ;
        RECT 4.400 466.800 595.600 466.840 ;
        RECT 4.400 465.480 597.015 466.800 ;
        RECT 4.400 465.440 595.600 465.480 ;
        RECT 3.285 464.080 595.600 465.440 ;
        RECT 3.285 463.440 597.015 464.080 ;
        RECT 4.400 462.760 597.015 463.440 ;
        RECT 4.400 462.040 595.600 462.760 ;
        RECT 3.285 461.360 595.600 462.040 ;
        RECT 3.285 460.040 597.015 461.360 ;
        RECT 4.400 458.640 595.600 460.040 ;
        RECT 3.285 457.320 597.015 458.640 ;
        RECT 3.285 456.640 595.600 457.320 ;
        RECT 4.400 455.920 595.600 456.640 ;
        RECT 4.400 455.240 597.015 455.920 ;
        RECT 3.285 454.600 597.015 455.240 ;
        RECT 3.285 453.240 595.600 454.600 ;
        RECT 4.400 453.200 595.600 453.240 ;
        RECT 4.400 451.880 597.015 453.200 ;
        RECT 4.400 451.840 595.600 451.880 ;
        RECT 3.285 450.480 595.600 451.840 ;
        RECT 3.285 449.840 597.015 450.480 ;
        RECT 4.400 449.160 597.015 449.840 ;
        RECT 4.400 448.440 595.600 449.160 ;
        RECT 3.285 447.760 595.600 448.440 ;
        RECT 3.285 446.440 597.015 447.760 ;
        RECT 4.400 445.040 595.600 446.440 ;
        RECT 3.285 443.720 597.015 445.040 ;
        RECT 3.285 443.040 595.600 443.720 ;
        RECT 4.400 442.320 595.600 443.040 ;
        RECT 4.400 441.640 597.015 442.320 ;
        RECT 3.285 441.000 597.015 441.640 ;
        RECT 3.285 439.640 595.600 441.000 ;
        RECT 4.400 439.600 595.600 439.640 ;
        RECT 4.400 438.280 597.015 439.600 ;
        RECT 4.400 438.240 595.600 438.280 ;
        RECT 3.285 436.880 595.600 438.240 ;
        RECT 3.285 436.240 597.015 436.880 ;
        RECT 4.400 435.560 597.015 436.240 ;
        RECT 4.400 434.840 595.600 435.560 ;
        RECT 3.285 434.160 595.600 434.840 ;
        RECT 3.285 432.840 597.015 434.160 ;
        RECT 4.400 431.440 595.600 432.840 ;
        RECT 3.285 430.120 597.015 431.440 ;
        RECT 3.285 429.440 595.600 430.120 ;
        RECT 4.400 428.720 595.600 429.440 ;
        RECT 4.400 428.040 597.015 428.720 ;
        RECT 3.285 427.400 597.015 428.040 ;
        RECT 3.285 426.040 595.600 427.400 ;
        RECT 4.400 426.000 595.600 426.040 ;
        RECT 4.400 424.680 597.015 426.000 ;
        RECT 4.400 424.640 595.600 424.680 ;
        RECT 3.285 423.280 595.600 424.640 ;
        RECT 3.285 422.640 597.015 423.280 ;
        RECT 4.400 421.960 597.015 422.640 ;
        RECT 4.400 421.240 595.600 421.960 ;
        RECT 3.285 420.560 595.600 421.240 ;
        RECT 3.285 419.240 597.015 420.560 ;
        RECT 4.400 417.840 595.600 419.240 ;
        RECT 3.285 416.520 597.015 417.840 ;
        RECT 3.285 415.840 595.600 416.520 ;
        RECT 4.400 415.120 595.600 415.840 ;
        RECT 4.400 414.440 597.015 415.120 ;
        RECT 3.285 413.800 597.015 414.440 ;
        RECT 3.285 412.440 595.600 413.800 ;
        RECT 4.400 412.400 595.600 412.440 ;
        RECT 4.400 411.080 597.015 412.400 ;
        RECT 4.400 411.040 595.600 411.080 ;
        RECT 3.285 409.680 595.600 411.040 ;
        RECT 3.285 409.040 597.015 409.680 ;
        RECT 4.400 407.680 597.015 409.040 ;
        RECT 4.400 407.640 595.600 407.680 ;
        RECT 3.285 406.280 595.600 407.640 ;
        RECT 3.285 405.640 597.015 406.280 ;
        RECT 4.400 404.960 597.015 405.640 ;
        RECT 4.400 404.240 595.600 404.960 ;
        RECT 3.285 403.560 595.600 404.240 ;
        RECT 3.285 402.240 597.015 403.560 ;
        RECT 4.400 400.840 595.600 402.240 ;
        RECT 3.285 399.520 597.015 400.840 ;
        RECT 3.285 398.840 595.600 399.520 ;
        RECT 4.400 398.120 595.600 398.840 ;
        RECT 4.400 397.440 597.015 398.120 ;
        RECT 3.285 396.800 597.015 397.440 ;
        RECT 3.285 395.440 595.600 396.800 ;
        RECT 4.400 395.400 595.600 395.440 ;
        RECT 4.400 394.080 597.015 395.400 ;
        RECT 4.400 394.040 595.600 394.080 ;
        RECT 3.285 392.680 595.600 394.040 ;
        RECT 3.285 392.040 597.015 392.680 ;
        RECT 4.400 391.360 597.015 392.040 ;
        RECT 4.400 390.640 595.600 391.360 ;
        RECT 3.285 389.960 595.600 390.640 ;
        RECT 3.285 388.640 597.015 389.960 ;
        RECT 4.400 387.240 595.600 388.640 ;
        RECT 3.285 385.920 597.015 387.240 ;
        RECT 3.285 385.240 595.600 385.920 ;
        RECT 4.400 384.520 595.600 385.240 ;
        RECT 4.400 383.840 597.015 384.520 ;
        RECT 3.285 383.200 597.015 383.840 ;
        RECT 3.285 381.840 595.600 383.200 ;
        RECT 4.400 381.800 595.600 381.840 ;
        RECT 4.400 380.480 597.015 381.800 ;
        RECT 4.400 380.440 595.600 380.480 ;
        RECT 3.285 379.080 595.600 380.440 ;
        RECT 3.285 378.440 597.015 379.080 ;
        RECT 4.400 377.760 597.015 378.440 ;
        RECT 4.400 377.040 595.600 377.760 ;
        RECT 3.285 376.360 595.600 377.040 ;
        RECT 3.285 375.040 597.015 376.360 ;
        RECT 4.400 373.640 595.600 375.040 ;
        RECT 3.285 372.320 597.015 373.640 ;
        RECT 3.285 371.640 595.600 372.320 ;
        RECT 4.400 370.920 595.600 371.640 ;
        RECT 4.400 370.240 597.015 370.920 ;
        RECT 3.285 369.600 597.015 370.240 ;
        RECT 3.285 368.200 595.600 369.600 ;
        RECT 3.285 367.560 597.015 368.200 ;
        RECT 4.400 366.880 597.015 367.560 ;
        RECT 4.400 366.160 595.600 366.880 ;
        RECT 3.285 365.480 595.600 366.160 ;
        RECT 3.285 364.160 597.015 365.480 ;
        RECT 4.400 362.760 595.600 364.160 ;
        RECT 3.285 361.440 597.015 362.760 ;
        RECT 3.285 360.760 595.600 361.440 ;
        RECT 4.400 360.040 595.600 360.760 ;
        RECT 4.400 359.360 597.015 360.040 ;
        RECT 3.285 358.720 597.015 359.360 ;
        RECT 3.285 357.360 595.600 358.720 ;
        RECT 4.400 357.320 595.600 357.360 ;
        RECT 4.400 356.000 597.015 357.320 ;
        RECT 4.400 355.960 595.600 356.000 ;
        RECT 3.285 354.600 595.600 355.960 ;
        RECT 3.285 353.960 597.015 354.600 ;
        RECT 4.400 353.280 597.015 353.960 ;
        RECT 4.400 352.560 595.600 353.280 ;
        RECT 3.285 351.880 595.600 352.560 ;
        RECT 3.285 350.560 597.015 351.880 ;
        RECT 4.400 349.160 595.600 350.560 ;
        RECT 3.285 347.840 597.015 349.160 ;
        RECT 3.285 347.160 595.600 347.840 ;
        RECT 4.400 346.440 595.600 347.160 ;
        RECT 4.400 345.760 597.015 346.440 ;
        RECT 3.285 345.120 597.015 345.760 ;
        RECT 3.285 343.760 595.600 345.120 ;
        RECT 4.400 343.720 595.600 343.760 ;
        RECT 4.400 342.400 597.015 343.720 ;
        RECT 4.400 342.360 595.600 342.400 ;
        RECT 3.285 341.000 595.600 342.360 ;
        RECT 3.285 340.360 597.015 341.000 ;
        RECT 4.400 339.680 597.015 340.360 ;
        RECT 4.400 338.960 595.600 339.680 ;
        RECT 3.285 338.280 595.600 338.960 ;
        RECT 3.285 336.960 597.015 338.280 ;
        RECT 4.400 335.560 595.600 336.960 ;
        RECT 3.285 334.240 597.015 335.560 ;
        RECT 3.285 333.560 595.600 334.240 ;
        RECT 4.400 332.840 595.600 333.560 ;
        RECT 4.400 332.160 597.015 332.840 ;
        RECT 3.285 331.520 597.015 332.160 ;
        RECT 3.285 330.160 595.600 331.520 ;
        RECT 4.400 330.120 595.600 330.160 ;
        RECT 4.400 328.760 597.015 330.120 ;
        RECT 3.285 328.120 597.015 328.760 ;
        RECT 3.285 326.760 595.600 328.120 ;
        RECT 4.400 326.720 595.600 326.760 ;
        RECT 4.400 325.400 597.015 326.720 ;
        RECT 4.400 325.360 595.600 325.400 ;
        RECT 3.285 324.000 595.600 325.360 ;
        RECT 3.285 323.360 597.015 324.000 ;
        RECT 4.400 322.680 597.015 323.360 ;
        RECT 4.400 321.960 595.600 322.680 ;
        RECT 3.285 321.280 595.600 321.960 ;
        RECT 3.285 319.960 597.015 321.280 ;
        RECT 4.400 318.560 595.600 319.960 ;
        RECT 3.285 317.240 597.015 318.560 ;
        RECT 3.285 316.560 595.600 317.240 ;
        RECT 4.400 315.840 595.600 316.560 ;
        RECT 4.400 315.160 597.015 315.840 ;
        RECT 3.285 314.520 597.015 315.160 ;
        RECT 3.285 313.160 595.600 314.520 ;
        RECT 4.400 313.120 595.600 313.160 ;
        RECT 4.400 311.800 597.015 313.120 ;
        RECT 4.400 311.760 595.600 311.800 ;
        RECT 3.285 310.400 595.600 311.760 ;
        RECT 3.285 309.760 597.015 310.400 ;
        RECT 4.400 309.080 597.015 309.760 ;
        RECT 4.400 308.360 595.600 309.080 ;
        RECT 3.285 307.680 595.600 308.360 ;
        RECT 3.285 306.360 597.015 307.680 ;
        RECT 4.400 304.960 595.600 306.360 ;
        RECT 3.285 303.640 597.015 304.960 ;
        RECT 3.285 302.960 595.600 303.640 ;
        RECT 4.400 302.240 595.600 302.960 ;
        RECT 4.400 301.560 597.015 302.240 ;
        RECT 3.285 300.920 597.015 301.560 ;
        RECT 3.285 299.560 595.600 300.920 ;
        RECT 4.400 299.520 595.600 299.560 ;
        RECT 4.400 298.200 597.015 299.520 ;
        RECT 4.400 298.160 595.600 298.200 ;
        RECT 3.285 296.800 595.600 298.160 ;
        RECT 3.285 296.160 597.015 296.800 ;
        RECT 4.400 295.480 597.015 296.160 ;
        RECT 4.400 294.760 595.600 295.480 ;
        RECT 3.285 294.080 595.600 294.760 ;
        RECT 3.285 292.760 597.015 294.080 ;
        RECT 4.400 291.360 595.600 292.760 ;
        RECT 3.285 290.040 597.015 291.360 ;
        RECT 3.285 289.360 595.600 290.040 ;
        RECT 4.400 288.640 595.600 289.360 ;
        RECT 4.400 287.960 597.015 288.640 ;
        RECT 3.285 287.320 597.015 287.960 ;
        RECT 3.285 285.960 595.600 287.320 ;
        RECT 4.400 285.920 595.600 285.960 ;
        RECT 4.400 284.600 597.015 285.920 ;
        RECT 4.400 284.560 595.600 284.600 ;
        RECT 3.285 283.200 595.600 284.560 ;
        RECT 3.285 282.560 597.015 283.200 ;
        RECT 4.400 281.880 597.015 282.560 ;
        RECT 4.400 281.160 595.600 281.880 ;
        RECT 3.285 280.480 595.600 281.160 ;
        RECT 3.285 279.160 597.015 280.480 ;
        RECT 4.400 277.760 595.600 279.160 ;
        RECT 3.285 276.440 597.015 277.760 ;
        RECT 3.285 275.760 595.600 276.440 ;
        RECT 4.400 275.040 595.600 275.760 ;
        RECT 4.400 274.360 597.015 275.040 ;
        RECT 3.285 273.720 597.015 274.360 ;
        RECT 3.285 272.360 595.600 273.720 ;
        RECT 4.400 272.320 595.600 272.360 ;
        RECT 4.400 271.000 597.015 272.320 ;
        RECT 4.400 270.960 595.600 271.000 ;
        RECT 3.285 269.600 595.600 270.960 ;
        RECT 3.285 268.960 597.015 269.600 ;
        RECT 4.400 268.280 597.015 268.960 ;
        RECT 4.400 267.560 595.600 268.280 ;
        RECT 3.285 266.880 595.600 267.560 ;
        RECT 3.285 265.560 597.015 266.880 ;
        RECT 4.400 264.160 595.600 265.560 ;
        RECT 3.285 262.840 597.015 264.160 ;
        RECT 3.285 262.160 595.600 262.840 ;
        RECT 4.400 261.440 595.600 262.160 ;
        RECT 4.400 260.760 597.015 261.440 ;
        RECT 3.285 260.120 597.015 260.760 ;
        RECT 3.285 258.760 595.600 260.120 ;
        RECT 4.400 258.720 595.600 258.760 ;
        RECT 4.400 257.400 597.015 258.720 ;
        RECT 4.400 257.360 595.600 257.400 ;
        RECT 3.285 256.000 595.600 257.360 ;
        RECT 3.285 255.360 597.015 256.000 ;
        RECT 4.400 254.680 597.015 255.360 ;
        RECT 4.400 253.960 595.600 254.680 ;
        RECT 3.285 253.280 595.600 253.960 ;
        RECT 3.285 251.960 597.015 253.280 ;
        RECT 4.400 250.560 595.600 251.960 ;
        RECT 3.285 249.240 597.015 250.560 ;
        RECT 3.285 248.560 595.600 249.240 ;
        RECT 4.400 247.840 595.600 248.560 ;
        RECT 4.400 247.160 597.015 247.840 ;
        RECT 3.285 245.840 597.015 247.160 ;
        RECT 3.285 244.480 595.600 245.840 ;
        RECT 4.400 244.440 595.600 244.480 ;
        RECT 4.400 243.120 597.015 244.440 ;
        RECT 4.400 243.080 595.600 243.120 ;
        RECT 3.285 241.720 595.600 243.080 ;
        RECT 3.285 241.080 597.015 241.720 ;
        RECT 4.400 240.400 597.015 241.080 ;
        RECT 4.400 239.680 595.600 240.400 ;
        RECT 3.285 239.000 595.600 239.680 ;
        RECT 3.285 237.680 597.015 239.000 ;
        RECT 4.400 236.280 595.600 237.680 ;
        RECT 3.285 234.960 597.015 236.280 ;
        RECT 3.285 234.280 595.600 234.960 ;
        RECT 4.400 233.560 595.600 234.280 ;
        RECT 4.400 232.880 597.015 233.560 ;
        RECT 3.285 232.240 597.015 232.880 ;
        RECT 3.285 230.880 595.600 232.240 ;
        RECT 4.400 230.840 595.600 230.880 ;
        RECT 4.400 229.520 597.015 230.840 ;
        RECT 4.400 229.480 595.600 229.520 ;
        RECT 3.285 228.120 595.600 229.480 ;
        RECT 3.285 227.480 597.015 228.120 ;
        RECT 4.400 226.800 597.015 227.480 ;
        RECT 4.400 226.080 595.600 226.800 ;
        RECT 3.285 225.400 595.600 226.080 ;
        RECT 3.285 224.080 597.015 225.400 ;
        RECT 4.400 222.680 595.600 224.080 ;
        RECT 3.285 221.360 597.015 222.680 ;
        RECT 3.285 220.680 595.600 221.360 ;
        RECT 4.400 219.960 595.600 220.680 ;
        RECT 4.400 219.280 597.015 219.960 ;
        RECT 3.285 218.640 597.015 219.280 ;
        RECT 3.285 217.280 595.600 218.640 ;
        RECT 4.400 217.240 595.600 217.280 ;
        RECT 4.400 215.920 597.015 217.240 ;
        RECT 4.400 215.880 595.600 215.920 ;
        RECT 3.285 214.520 595.600 215.880 ;
        RECT 3.285 213.880 597.015 214.520 ;
        RECT 4.400 213.200 597.015 213.880 ;
        RECT 4.400 212.480 595.600 213.200 ;
        RECT 3.285 211.800 595.600 212.480 ;
        RECT 3.285 210.480 597.015 211.800 ;
        RECT 4.400 209.080 595.600 210.480 ;
        RECT 3.285 207.760 597.015 209.080 ;
        RECT 3.285 207.080 595.600 207.760 ;
        RECT 4.400 206.360 595.600 207.080 ;
        RECT 4.400 205.680 597.015 206.360 ;
        RECT 3.285 205.040 597.015 205.680 ;
        RECT 3.285 203.680 595.600 205.040 ;
        RECT 4.400 203.640 595.600 203.680 ;
        RECT 4.400 202.320 597.015 203.640 ;
        RECT 4.400 202.280 595.600 202.320 ;
        RECT 3.285 200.920 595.600 202.280 ;
        RECT 3.285 200.280 597.015 200.920 ;
        RECT 4.400 199.600 597.015 200.280 ;
        RECT 4.400 198.880 595.600 199.600 ;
        RECT 3.285 198.200 595.600 198.880 ;
        RECT 3.285 196.880 597.015 198.200 ;
        RECT 4.400 195.480 595.600 196.880 ;
        RECT 3.285 194.160 597.015 195.480 ;
        RECT 3.285 193.480 595.600 194.160 ;
        RECT 4.400 192.760 595.600 193.480 ;
        RECT 4.400 192.080 597.015 192.760 ;
        RECT 3.285 191.440 597.015 192.080 ;
        RECT 3.285 190.080 595.600 191.440 ;
        RECT 4.400 190.040 595.600 190.080 ;
        RECT 4.400 188.720 597.015 190.040 ;
        RECT 4.400 188.680 595.600 188.720 ;
        RECT 3.285 187.320 595.600 188.680 ;
        RECT 3.285 186.680 597.015 187.320 ;
        RECT 4.400 186.000 597.015 186.680 ;
        RECT 4.400 185.280 595.600 186.000 ;
        RECT 3.285 184.600 595.600 185.280 ;
        RECT 3.285 183.280 597.015 184.600 ;
        RECT 4.400 181.880 595.600 183.280 ;
        RECT 3.285 180.560 597.015 181.880 ;
        RECT 3.285 179.880 595.600 180.560 ;
        RECT 4.400 179.160 595.600 179.880 ;
        RECT 4.400 178.480 597.015 179.160 ;
        RECT 3.285 177.840 597.015 178.480 ;
        RECT 3.285 176.480 595.600 177.840 ;
        RECT 4.400 176.440 595.600 176.480 ;
        RECT 4.400 175.120 597.015 176.440 ;
        RECT 4.400 175.080 595.600 175.120 ;
        RECT 3.285 173.720 595.600 175.080 ;
        RECT 3.285 173.080 597.015 173.720 ;
        RECT 4.400 172.400 597.015 173.080 ;
        RECT 4.400 171.680 595.600 172.400 ;
        RECT 3.285 171.000 595.600 171.680 ;
        RECT 3.285 169.680 597.015 171.000 ;
        RECT 4.400 168.280 595.600 169.680 ;
        RECT 3.285 166.960 597.015 168.280 ;
        RECT 3.285 166.280 595.600 166.960 ;
        RECT 4.400 165.560 595.600 166.280 ;
        RECT 4.400 164.880 597.015 165.560 ;
        RECT 3.285 163.560 597.015 164.880 ;
        RECT 3.285 162.880 595.600 163.560 ;
        RECT 4.400 162.160 595.600 162.880 ;
        RECT 4.400 161.480 597.015 162.160 ;
        RECT 3.285 160.840 597.015 161.480 ;
        RECT 3.285 159.480 595.600 160.840 ;
        RECT 4.400 159.440 595.600 159.480 ;
        RECT 4.400 158.120 597.015 159.440 ;
        RECT 4.400 158.080 595.600 158.120 ;
        RECT 3.285 156.720 595.600 158.080 ;
        RECT 3.285 156.080 597.015 156.720 ;
        RECT 4.400 155.400 597.015 156.080 ;
        RECT 4.400 154.680 595.600 155.400 ;
        RECT 3.285 154.000 595.600 154.680 ;
        RECT 3.285 152.680 597.015 154.000 ;
        RECT 4.400 151.280 595.600 152.680 ;
        RECT 3.285 149.960 597.015 151.280 ;
        RECT 3.285 149.280 595.600 149.960 ;
        RECT 4.400 148.560 595.600 149.280 ;
        RECT 4.400 147.880 597.015 148.560 ;
        RECT 3.285 147.240 597.015 147.880 ;
        RECT 3.285 145.880 595.600 147.240 ;
        RECT 4.400 145.840 595.600 145.880 ;
        RECT 4.400 144.520 597.015 145.840 ;
        RECT 4.400 144.480 595.600 144.520 ;
        RECT 3.285 143.120 595.600 144.480 ;
        RECT 3.285 142.480 597.015 143.120 ;
        RECT 4.400 141.800 597.015 142.480 ;
        RECT 4.400 141.080 595.600 141.800 ;
        RECT 3.285 140.400 595.600 141.080 ;
        RECT 3.285 139.080 597.015 140.400 ;
        RECT 4.400 137.680 595.600 139.080 ;
        RECT 3.285 136.360 597.015 137.680 ;
        RECT 3.285 135.680 595.600 136.360 ;
        RECT 4.400 134.960 595.600 135.680 ;
        RECT 4.400 134.280 597.015 134.960 ;
        RECT 3.285 133.640 597.015 134.280 ;
        RECT 3.285 132.280 595.600 133.640 ;
        RECT 4.400 132.240 595.600 132.280 ;
        RECT 4.400 130.920 597.015 132.240 ;
        RECT 4.400 130.880 595.600 130.920 ;
        RECT 3.285 129.520 595.600 130.880 ;
        RECT 3.285 128.880 597.015 129.520 ;
        RECT 4.400 128.200 597.015 128.880 ;
        RECT 4.400 127.480 595.600 128.200 ;
        RECT 3.285 126.800 595.600 127.480 ;
        RECT 3.285 125.480 597.015 126.800 ;
        RECT 4.400 124.080 595.600 125.480 ;
        RECT 3.285 122.760 597.015 124.080 ;
        RECT 3.285 121.400 595.600 122.760 ;
        RECT 4.400 121.360 595.600 121.400 ;
        RECT 4.400 120.040 597.015 121.360 ;
        RECT 4.400 120.000 595.600 120.040 ;
        RECT 3.285 118.640 595.600 120.000 ;
        RECT 3.285 118.000 597.015 118.640 ;
        RECT 4.400 117.320 597.015 118.000 ;
        RECT 4.400 116.600 595.600 117.320 ;
        RECT 3.285 115.920 595.600 116.600 ;
        RECT 3.285 114.600 597.015 115.920 ;
        RECT 4.400 113.200 595.600 114.600 ;
        RECT 3.285 111.880 597.015 113.200 ;
        RECT 3.285 111.200 595.600 111.880 ;
        RECT 4.400 110.480 595.600 111.200 ;
        RECT 4.400 109.800 597.015 110.480 ;
        RECT 3.285 109.160 597.015 109.800 ;
        RECT 3.285 107.800 595.600 109.160 ;
        RECT 4.400 107.760 595.600 107.800 ;
        RECT 4.400 106.440 597.015 107.760 ;
        RECT 4.400 106.400 595.600 106.440 ;
        RECT 3.285 105.040 595.600 106.400 ;
        RECT 3.285 104.400 597.015 105.040 ;
        RECT 4.400 103.720 597.015 104.400 ;
        RECT 4.400 103.000 595.600 103.720 ;
        RECT 3.285 102.320 595.600 103.000 ;
        RECT 3.285 101.000 597.015 102.320 ;
        RECT 4.400 99.600 595.600 101.000 ;
        RECT 3.285 98.280 597.015 99.600 ;
        RECT 3.285 97.600 595.600 98.280 ;
        RECT 4.400 96.880 595.600 97.600 ;
        RECT 4.400 96.200 597.015 96.880 ;
        RECT 3.285 95.560 597.015 96.200 ;
        RECT 3.285 94.200 595.600 95.560 ;
        RECT 4.400 94.160 595.600 94.200 ;
        RECT 4.400 92.840 597.015 94.160 ;
        RECT 4.400 92.800 595.600 92.840 ;
        RECT 3.285 91.440 595.600 92.800 ;
        RECT 3.285 90.800 597.015 91.440 ;
        RECT 4.400 90.120 597.015 90.800 ;
        RECT 4.400 89.400 595.600 90.120 ;
        RECT 3.285 88.720 595.600 89.400 ;
        RECT 3.285 87.400 597.015 88.720 ;
        RECT 4.400 86.000 595.600 87.400 ;
        RECT 3.285 84.680 597.015 86.000 ;
        RECT 3.285 84.000 595.600 84.680 ;
        RECT 4.400 83.280 595.600 84.000 ;
        RECT 4.400 82.600 597.015 83.280 ;
        RECT 3.285 81.280 597.015 82.600 ;
        RECT 3.285 80.600 595.600 81.280 ;
        RECT 4.400 79.880 595.600 80.600 ;
        RECT 4.400 79.200 597.015 79.880 ;
        RECT 3.285 78.560 597.015 79.200 ;
        RECT 3.285 77.200 595.600 78.560 ;
        RECT 4.400 77.160 595.600 77.200 ;
        RECT 4.400 75.840 597.015 77.160 ;
        RECT 4.400 75.800 595.600 75.840 ;
        RECT 3.285 74.440 595.600 75.800 ;
        RECT 3.285 73.800 597.015 74.440 ;
        RECT 4.400 73.120 597.015 73.800 ;
        RECT 4.400 72.400 595.600 73.120 ;
        RECT 3.285 71.720 595.600 72.400 ;
        RECT 3.285 70.400 597.015 71.720 ;
        RECT 4.400 69.000 595.600 70.400 ;
        RECT 3.285 67.680 597.015 69.000 ;
        RECT 3.285 67.000 595.600 67.680 ;
        RECT 4.400 66.280 595.600 67.000 ;
        RECT 4.400 65.600 597.015 66.280 ;
        RECT 3.285 64.960 597.015 65.600 ;
        RECT 3.285 63.600 595.600 64.960 ;
        RECT 4.400 63.560 595.600 63.600 ;
        RECT 4.400 62.240 597.015 63.560 ;
        RECT 4.400 62.200 595.600 62.240 ;
        RECT 3.285 60.840 595.600 62.200 ;
        RECT 3.285 60.200 597.015 60.840 ;
        RECT 4.400 59.520 597.015 60.200 ;
        RECT 4.400 58.800 595.600 59.520 ;
        RECT 3.285 58.120 595.600 58.800 ;
        RECT 3.285 56.800 597.015 58.120 ;
        RECT 4.400 55.400 595.600 56.800 ;
        RECT 3.285 54.080 597.015 55.400 ;
        RECT 3.285 53.400 595.600 54.080 ;
        RECT 4.400 52.680 595.600 53.400 ;
        RECT 4.400 52.000 597.015 52.680 ;
        RECT 3.285 51.360 597.015 52.000 ;
        RECT 3.285 50.000 595.600 51.360 ;
        RECT 4.400 49.960 595.600 50.000 ;
        RECT 4.400 48.640 597.015 49.960 ;
        RECT 4.400 48.600 595.600 48.640 ;
        RECT 3.285 47.240 595.600 48.600 ;
        RECT 3.285 46.600 597.015 47.240 ;
        RECT 4.400 45.920 597.015 46.600 ;
        RECT 4.400 45.200 595.600 45.920 ;
        RECT 3.285 44.520 595.600 45.200 ;
        RECT 3.285 43.200 597.015 44.520 ;
        RECT 4.400 41.800 595.600 43.200 ;
        RECT 3.285 40.480 597.015 41.800 ;
        RECT 3.285 39.800 595.600 40.480 ;
        RECT 4.400 39.080 595.600 39.800 ;
        RECT 4.400 38.400 597.015 39.080 ;
        RECT 3.285 37.760 597.015 38.400 ;
        RECT 3.285 36.400 595.600 37.760 ;
        RECT 4.400 36.360 595.600 36.400 ;
        RECT 4.400 35.040 597.015 36.360 ;
        RECT 4.400 35.000 595.600 35.040 ;
        RECT 3.285 33.640 595.600 35.000 ;
        RECT 3.285 33.000 597.015 33.640 ;
        RECT 4.400 32.320 597.015 33.000 ;
        RECT 4.400 31.600 595.600 32.320 ;
        RECT 3.285 30.920 595.600 31.600 ;
        RECT 3.285 29.600 597.015 30.920 ;
        RECT 4.400 28.200 595.600 29.600 ;
        RECT 3.285 26.880 597.015 28.200 ;
        RECT 3.285 26.200 595.600 26.880 ;
        RECT 4.400 25.480 595.600 26.200 ;
        RECT 4.400 24.800 597.015 25.480 ;
        RECT 3.285 24.160 597.015 24.800 ;
        RECT 3.285 22.800 595.600 24.160 ;
        RECT 4.400 22.760 595.600 22.800 ;
        RECT 4.400 21.440 597.015 22.760 ;
        RECT 4.400 21.400 595.600 21.440 ;
        RECT 3.285 20.040 595.600 21.400 ;
        RECT 3.285 19.400 597.015 20.040 ;
        RECT 4.400 18.720 597.015 19.400 ;
        RECT 4.400 18.000 595.600 18.720 ;
        RECT 3.285 17.320 595.600 18.000 ;
        RECT 3.285 16.000 597.015 17.320 ;
        RECT 4.400 14.600 595.600 16.000 ;
        RECT 3.285 13.280 597.015 14.600 ;
        RECT 3.285 12.600 595.600 13.280 ;
        RECT 4.400 11.880 595.600 12.600 ;
        RECT 4.400 11.200 597.015 11.880 ;
        RECT 3.285 10.560 597.015 11.200 ;
        RECT 3.285 9.200 595.600 10.560 ;
        RECT 4.400 9.160 595.600 9.200 ;
        RECT 4.400 7.840 597.015 9.160 ;
        RECT 4.400 7.800 595.600 7.840 ;
        RECT 3.285 6.440 595.600 7.800 ;
        RECT 3.285 5.800 597.015 6.440 ;
        RECT 4.400 5.120 597.015 5.800 ;
        RECT 4.400 4.400 595.600 5.120 ;
        RECT 3.285 3.720 595.600 4.400 ;
        RECT 3.285 2.400 597.015 3.720 ;
        RECT 4.400 1.535 595.600 2.400 ;
      LAYER met4 ;
        RECT 9.495 10.240 20.640 441.825 ;
        RECT 23.040 10.240 97.440 441.825 ;
        RECT 99.840 10.240 174.240 441.825 ;
        RECT 176.640 10.240 251.040 441.825 ;
        RECT 253.440 10.240 327.840 441.825 ;
        RECT 330.240 10.240 404.640 441.825 ;
        RECT 407.040 10.240 481.440 441.825 ;
        RECT 483.840 10.240 558.240 441.825 ;
        RECT 560.640 10.240 586.665 441.825 ;
        RECT 9.495 4.255 586.665 10.240 ;
  END
END main_controller
END LIBRARY

