VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1375.380 2924.800 1376.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 3517.600 2266.930 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 3517.600 1959.650 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 3517.600 1652.370 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 3517.600 1344.630 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 3517.600 1037.350 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 3517.600 730.070 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 3517.600 422.790 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3487.460 2.400 3488.660 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3235.860 2.400 3237.060 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2984.940 2.400 2986.140 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1631.060 2924.800 1632.260 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2733.340 2.400 2734.540 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2481.740 2.400 2482.940 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2230.820 2.400 2232.020 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1979.220 2.400 1980.420 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1727.620 2.400 1728.820 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1476.020 2.400 1477.220 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1225.100 2.400 1226.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 973.500 2.400 974.700 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 721.900 2.400 723.100 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1887.420 2924.800 1888.620 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2143.100 2924.800 2144.300 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2399.460 2924.800 2400.660 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2655.140 2924.800 2656.340 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2910.820 2924.800 2912.020 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3167.180 2924.800 3168.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2880.930 3517.600 2881.490 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 3517.600 2574.210 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 31.700 2924.800 32.900 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2207.020 2924.800 2208.220 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2463.380 2924.800 2464.580 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2719.060 2924.800 2720.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2975.420 2924.800 2976.620 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3231.100 2924.800 3232.300 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 3517.600 2804.670 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 3517.600 2497.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 3517.600 2190.110 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 3517.600 1882.830 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 3517.600 1575.550 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 223.460 2924.800 224.660 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 3517.600 1267.810 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 3517.600 960.530 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 3517.600 653.250 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 3517.600 345.970 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3424.900 2.400 3426.100 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3173.300 2.400 3174.500 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2921.700 2.400 2922.900 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2670.780 2.400 2671.980 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2419.180 2.400 2420.380 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2167.580 2.400 2168.780 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 415.220 2924.800 416.420 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1915.980 2.400 1917.180 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1665.060 2.400 1666.260 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1413.460 2.400 1414.660 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1161.860 2.400 1163.060 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 910.940 2.400 912.140 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 659.340 2.400 660.540 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 470.980 2.400 472.180 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 281.940 2.400 283.140 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 606.980 2924.800 608.180 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 799.420 2924.800 800.620 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 991.180 2924.800 992.380 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1182.940 2924.800 1184.140 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1439.300 2924.800 1440.500 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1694.980 2924.800 1696.180 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1951.340 2924.800 1952.540 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 159.540 2924.800 160.740 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2334.860 2924.800 2336.060 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2591.220 2924.800 2592.420 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2846.900 2924.800 2848.100 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3103.260 2924.800 3104.460 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3358.940 2924.800 3360.140 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 3517.600 2651.030 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 3517.600 2343.750 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 3517.600 2036.470 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 3517.600 1729.190 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.890 3517.600 1421.450 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 351.300 2924.800 352.500 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 3517.600 1114.170 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 3517.600 806.890 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 3517.600 499.610 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 3517.600 192.330 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3299.100 2.400 3300.300 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3047.500 2.400 3048.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2795.900 2.400 2797.100 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2544.980 2.400 2546.180 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2293.380 2.400 2294.580 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2041.780 2.400 2042.980 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 543.060 2924.800 544.260 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1790.860 2.400 1792.060 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1539.260 2.400 1540.460 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1287.660 2.400 1288.860 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1036.060 2.400 1037.260 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 785.140 2.400 786.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 533.540 2.400 534.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 345.180 2.400 346.380 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 156.140 2.400 157.340 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 735.500 2924.800 736.700 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 927.260 2924.800 928.460 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1119.020 2924.800 1120.220 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1311.460 2924.800 1312.660 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1567.140 2924.800 1568.340 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1823.500 2924.800 1824.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2079.180 2924.800 2080.380 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 95.620 2924.800 96.820 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2270.940 2924.800 2272.140 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2527.300 2924.800 2528.500 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2782.980 2924.800 2784.180 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3039.340 2924.800 3040.540 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3295.020 2924.800 3296.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 3517.600 2727.850 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 3517.600 2420.570 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 3517.600 2113.290 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 3517.600 1806.010 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 3517.600 1498.730 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 287.380 2924.800 288.580 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 3517.600 1190.990 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 3517.600 883.710 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 3517.600 576.430 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 3517.600 269.150 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3361.660 2.400 3362.860 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3110.740 2.400 3111.940 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2859.140 2.400 2860.340 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2607.540 2.400 2608.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2355.940 2.400 2357.140 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2105.020 2.400 2106.220 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 479.140 2924.800 480.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1853.420 2.400 1854.620 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1601.820 2.400 1603.020 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1350.900 2.400 1352.100 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1099.300 2.400 1100.500 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 847.700 2.400 848.900 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 596.100 2.400 597.300 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 407.740 2.400 408.940 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 219.380 2.400 220.580 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 671.580 2924.800 672.780 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 863.340 2924.800 864.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1055.100 2924.800 1056.300 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1247.540 2924.800 1248.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1503.220 2924.800 1504.420 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2015.260 2924.800 2016.460 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.470 -4.800 627.030 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.870 -4.800 2393.430 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2410.350 -4.800 2410.910 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2427.830 -4.800 2428.390 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2445.770 -4.800 2446.330 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.250 -4.800 2463.810 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2481.190 -4.800 2481.750 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2498.670 -4.800 2499.230 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.150 -4.800 2516.710 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2534.090 -4.800 2534.650 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2551.570 -4.800 2552.130 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.110 -4.800 803.670 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2569.510 -4.800 2570.070 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2586.990 -4.800 2587.550 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2604.470 -4.800 2605.030 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2622.410 -4.800 2622.970 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2639.890 -4.800 2640.450 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2657.830 -4.800 2658.390 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2675.310 -4.800 2675.870 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2692.790 -4.800 2693.350 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2710.730 -4.800 2711.290 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2728.210 -4.800 2728.770 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.590 -4.800 821.150 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2746.150 -4.800 2746.710 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.630 -4.800 2764.190 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2781.110 -4.800 2781.670 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2799.050 -4.800 2799.610 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.530 -4.800 2817.090 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.470 -4.800 2835.030 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.950 -4.800 2852.510 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.530 -4.800 839.090 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.010 -4.800 856.570 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.950 -4.800 874.510 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.430 -4.800 891.990 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.910 -4.800 909.470 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.850 -4.800 927.410 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.330 -4.800 944.890 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.270 -4.800 962.830 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.410 -4.800 644.970 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.750 -4.800 980.310 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.230 -4.800 997.790 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.170 -4.800 1015.730 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.650 -4.800 1033.210 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.590 -4.800 1051.150 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.070 -4.800 1068.630 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.550 -4.800 1086.110 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.490 -4.800 1104.050 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.970 -4.800 1121.530 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.910 -4.800 1139.470 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.890 -4.800 662.450 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.290 -4.800 1209.850 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.230 -4.800 1227.790 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.710 -4.800 1245.270 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.190 -4.800 1262.750 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.130 -4.800 1280.690 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.610 -4.800 1298.170 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.550 -4.800 1316.110 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.370 -4.800 679.930 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.030 -4.800 1333.590 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.510 -4.800 1351.070 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.450 -4.800 1369.010 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.930 -4.800 1386.490 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.870 -4.800 1404.430 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.730 -4.800 1492.290 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.310 -4.800 697.870 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.150 -4.800 1527.710 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.570 -4.800 1563.130 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.050 -4.800 1580.610 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.990 -4.800 1598.550 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.470 -4.800 1616.030 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.410 -4.800 1633.970 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.890 -4.800 1651.450 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.370 -4.800 1668.930 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.790 -4.800 715.350 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.310 -4.800 1686.870 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.790 -4.800 1704.350 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.730 -4.800 1722.290 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.110 -4.800 1792.670 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.050 -4.800 1810.610 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.530 -4.800 1828.090 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.010 -4.800 1845.570 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.730 -4.800 733.290 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.950 -4.800 1863.510 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.430 -4.800 1880.990 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.370 -4.800 1898.930 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.850 -4.800 1916.410 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.330 -4.800 1933.890 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.270 -4.800 1951.830 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.750 -4.800 1969.310 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.690 -4.800 1987.250 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2004.170 -4.800 2004.730 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.650 -4.800 2022.210 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.210 -4.800 750.770 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.590 -4.800 2040.150 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.070 -4.800 2057.630 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.010 -4.800 2075.570 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.490 -4.800 2093.050 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.970 -4.800 2110.530 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2127.910 -4.800 2128.470 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.390 -4.800 2145.950 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.330 -4.800 2163.890 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.810 -4.800 2181.370 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.290 -4.800 2198.850 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.690 -4.800 768.250 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2216.230 -4.800 2216.790 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2233.710 -4.800 2234.270 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.190 -4.800 2251.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2269.130 -4.800 2269.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.610 -4.800 2287.170 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.550 -4.800 2305.110 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.930 -4.800 2375.490 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.630 -4.800 786.190 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.450 -4.800 633.010 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.390 -4.800 2398.950 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.330 -4.800 2416.890 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.810 -4.800 2434.370 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2451.750 -4.800 2452.310 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2469.230 -4.800 2469.790 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2486.710 -4.800 2487.270 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2504.650 -4.800 2505.210 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2522.130 -4.800 2522.690 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2540.070 -4.800 2540.630 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2557.550 -4.800 2558.110 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.090 -4.800 809.650 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.030 -4.800 2575.590 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2592.970 -4.800 2593.530 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2610.450 -4.800 2611.010 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2628.390 -4.800 2628.950 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2645.870 -4.800 2646.430 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2663.350 -4.800 2663.910 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2681.290 -4.800 2681.850 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2698.770 -4.800 2699.330 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2716.710 -4.800 2717.270 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2734.190 -4.800 2734.750 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.570 -4.800 827.130 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.670 -4.800 2752.230 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2769.610 -4.800 2770.170 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2787.090 -4.800 2787.650 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2805.030 -4.800 2805.590 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.510 -4.800 2823.070 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.930 -4.800 2858.490 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.510 -4.800 845.070 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.990 -4.800 862.550 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.470 -4.800 880.030 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.410 -4.800 897.970 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.890 -4.800 915.450 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.830 -4.800 933.390 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.310 -4.800 950.870 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.790 -4.800 968.350 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.930 -4.800 650.490 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.730 -4.800 986.290 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.210 -4.800 1003.770 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.150 -4.800 1021.710 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.630 -4.800 1039.190 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.110 -4.800 1056.670 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.050 -4.800 1074.610 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.530 -4.800 1092.090 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.470 -4.800 1110.030 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.950 -4.800 1127.510 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.870 -4.800 668.430 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.270 -4.800 1215.830 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.750 -4.800 1233.310 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.690 -4.800 1251.250 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.170 -4.800 1268.730 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.110 -4.800 1286.670 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.590 -4.800 1304.150 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.070 -4.800 1321.630 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.350 -4.800 685.910 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.010 -4.800 1339.570 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.490 -4.800 1357.050 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.430 -4.800 1374.990 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.910 -4.800 1392.470 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.330 -4.800 1427.890 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.710 -4.800 1498.270 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.290 -4.800 703.850 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.130 -4.800 1533.690 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.610 -4.800 1551.170 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.550 -4.800 1569.110 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.030 -4.800 1586.590 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.970 -4.800 1604.530 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.450 -4.800 1622.010 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.930 -4.800 1639.490 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.870 -4.800 1657.430 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.350 -4.800 1674.910 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.770 -4.800 721.330 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.290 -4.800 1692.850 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.770 -4.800 1710.330 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.090 -4.800 1798.650 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.570 -4.800 1816.130 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1833.510 -4.800 1834.070 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.990 -4.800 1851.550 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.250 -4.800 738.810 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.930 -4.800 1869.490 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.410 -4.800 1886.970 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.890 -4.800 1904.450 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.830 -4.800 1922.390 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1939.310 -4.800 1939.870 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.250 -4.800 1957.810 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1974.730 -4.800 1975.290 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1992.210 -4.800 1992.770 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2010.150 -4.800 2010.710 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.630 -4.800 2028.190 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.190 -4.800 756.750 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.570 -4.800 2046.130 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.050 -4.800 2063.610 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.530 -4.800 2081.090 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.470 -4.800 2099.030 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.950 -4.800 2116.510 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2133.890 -4.800 2134.450 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.370 -4.800 2151.930 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.850 -4.800 2169.410 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.790 -4.800 2187.350 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.270 -4.800 2204.830 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.670 -4.800 774.230 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.750 -4.800 2222.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2239.690 -4.800 2240.250 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.170 -4.800 2257.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2275.110 -4.800 2275.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.590 -4.800 2293.150 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2380.910 -4.800 2381.470 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.150 -4.800 791.710 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.430 -4.800 638.990 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2404.370 -4.800 2404.930 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.310 -4.800 2422.870 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.790 -4.800 2440.350 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2457.270 -4.800 2457.830 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2475.210 -4.800 2475.770 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.690 -4.800 2493.250 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2510.630 -4.800 2511.190 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2528.110 -4.800 2528.670 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2545.590 -4.800 2546.150 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2563.530 -4.800 2564.090 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.070 -4.800 815.630 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2581.010 -4.800 2581.570 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2598.950 -4.800 2599.510 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2616.430 -4.800 2616.990 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2633.910 -4.800 2634.470 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2651.850 -4.800 2652.410 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2669.330 -4.800 2669.890 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2687.270 -4.800 2687.830 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2704.750 -4.800 2705.310 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2722.230 -4.800 2722.790 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2740.170 -4.800 2740.730 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.550 -4.800 833.110 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.650 -4.800 2758.210 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2775.590 -4.800 2776.150 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2793.070 -4.800 2793.630 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.550 -4.800 2811.110 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.490 -4.800 2829.050 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.970 -4.800 2846.530 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.910 -4.800 2864.470 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.030 -4.800 850.590 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.970 -4.800 868.530 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.450 -4.800 886.010 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.390 -4.800 903.950 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.870 -4.800 921.430 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.350 -4.800 938.910 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.290 -4.800 956.850 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.770 -4.800 974.330 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.910 -4.800 656.470 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.710 -4.800 992.270 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.190 -4.800 1009.750 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.670 -4.800 1027.230 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.610 -4.800 1045.170 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.090 -4.800 1062.650 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.030 -4.800 1080.590 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.510 -4.800 1098.070 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.990 -4.800 1115.550 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.930 -4.800 1133.490 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.850 -4.800 674.410 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.310 -4.800 1203.870 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.250 -4.800 1221.810 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.730 -4.800 1239.290 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.670 -4.800 1257.230 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.150 -4.800 1274.710 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.630 -4.800 1292.190 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.570 -4.800 1310.130 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.050 -4.800 1327.610 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.330 -4.800 691.890 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.990 -4.800 1345.550 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.470 -4.800 1363.030 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.890 -4.800 1398.450 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.310 -4.800 1433.870 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.810 -4.800 709.370 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.170 -4.800 1521.730 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.110 -4.800 1539.670 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.590 -4.800 1557.150 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.530 -4.800 1575.090 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.010 -4.800 1592.570 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.490 -4.800 1610.050 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.430 -4.800 1627.990 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.910 -4.800 1645.470 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.850 -4.800 1663.410 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.330 -4.800 1680.890 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.750 -4.800 727.310 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.810 -4.800 1698.370 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.750 -4.800 1716.310 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.130 -4.800 1786.690 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.070 -4.800 1804.630 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.550 -4.800 1822.110 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.490 -4.800 1840.050 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1856.970 -4.800 1857.530 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.230 -4.800 744.790 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.450 -4.800 1875.010 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.390 -4.800 1892.950 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.870 -4.800 1910.430 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.810 -4.800 1928.370 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.290 -4.800 1945.850 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.770 -4.800 1963.330 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.710 -4.800 1981.270 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.190 -4.800 1998.750 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2016.130 -4.800 2016.690 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.610 -4.800 2034.170 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.710 -4.800 762.270 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.090 -4.800 2051.650 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.030 -4.800 2069.590 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.510 -4.800 2087.070 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2104.450 -4.800 2105.010 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.930 -4.800 2122.490 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2139.410 -4.800 2139.970 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.350 -4.800 2157.910 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.830 -4.800 2175.390 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.770 -4.800 2193.330 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.250 -4.800 2210.810 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.650 -4.800 780.210 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2227.730 -4.800 2228.290 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2245.670 -4.800 2246.230 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.150 -4.800 2263.710 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.630 -4.800 2281.190 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.570 -4.800 2299.130 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.950 -4.800 2369.510 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.890 -4.800 2387.450 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.130 -4.800 797.690 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2887.370 -4.800 2887.930 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2893.350 -4.800 2893.910 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.330 2934.450 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 194.330 2934.450 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 374.330 2934.450 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 554.330 2934.450 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 734.330 2934.450 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 914.330 2934.450 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1094.330 2934.450 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1274.330 2934.450 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1454.330 2934.450 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1634.330 2934.450 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1814.330 2934.450 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1994.330 2934.450 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2174.330 2934.450 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2354.330 2934.450 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2534.330 2934.450 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2714.330 2934.450 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 368.970 2809.030 1272.070 2812.130 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2894.330 2934.450 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3074.330 2934.450 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3254.330 2934.450 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3434.330 2934.450 3437.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -9.470 372.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -9.470 552.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -9.470 732.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -9.470 912.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -9.470 1092.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -9.470 1272.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -9.470 1452.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -9.470 1632.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -9.470 1992.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -9.470 2172.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -9.470 2352.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -9.470 2532.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 651.540 372.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 651.540 552.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 651.540 732.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 651.540 912.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 651.540 1092.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 651.540 1272.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 651.540 1452.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 651.540 1632.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 651.540 1992.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 651.540 2172.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 651.540 2352.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 651.540 2532.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1201.540 372.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1201.540 552.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1201.540 732.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 1201.540 912.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 1201.540 1092.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 1201.540 1272.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 1201.540 1452.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 1201.540 1632.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 1201.540 1992.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1201.540 2172.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1201.540 2352.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1201.540 2532.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1751.540 372.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1751.540 552.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1751.540 732.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 1751.540 912.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 1751.540 1092.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 1751.540 1272.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 1751.540 1452.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 1751.540 1632.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 1751.540 1992.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1751.540 2172.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1751.540 2352.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1751.540 2532.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2301.540 372.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2301.540 552.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2301.540 732.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 2301.540 912.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 2301.540 1092.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 2301.540 1272.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 2301.540 1452.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 2301.540 1632.070 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -9.470 1812.070 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 2301.540 1992.070 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2785.000 372.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2785.000 552.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2785.000 732.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 2785.000 912.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 2785.000 1092.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 2785.000 1272.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 2301.540 2352.070 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 2301.540 2532.070 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -9.470 192.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 3200.495 372.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 3200.495 552.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 3200.495 732.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 3200.495 912.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 3200.495 1092.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 3200.495 1272.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 2785.000 1452.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 3240.165 1632.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 3240.165 1812.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 3240.165 1992.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 2301.540 2172.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 3185.000 2352.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 3185.000 2532.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -9.470 2712.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -9.470 2892.070 3529.150 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 114.950 3517.600 115.510 3524.800 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 32.930 2944.050 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 212.930 2944.050 216.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 392.930 2944.050 396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 572.930 2944.050 576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 752.930 2944.050 756.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 932.930 2944.050 936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1112.930 2944.050 1116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1472.930 2944.050 1476.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1652.930 2944.050 1656.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2012.930 2944.050 2016.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2192.930 2944.050 2196.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2372.930 2944.050 2376.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 387.570 2827.630 1290.670 2830.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2912.930 2944.050 2916.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3092.930 2944.050 3096.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3272.930 2944.050 3276.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3452.930 2944.050 3456.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 -19.070 390.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 -19.070 570.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 -19.070 750.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 -19.070 930.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 -19.070 1110.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 -19.070 1290.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 -19.070 1470.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 -19.070 1650.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 -19.070 2010.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 -19.070 2190.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 -19.070 2370.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 -19.070 2550.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 651.540 390.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 651.540 570.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 651.540 750.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 651.540 930.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 651.540 1110.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 651.540 1290.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 651.540 1470.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 651.540 1650.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 651.540 2010.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 651.540 2190.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 651.540 2370.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 651.540 2550.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 1201.540 390.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 1201.540 570.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 1201.540 750.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 1201.540 930.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 1201.540 1110.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 1201.540 1290.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 1201.540 1470.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 1201.540 1650.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 1201.540 2010.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 1201.540 2190.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 1201.540 2370.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 1201.540 2550.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 1751.540 390.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 1751.540 570.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 1751.540 750.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 1751.540 930.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 1751.540 1110.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 1751.540 1290.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 1751.540 1470.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 1751.540 1650.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 1751.540 2010.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 1751.540 2190.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 1751.540 2370.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 1751.540 2550.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 2301.540 390.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 2301.540 570.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 2301.540 750.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 2301.540 930.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 2301.540 1110.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 2301.540 1290.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 2301.540 1470.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 2301.540 1650.670 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 -19.070 1830.670 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 2301.540 2010.670 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 2785.000 390.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 2785.000 570.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 2785.000 750.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 2785.000 930.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 2785.000 1110.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 2785.000 1290.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 2301.540 2370.670 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 2301.540 2550.670 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 -19.070 210.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 3200.495 390.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 3200.495 570.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 3200.495 750.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 3200.495 930.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 3200.495 1110.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 3200.495 1290.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 2785.000 1470.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 3240.165 1650.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 3240.165 1830.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 3240.165 2010.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 2301.540 2190.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 3185.000 2370.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 3185.000 2550.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 -19.070 2730.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.570 -19.070 2910.670 3538.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 51.530 2953.650 54.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 231.530 2953.650 234.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 411.530 2953.650 414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 591.530 2953.650 594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 406.170 686.230 2569.270 689.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 771.530 2953.650 774.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 951.530 2953.650 954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1131.530 2953.650 1134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1491.530 2953.650 1494.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1671.530 2953.650 1674.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2031.530 2953.650 2034.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2211.530 2953.650 2214.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2391.530 2953.650 2394.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 406.170 2836.830 1309.270 2839.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2931.530 2953.650 2934.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3111.530 2953.650 3114.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3291.530 2953.650 3294.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3471.530 2953.650 3474.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 -28.670 409.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 -28.670 589.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 -28.670 769.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 -28.670 949.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 -28.670 1129.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 -28.670 1309.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 -28.670 1489.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 -28.670 1669.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 -28.670 2029.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 -28.670 2209.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 -28.670 2389.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 -28.670 2569.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 651.540 409.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 651.540 589.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 651.540 769.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 651.540 949.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 651.540 1129.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 651.540 1309.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 651.540 1489.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 651.540 1669.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 651.540 2029.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 651.540 2209.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 651.540 2389.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 651.540 2569.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 1201.540 409.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 1201.540 589.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 1201.540 769.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 1201.540 949.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 1201.540 1129.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 1201.540 1309.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 1201.540 1489.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 1201.540 1669.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 1201.540 2029.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 1201.540 2209.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 1201.540 2389.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 1201.540 2569.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 1751.540 409.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 1751.540 589.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 1751.540 769.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 1751.540 949.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 1751.540 1129.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 1751.540 1309.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 1751.540 1489.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 1751.540 1669.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 1751.540 2029.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 1751.540 2209.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 1751.540 2389.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 1751.540 2569.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 2301.540 409.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 2301.540 589.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 2301.540 769.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 2301.540 949.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 2301.540 1129.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 2301.540 1309.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 2301.540 1489.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 2301.540 1669.270 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 -28.670 1849.270 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 2301.540 2029.270 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 2785.000 409.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 2785.000 589.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 2785.000 769.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 2785.000 949.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 2785.000 1129.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 2785.000 1309.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 2301.540 2389.270 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 -28.670 229.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 3200.495 409.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 3200.495 589.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 3200.495 769.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 3200.495 949.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 3200.495 1129.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 3200.495 1309.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 2785.000 1489.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 3240.165 1669.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 3240.165 1849.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 3240.165 2029.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 2301.540 2209.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 3185.000 2389.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 2301.540 2569.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 -28.670 2749.270 3548.350 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3422.860 2924.800 3424.060 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 250.130 2963.250 253.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 430.130 2963.250 433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 610.130 2963.250 613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 424.770 704.830 2587.870 707.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 790.130 2963.250 793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.130 2963.250 973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 424.770 1244.830 2587.870 1247.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 424.770 1784.830 2587.870 1787.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 424.770 2855.430 1327.870 2858.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 -38.270 427.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 -38.270 607.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 -38.270 787.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 -38.270 967.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 -38.270 1147.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 -38.270 1327.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 -38.270 1507.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 -38.270 1687.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 -38.270 2047.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 -38.270 2227.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 -38.270 2407.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 -38.270 2587.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 651.540 427.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 651.540 607.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 651.540 787.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 651.540 967.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 651.540 1147.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 651.540 1327.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 651.540 1507.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 651.540 1687.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 651.540 2047.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 651.540 2227.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 651.540 2407.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 651.540 2587.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 1201.540 427.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 1201.540 607.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 1201.540 787.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 1201.540 967.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 1201.540 1147.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 1201.540 1327.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 1201.540 1507.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 1201.540 1687.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 1201.540 2047.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 1201.540 2227.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 1201.540 2407.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 1201.540 2587.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 1751.540 427.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 1751.540 607.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 1751.540 787.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 1751.540 967.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 1751.540 1147.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 1751.540 1327.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 1751.540 1507.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 1751.540 1687.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 1751.540 2047.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 1751.540 2227.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 1751.540 2407.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 1751.540 2587.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 2301.540 427.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 2301.540 607.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 2301.540 787.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 2301.540 967.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 2301.540 1147.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 2301.540 1327.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 2301.540 1507.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 2301.540 1687.870 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 -38.270 1867.870 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 2301.540 2047.870 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 2785.000 427.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 2785.000 607.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 2785.000 787.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 2785.000 967.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 2785.000 1147.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 2785.000 1327.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 2301.540 2407.870 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 -38.270 247.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 3200.495 427.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 3200.495 607.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 3200.495 787.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 3200.495 967.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 3200.495 1147.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 3200.495 1327.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 2785.000 1507.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 3240.165 1687.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 3240.165 1867.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 3240.165 2047.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 2301.540 2227.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 3185.000 2407.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 2301.540 2587.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 -38.270 2767.870 3557.950 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 38.130 3517.600 38.690 3524.800 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 141.530 2953.650 144.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 321.530 2953.650 324.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 501.530 2953.650 504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 681.530 2953.650 684.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 861.530 2953.650 864.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1041.530 2953.650 1044.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1221.530 2953.650 1224.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1581.530 2953.650 1584.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1761.530 2953.650 1764.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2121.530 2953.650 2124.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 316.170 2386.830 1399.270 2389.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2481.530 2953.650 2484.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2661.530 2953.650 2664.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2841.530 2953.650 2844.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3021.530 2953.650 3024.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3381.530 2953.650 3384.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 -28.670 319.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 -28.670 499.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 -28.670 679.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 -28.670 859.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 -28.670 1219.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 -28.670 1399.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 -28.670 1579.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 -28.670 1759.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 -28.670 1939.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 -28.670 2119.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 -28.670 2299.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 -28.670 2479.270 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 651.540 319.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 651.540 499.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 651.540 679.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 651.540 859.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 651.540 1219.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 651.540 1399.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 651.540 1579.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 651.540 1759.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 651.540 1939.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 651.540 2119.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 651.540 2299.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 651.540 2479.270 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 1201.540 319.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 1201.540 499.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 1201.540 679.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 1201.540 859.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 1201.540 1219.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 1201.540 1399.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 1201.540 1579.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 1201.540 1759.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 1201.540 1939.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 1201.540 2119.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 1201.540 2299.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 1201.540 2479.270 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 1751.540 319.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 1751.540 499.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 1751.540 679.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 1751.540 859.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 1751.540 1219.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 1751.540 1399.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 1751.540 1579.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 1751.540 1759.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 1751.540 1939.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 1751.540 2119.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 1751.540 2299.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 1751.540 2479.270 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 2301.540 319.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 2301.540 499.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 2301.540 679.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 2301.540 859.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1036.170 -28.670 1039.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 2301.540 1219.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 2301.540 1399.270 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 2301.540 1759.270 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 2301.540 1939.270 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 2301.540 2119.270 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 2785.000 319.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 2785.000 499.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 2785.000 859.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 2785.000 1219.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 2785.000 1399.270 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 2301.540 2299.270 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 2301.540 2479.270 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.170 -28.670 139.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 3200.495 319.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 3200.495 499.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 2785.000 679.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 3200.495 859.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1036.170 2785.000 1039.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 3200.495 1219.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 3200.495 1399.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 2301.540 1579.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 3240.165 1759.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 3240.165 1939.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 3240.165 2119.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 3185.000 2299.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 3185.000 2479.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.170 -28.670 2659.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.170 -28.670 2839.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 160.130 2963.250 163.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 340.130 2963.250 343.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 520.130 2963.250 523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 700.130 2963.250 703.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 880.130 2963.250 883.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1060.130 2963.250 1063.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1240.130 2963.250 1243.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1600.130 2963.250 1603.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1780.130 2963.250 1783.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2140.130 2963.250 2143.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2500.130 2963.250 2503.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2680.130 2963.250 2683.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2860.130 2963.250 2863.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3040.130 2963.250 3043.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3400.130 2963.250 3403.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 -38.270 337.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 -38.270 517.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 -38.270 697.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 -38.270 877.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 -38.270 1237.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 -38.270 1417.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 -38.270 1597.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 -38.270 1777.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 -38.270 1957.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 -38.270 2137.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 -38.270 2317.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 -38.270 2497.870 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 651.540 337.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 651.540 517.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 651.540 697.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 651.540 877.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 651.540 1237.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 651.540 1417.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 651.540 1597.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 651.540 1777.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 651.540 1957.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 651.540 2137.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 651.540 2317.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 651.540 2497.870 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 1201.540 337.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 1201.540 517.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 1201.540 697.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 1201.540 877.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 1201.540 1237.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 1201.540 1417.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 1201.540 1597.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 1201.540 1777.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 1201.540 1957.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 1201.540 2137.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 1201.540 2317.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 1201.540 2497.870 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 1751.540 337.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 1751.540 517.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 1751.540 697.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 1751.540 877.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 1751.540 1237.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 1751.540 1417.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 1751.540 1597.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 1751.540 1777.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 1751.540 1957.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 1751.540 2137.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 1751.540 2317.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 1751.540 2497.870 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 2301.540 337.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 2301.540 517.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 2301.540 697.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 2301.540 877.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.770 -38.270 1057.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 2301.540 1237.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 2301.540 1417.870 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 2301.540 1597.870 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 2301.540 1777.870 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 2301.540 1957.870 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 2301.540 2137.870 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 2785.000 337.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 2785.000 517.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 2785.000 697.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 2785.000 877.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 2785.000 1237.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 2785.000 1417.870 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 2301.540 2317.870 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 2301.540 2497.870 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.770 -38.270 157.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 3200.495 337.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 3200.495 517.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 3200.495 697.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 3200.495 877.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.770 2785.000 1057.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 3200.495 1237.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 3200.495 1417.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 3240.165 1597.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 3240.165 1777.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 3240.165 1957.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 3240.165 2137.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 3185.000 2317.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 3185.000 2497.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.770 -38.270 2677.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.770 -38.270 2857.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3486.780 2924.800 3487.980 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 104.330 2934.450 107.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 284.330 2934.450 287.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 464.330 2934.450 467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 644.330 2934.450 647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 458.970 729.630 2442.070 732.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 824.330 2934.450 827.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1004.330 2934.450 1007.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1184.330 2934.450 1187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 458.970 1269.630 2442.070 1272.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1364.330 2934.450 1367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1544.330 2934.450 1547.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1724.330 2934.450 1727.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 458.970 1809.630 2442.070 1812.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1904.330 2934.450 1907.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2084.330 2934.450 2087.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2264.330 2934.450 2267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2444.330 2934.450 2447.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2624.330 2934.450 2627.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2804.330 2934.450 2807.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2984.330 2934.450 2987.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3164.330 2934.450 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3344.330 2934.450 3347.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 -9.470 462.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 -9.470 642.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 -9.470 822.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 -9.470 1182.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 -9.470 1362.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 -9.470 1542.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 -9.470 1722.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 -9.470 1902.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 -9.470 2082.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -9.470 2262.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 -9.470 2442.070 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 651.540 462.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 651.540 642.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 651.540 822.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 651.540 1182.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 651.540 1362.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 651.540 1542.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 651.540 1722.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 651.540 1902.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 651.540 2082.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 651.540 2262.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 651.540 2442.070 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1201.540 462.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1201.540 642.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 1201.540 822.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 1201.540 1182.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 1201.540 1362.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 1201.540 1542.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 1201.540 1722.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 1201.540 1902.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 1201.540 2082.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1201.540 2262.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1201.540 2442.070 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1751.540 462.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1751.540 642.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 1751.540 822.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 1751.540 1182.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 1751.540 1362.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 1751.540 1542.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 1751.540 1722.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 1751.540 1902.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 1751.540 2082.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1751.540 2262.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1751.540 2442.070 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2301.540 462.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2301.540 642.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 2301.540 822.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 -9.470 1002.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 2301.540 1182.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 2301.540 1362.070 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 2301.540 1722.070 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 2301.540 1902.070 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 2301.540 2082.070 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2785.000 462.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 2785.000 822.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 2785.000 1002.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 2785.000 1182.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 2785.000 1362.070 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 2301.540 2442.070 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 -9.470 102.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 -9.470 282.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 3200.495 462.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2785.000 642.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 3200.495 822.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 3200.495 1002.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 3200.495 1182.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 3200.495 1362.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 2301.540 1542.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 3240.165 1722.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 3240.165 1902.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 3240.165 2082.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2301.540 2262.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 3185.000 2442.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 -9.470 2622.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 -9.470 2802.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -4.800 93.580 2.400 94.780 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 122.930 2944.050 126.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 302.930 2944.050 306.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 482.930 2944.050 486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 662.930 2944.050 666.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 842.930 2944.050 846.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1022.930 2944.050 1026.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1202.930 2944.050 1206.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1562.930 2944.050 1566.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1742.930 2944.050 1746.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 297.570 1828.230 2460.670 1831.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2102.930 2944.050 2106.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 297.570 2377.630 1380.670 2380.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2462.930 2944.050 2466.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2642.930 2944.050 2646.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2822.930 2944.050 2826.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3002.930 2944.050 3006.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3362.930 2944.050 3366.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 -19.070 300.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 -19.070 480.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 -19.070 660.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 -19.070 840.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 -19.070 1200.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 -19.070 1380.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 -19.070 1560.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 -19.070 1740.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 -19.070 1920.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 -19.070 2100.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 -19.070 2280.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 -19.070 2460.670 215.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 651.540 300.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 651.540 480.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 651.540 660.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 651.540 840.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 651.540 1200.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 651.540 1380.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 651.540 1560.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 651.540 1740.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 651.540 1920.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 651.540 2100.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 651.540 2280.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 651.540 2460.670 765.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 1201.540 300.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 1201.540 480.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 1201.540 660.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 1201.540 840.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 1201.540 1200.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 1201.540 1380.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 1201.540 1560.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 1201.540 1740.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 1201.540 1920.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 1201.540 2100.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 1201.540 2280.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 1201.540 2460.670 1315.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 1751.540 300.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 1751.540 480.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 1751.540 660.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 1751.540 840.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 1751.540 1200.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 1751.540 1380.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 1751.540 1560.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 1751.540 1740.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 1751.540 1920.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 1751.540 2100.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 1751.540 2280.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 1751.540 2460.670 1865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 2301.540 300.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 2301.540 480.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 2301.540 660.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 2301.540 840.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.570 -19.070 1020.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 2301.540 1200.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 2301.540 1380.670 2465.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 2301.540 1740.670 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 2301.540 1920.670 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 2301.540 2100.670 2665.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 2785.000 300.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 2785.000 480.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 2785.000 840.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 2785.000 1200.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 2785.000 1380.670 2865.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 2301.540 2460.670 2915.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.570 -19.070 120.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 3200.495 300.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 3200.495 480.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 2785.000 660.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 3200.495 840.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.570 2785.000 1020.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 3200.495 1200.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 3200.495 1380.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 2301.540 1560.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 3240.165 1740.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 3240.165 1920.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 3240.165 2100.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 2301.540 2280.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 3185.000 2460.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.570 -19.070 2640.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.570 -19.070 2820.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.020 2.400 32.220 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.670 -4.800 38.230 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.770 -4.800 238.330 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.710 -4.800 256.270 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.190 -4.800 273.750 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.130 -4.800 291.690 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.610 -4.800 309.170 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.090 -4.800 326.650 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.030 -4.800 344.590 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.510 -4.800 362.070 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.450 -4.800 380.010 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.930 -4.800 397.490 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 -4.800 61.690 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.410 -4.800 414.970 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.350 -4.800 432.910 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.830 -4.800 450.390 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.770 -4.800 468.330 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.250 -4.800 485.810 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.730 -4.800 503.290 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.670 -4.800 521.230 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.150 -4.800 538.710 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.090 -4.800 556.650 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.510 -4.800 109.070 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 -4.800 132.530 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 -4.800 150.010 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 -4.800 167.950 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.870 -4.800 185.430 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.810 -4.800 203.370 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.290 -4.800 220.850 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.750 -4.800 244.310 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.690 -4.800 262.250 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.170 -4.800 279.730 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.650 -4.800 297.210 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.590 -4.800 315.150 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.070 -4.800 332.630 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.010 -4.800 350.570 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.490 -4.800 368.050 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.970 -4.800 385.530 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.910 -4.800 403.470 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 -4.800 67.670 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.390 -4.800 420.950 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.330 -4.800 438.890 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.810 -4.800 456.370 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.290 -4.800 473.850 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.230 -4.800 491.790 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.710 -4.800 509.270 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.650 -4.800 527.210 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.130 -4.800 544.690 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.570 -4.800 91.130 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.490 -4.800 115.050 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 -4.800 138.510 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 -4.800 155.990 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.370 -4.800 173.930 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.850 -4.800 191.410 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.330 -4.800 208.890 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.270 -4.800 226.830 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.730 -4.800 250.290 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.210 -4.800 267.770 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.150 -4.800 285.710 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 -4.800 303.190 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.570 -4.800 321.130 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.050 -4.800 338.610 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.530 -4.800 356.090 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.470 -4.800 374.030 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.950 -4.800 391.510 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.890 -4.800 409.450 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.090 -4.800 73.650 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.370 -4.800 426.930 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.850 -4.800 444.410 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.790 -4.800 462.350 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.270 -4.800 479.830 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.210 -4.800 497.770 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.690 -4.800 515.250 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.170 -4.800 532.730 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.110 -4.800 550.670 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 -4.800 97.110 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.490 -4.800 621.050 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.010 -4.800 120.570 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.930 -4.800 144.490 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.410 -4.800 161.970 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.890 -4.800 179.450 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.830 -4.800 197.390 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.310 -4.800 214.870 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.250 -4.800 232.810 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 -4.800 79.630 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.530 -4.800 103.090 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 -4.800 126.550 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.690 -4.800 32.250 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 305.520 2485.795 2544.260 3219.085 ;
      LAYER met1 ;
        RECT 2.830 17.040 2902.530 3505.020 ;
      LAYER met2 ;
        RECT 2.860 3517.320 37.850 3518.050 ;
        RECT 38.970 3517.320 114.670 3518.050 ;
        RECT 115.790 3517.320 191.490 3518.050 ;
        RECT 192.610 3517.320 268.310 3518.050 ;
        RECT 269.430 3517.320 345.130 3518.050 ;
        RECT 346.250 3517.320 421.950 3518.050 ;
        RECT 423.070 3517.320 498.770 3518.050 ;
        RECT 499.890 3517.320 575.590 3518.050 ;
        RECT 576.710 3517.320 652.410 3518.050 ;
        RECT 653.530 3517.320 729.230 3518.050 ;
        RECT 730.350 3517.320 806.050 3518.050 ;
        RECT 807.170 3517.320 882.870 3518.050 ;
        RECT 883.990 3517.320 959.690 3518.050 ;
        RECT 960.810 3517.320 1036.510 3518.050 ;
        RECT 1037.630 3517.320 1113.330 3518.050 ;
        RECT 1114.450 3517.320 1190.150 3518.050 ;
        RECT 1191.270 3517.320 1266.970 3518.050 ;
        RECT 1268.090 3517.320 1343.790 3518.050 ;
        RECT 1344.910 3517.320 1420.610 3518.050 ;
        RECT 1421.730 3517.320 1497.890 3518.050 ;
        RECT 1499.010 3517.320 1574.710 3518.050 ;
        RECT 1575.830 3517.320 1651.530 3518.050 ;
        RECT 1652.650 3517.320 1728.350 3518.050 ;
        RECT 1729.470 3517.320 1805.170 3518.050 ;
        RECT 1806.290 3517.320 1881.990 3518.050 ;
        RECT 1883.110 3517.320 1958.810 3518.050 ;
        RECT 1959.930 3517.320 2035.630 3518.050 ;
        RECT 2036.750 3517.320 2112.450 3518.050 ;
        RECT 2113.570 3517.320 2189.270 3518.050 ;
        RECT 2190.390 3517.320 2266.090 3518.050 ;
        RECT 2267.210 3517.320 2342.910 3518.050 ;
        RECT 2344.030 3517.320 2419.730 3518.050 ;
        RECT 2420.850 3517.320 2496.550 3518.050 ;
        RECT 2497.670 3517.320 2573.370 3518.050 ;
        RECT 2574.490 3517.320 2650.190 3518.050 ;
        RECT 2651.310 3517.320 2727.010 3518.050 ;
        RECT 2728.130 3517.320 2803.830 3518.050 ;
        RECT 2804.950 3517.320 2880.650 3518.050 ;
        RECT 2881.770 3517.320 2904.810 3518.050 ;
        RECT 2.860 2.680 2904.810 3517.320 ;
        RECT 3.550 2.400 7.950 2.680 ;
        RECT 9.070 2.400 13.930 2.680 ;
        RECT 15.050 2.400 19.910 2.680 ;
        RECT 21.030 2.400 25.890 2.680 ;
        RECT 27.010 2.400 31.410 2.680 ;
        RECT 32.530 2.400 37.390 2.680 ;
        RECT 38.510 2.400 43.370 2.680 ;
        RECT 44.490 2.400 49.350 2.680 ;
        RECT 50.470 2.400 55.330 2.680 ;
        RECT 56.450 2.400 60.850 2.680 ;
        RECT 61.970 2.400 66.830 2.680 ;
        RECT 67.950 2.400 72.810 2.680 ;
        RECT 73.930 2.400 78.790 2.680 ;
        RECT 79.910 2.400 84.770 2.680 ;
        RECT 85.890 2.400 90.290 2.680 ;
        RECT 91.410 2.400 96.270 2.680 ;
        RECT 97.390 2.400 102.250 2.680 ;
        RECT 103.370 2.400 108.230 2.680 ;
        RECT 109.350 2.400 114.210 2.680 ;
        RECT 115.330 2.400 119.730 2.680 ;
        RECT 120.850 2.400 125.710 2.680 ;
        RECT 126.830 2.400 131.690 2.680 ;
        RECT 132.810 2.400 137.670 2.680 ;
        RECT 138.790 2.400 143.650 2.680 ;
        RECT 144.770 2.400 149.170 2.680 ;
        RECT 150.290 2.400 155.150 2.680 ;
        RECT 156.270 2.400 161.130 2.680 ;
        RECT 162.250 2.400 167.110 2.680 ;
        RECT 168.230 2.400 173.090 2.680 ;
        RECT 174.210 2.400 178.610 2.680 ;
        RECT 179.730 2.400 184.590 2.680 ;
        RECT 185.710 2.400 190.570 2.680 ;
        RECT 191.690 2.400 196.550 2.680 ;
        RECT 197.670 2.400 202.530 2.680 ;
        RECT 203.650 2.400 208.050 2.680 ;
        RECT 209.170 2.400 214.030 2.680 ;
        RECT 215.150 2.400 220.010 2.680 ;
        RECT 221.130 2.400 225.990 2.680 ;
        RECT 227.110 2.400 231.970 2.680 ;
        RECT 233.090 2.400 237.490 2.680 ;
        RECT 238.610 2.400 243.470 2.680 ;
        RECT 244.590 2.400 249.450 2.680 ;
        RECT 250.570 2.400 255.430 2.680 ;
        RECT 256.550 2.400 261.410 2.680 ;
        RECT 262.530 2.400 266.930 2.680 ;
        RECT 268.050 2.400 272.910 2.680 ;
        RECT 274.030 2.400 278.890 2.680 ;
        RECT 280.010 2.400 284.870 2.680 ;
        RECT 285.990 2.400 290.850 2.680 ;
        RECT 291.970 2.400 296.370 2.680 ;
        RECT 297.490 2.400 302.350 2.680 ;
        RECT 303.470 2.400 308.330 2.680 ;
        RECT 309.450 2.400 314.310 2.680 ;
        RECT 315.430 2.400 320.290 2.680 ;
        RECT 321.410 2.400 325.810 2.680 ;
        RECT 326.930 2.400 331.790 2.680 ;
        RECT 332.910 2.400 337.770 2.680 ;
        RECT 338.890 2.400 343.750 2.680 ;
        RECT 344.870 2.400 349.730 2.680 ;
        RECT 350.850 2.400 355.250 2.680 ;
        RECT 356.370 2.400 361.230 2.680 ;
        RECT 362.350 2.400 367.210 2.680 ;
        RECT 368.330 2.400 373.190 2.680 ;
        RECT 374.310 2.400 379.170 2.680 ;
        RECT 380.290 2.400 384.690 2.680 ;
        RECT 385.810 2.400 390.670 2.680 ;
        RECT 391.790 2.400 396.650 2.680 ;
        RECT 397.770 2.400 402.630 2.680 ;
        RECT 403.750 2.400 408.610 2.680 ;
        RECT 409.730 2.400 414.130 2.680 ;
        RECT 415.250 2.400 420.110 2.680 ;
        RECT 421.230 2.400 426.090 2.680 ;
        RECT 427.210 2.400 432.070 2.680 ;
        RECT 433.190 2.400 438.050 2.680 ;
        RECT 439.170 2.400 443.570 2.680 ;
        RECT 444.690 2.400 449.550 2.680 ;
        RECT 450.670 2.400 455.530 2.680 ;
        RECT 456.650 2.400 461.510 2.680 ;
        RECT 462.630 2.400 467.490 2.680 ;
        RECT 468.610 2.400 473.010 2.680 ;
        RECT 474.130 2.400 478.990 2.680 ;
        RECT 480.110 2.400 484.970 2.680 ;
        RECT 486.090 2.400 490.950 2.680 ;
        RECT 492.070 2.400 496.930 2.680 ;
        RECT 498.050 2.400 502.450 2.680 ;
        RECT 503.570 2.400 508.430 2.680 ;
        RECT 509.550 2.400 514.410 2.680 ;
        RECT 515.530 2.400 520.390 2.680 ;
        RECT 521.510 2.400 526.370 2.680 ;
        RECT 527.490 2.400 531.890 2.680 ;
        RECT 533.010 2.400 537.870 2.680 ;
        RECT 538.990 2.400 543.850 2.680 ;
        RECT 544.970 2.400 549.830 2.680 ;
        RECT 550.950 2.400 555.810 2.680 ;
        RECT 556.930 2.400 561.330 2.680 ;
        RECT 562.450 2.400 567.310 2.680 ;
        RECT 568.430 2.400 573.290 2.680 ;
        RECT 574.410 2.400 579.270 2.680 ;
        RECT 580.390 2.400 585.250 2.680 ;
        RECT 586.370 2.400 590.770 2.680 ;
        RECT 591.890 2.400 596.750 2.680 ;
        RECT 597.870 2.400 602.730 2.680 ;
        RECT 603.850 2.400 608.710 2.680 ;
        RECT 609.830 2.400 614.690 2.680 ;
        RECT 615.810 2.400 620.210 2.680 ;
        RECT 621.330 2.400 626.190 2.680 ;
        RECT 627.310 2.400 632.170 2.680 ;
        RECT 633.290 2.400 638.150 2.680 ;
        RECT 639.270 2.400 644.130 2.680 ;
        RECT 645.250 2.400 649.650 2.680 ;
        RECT 650.770 2.400 655.630 2.680 ;
        RECT 656.750 2.400 661.610 2.680 ;
        RECT 662.730 2.400 667.590 2.680 ;
        RECT 668.710 2.400 673.570 2.680 ;
        RECT 674.690 2.400 679.090 2.680 ;
        RECT 680.210 2.400 685.070 2.680 ;
        RECT 686.190 2.400 691.050 2.680 ;
        RECT 692.170 2.400 697.030 2.680 ;
        RECT 698.150 2.400 703.010 2.680 ;
        RECT 704.130 2.400 708.530 2.680 ;
        RECT 709.650 2.400 714.510 2.680 ;
        RECT 715.630 2.400 720.490 2.680 ;
        RECT 721.610 2.400 726.470 2.680 ;
        RECT 727.590 2.400 732.450 2.680 ;
        RECT 733.570 2.400 737.970 2.680 ;
        RECT 739.090 2.400 743.950 2.680 ;
        RECT 745.070 2.400 749.930 2.680 ;
        RECT 751.050 2.400 755.910 2.680 ;
        RECT 757.030 2.400 761.430 2.680 ;
        RECT 762.550 2.400 767.410 2.680 ;
        RECT 768.530 2.400 773.390 2.680 ;
        RECT 774.510 2.400 779.370 2.680 ;
        RECT 780.490 2.400 785.350 2.680 ;
        RECT 786.470 2.400 790.870 2.680 ;
        RECT 791.990 2.400 796.850 2.680 ;
        RECT 797.970 2.400 802.830 2.680 ;
        RECT 803.950 2.400 808.810 2.680 ;
        RECT 809.930 2.400 814.790 2.680 ;
        RECT 815.910 2.400 820.310 2.680 ;
        RECT 821.430 2.400 826.290 2.680 ;
        RECT 827.410 2.400 832.270 2.680 ;
        RECT 833.390 2.400 838.250 2.680 ;
        RECT 839.370 2.400 844.230 2.680 ;
        RECT 845.350 2.400 849.750 2.680 ;
        RECT 850.870 2.400 855.730 2.680 ;
        RECT 856.850 2.400 861.710 2.680 ;
        RECT 862.830 2.400 867.690 2.680 ;
        RECT 868.810 2.400 873.670 2.680 ;
        RECT 874.790 2.400 879.190 2.680 ;
        RECT 880.310 2.400 885.170 2.680 ;
        RECT 886.290 2.400 891.150 2.680 ;
        RECT 892.270 2.400 897.130 2.680 ;
        RECT 898.250 2.400 903.110 2.680 ;
        RECT 904.230 2.400 908.630 2.680 ;
        RECT 909.750 2.400 914.610 2.680 ;
        RECT 915.730 2.400 920.590 2.680 ;
        RECT 921.710 2.400 926.570 2.680 ;
        RECT 927.690 2.400 932.550 2.680 ;
        RECT 933.670 2.400 938.070 2.680 ;
        RECT 939.190 2.400 944.050 2.680 ;
        RECT 945.170 2.400 950.030 2.680 ;
        RECT 951.150 2.400 956.010 2.680 ;
        RECT 957.130 2.400 961.990 2.680 ;
        RECT 963.110 2.400 967.510 2.680 ;
        RECT 968.630 2.400 973.490 2.680 ;
        RECT 974.610 2.400 979.470 2.680 ;
        RECT 980.590 2.400 985.450 2.680 ;
        RECT 986.570 2.400 991.430 2.680 ;
        RECT 992.550 2.400 996.950 2.680 ;
        RECT 998.070 2.400 1002.930 2.680 ;
        RECT 1004.050 2.400 1008.910 2.680 ;
        RECT 1010.030 2.400 1014.890 2.680 ;
        RECT 1016.010 2.400 1020.870 2.680 ;
        RECT 1021.990 2.400 1026.390 2.680 ;
        RECT 1027.510 2.400 1032.370 2.680 ;
        RECT 1033.490 2.400 1038.350 2.680 ;
        RECT 1039.470 2.400 1044.330 2.680 ;
        RECT 1045.450 2.400 1050.310 2.680 ;
        RECT 1051.430 2.400 1055.830 2.680 ;
        RECT 1056.950 2.400 1061.810 2.680 ;
        RECT 1062.930 2.400 1067.790 2.680 ;
        RECT 1068.910 2.400 1073.770 2.680 ;
        RECT 1074.890 2.400 1079.750 2.680 ;
        RECT 1080.870 2.400 1085.270 2.680 ;
        RECT 1086.390 2.400 1091.250 2.680 ;
        RECT 1092.370 2.400 1097.230 2.680 ;
        RECT 1098.350 2.400 1103.210 2.680 ;
        RECT 1104.330 2.400 1109.190 2.680 ;
        RECT 1110.310 2.400 1114.710 2.680 ;
        RECT 1115.830 2.400 1120.690 2.680 ;
        RECT 1121.810 2.400 1126.670 2.680 ;
        RECT 1127.790 2.400 1132.650 2.680 ;
        RECT 1133.770 2.400 1138.630 2.680 ;
        RECT 1139.750 2.400 1144.150 2.680 ;
        RECT 1145.270 2.400 1150.130 2.680 ;
        RECT 1151.250 2.400 1156.110 2.680 ;
        RECT 1157.230 2.400 1162.090 2.680 ;
        RECT 1163.210 2.400 1168.070 2.680 ;
        RECT 1169.190 2.400 1173.590 2.680 ;
        RECT 1174.710 2.400 1179.570 2.680 ;
        RECT 1180.690 2.400 1185.550 2.680 ;
        RECT 1186.670 2.400 1191.530 2.680 ;
        RECT 1192.650 2.400 1197.510 2.680 ;
        RECT 1198.630 2.400 1203.030 2.680 ;
        RECT 1204.150 2.400 1209.010 2.680 ;
        RECT 1210.130 2.400 1214.990 2.680 ;
        RECT 1216.110 2.400 1220.970 2.680 ;
        RECT 1222.090 2.400 1226.950 2.680 ;
        RECT 1228.070 2.400 1232.470 2.680 ;
        RECT 1233.590 2.400 1238.450 2.680 ;
        RECT 1239.570 2.400 1244.430 2.680 ;
        RECT 1245.550 2.400 1250.410 2.680 ;
        RECT 1251.530 2.400 1256.390 2.680 ;
        RECT 1257.510 2.400 1261.910 2.680 ;
        RECT 1263.030 2.400 1267.890 2.680 ;
        RECT 1269.010 2.400 1273.870 2.680 ;
        RECT 1274.990 2.400 1279.850 2.680 ;
        RECT 1280.970 2.400 1285.830 2.680 ;
        RECT 1286.950 2.400 1291.350 2.680 ;
        RECT 1292.470 2.400 1297.330 2.680 ;
        RECT 1298.450 2.400 1303.310 2.680 ;
        RECT 1304.430 2.400 1309.290 2.680 ;
        RECT 1310.410 2.400 1315.270 2.680 ;
        RECT 1316.390 2.400 1320.790 2.680 ;
        RECT 1321.910 2.400 1326.770 2.680 ;
        RECT 1327.890 2.400 1332.750 2.680 ;
        RECT 1333.870 2.400 1338.730 2.680 ;
        RECT 1339.850 2.400 1344.710 2.680 ;
        RECT 1345.830 2.400 1350.230 2.680 ;
        RECT 1351.350 2.400 1356.210 2.680 ;
        RECT 1357.330 2.400 1362.190 2.680 ;
        RECT 1363.310 2.400 1368.170 2.680 ;
        RECT 1369.290 2.400 1374.150 2.680 ;
        RECT 1375.270 2.400 1379.670 2.680 ;
        RECT 1380.790 2.400 1385.650 2.680 ;
        RECT 1386.770 2.400 1391.630 2.680 ;
        RECT 1392.750 2.400 1397.610 2.680 ;
        RECT 1398.730 2.400 1403.590 2.680 ;
        RECT 1404.710 2.400 1409.110 2.680 ;
        RECT 1410.230 2.400 1415.090 2.680 ;
        RECT 1416.210 2.400 1421.070 2.680 ;
        RECT 1422.190 2.400 1427.050 2.680 ;
        RECT 1428.170 2.400 1433.030 2.680 ;
        RECT 1434.150 2.400 1438.550 2.680 ;
        RECT 1439.670 2.400 1444.530 2.680 ;
        RECT 1445.650 2.400 1450.510 2.680 ;
        RECT 1451.630 2.400 1456.490 2.680 ;
        RECT 1457.610 2.400 1462.470 2.680 ;
        RECT 1463.590 2.400 1467.990 2.680 ;
        RECT 1469.110 2.400 1473.970 2.680 ;
        RECT 1475.090 2.400 1479.950 2.680 ;
        RECT 1481.070 2.400 1485.930 2.680 ;
        RECT 1487.050 2.400 1491.450 2.680 ;
        RECT 1492.570 2.400 1497.430 2.680 ;
        RECT 1498.550 2.400 1503.410 2.680 ;
        RECT 1504.530 2.400 1509.390 2.680 ;
        RECT 1510.510 2.400 1515.370 2.680 ;
        RECT 1516.490 2.400 1520.890 2.680 ;
        RECT 1522.010 2.400 1526.870 2.680 ;
        RECT 1527.990 2.400 1532.850 2.680 ;
        RECT 1533.970 2.400 1538.830 2.680 ;
        RECT 1539.950 2.400 1544.810 2.680 ;
        RECT 1545.930 2.400 1550.330 2.680 ;
        RECT 1551.450 2.400 1556.310 2.680 ;
        RECT 1557.430 2.400 1562.290 2.680 ;
        RECT 1563.410 2.400 1568.270 2.680 ;
        RECT 1569.390 2.400 1574.250 2.680 ;
        RECT 1575.370 2.400 1579.770 2.680 ;
        RECT 1580.890 2.400 1585.750 2.680 ;
        RECT 1586.870 2.400 1591.730 2.680 ;
        RECT 1592.850 2.400 1597.710 2.680 ;
        RECT 1598.830 2.400 1603.690 2.680 ;
        RECT 1604.810 2.400 1609.210 2.680 ;
        RECT 1610.330 2.400 1615.190 2.680 ;
        RECT 1616.310 2.400 1621.170 2.680 ;
        RECT 1622.290 2.400 1627.150 2.680 ;
        RECT 1628.270 2.400 1633.130 2.680 ;
        RECT 1634.250 2.400 1638.650 2.680 ;
        RECT 1639.770 2.400 1644.630 2.680 ;
        RECT 1645.750 2.400 1650.610 2.680 ;
        RECT 1651.730 2.400 1656.590 2.680 ;
        RECT 1657.710 2.400 1662.570 2.680 ;
        RECT 1663.690 2.400 1668.090 2.680 ;
        RECT 1669.210 2.400 1674.070 2.680 ;
        RECT 1675.190 2.400 1680.050 2.680 ;
        RECT 1681.170 2.400 1686.030 2.680 ;
        RECT 1687.150 2.400 1692.010 2.680 ;
        RECT 1693.130 2.400 1697.530 2.680 ;
        RECT 1698.650 2.400 1703.510 2.680 ;
        RECT 1704.630 2.400 1709.490 2.680 ;
        RECT 1710.610 2.400 1715.470 2.680 ;
        RECT 1716.590 2.400 1721.450 2.680 ;
        RECT 1722.570 2.400 1726.970 2.680 ;
        RECT 1728.090 2.400 1732.950 2.680 ;
        RECT 1734.070 2.400 1738.930 2.680 ;
        RECT 1740.050 2.400 1744.910 2.680 ;
        RECT 1746.030 2.400 1750.890 2.680 ;
        RECT 1752.010 2.400 1756.410 2.680 ;
        RECT 1757.530 2.400 1762.390 2.680 ;
        RECT 1763.510 2.400 1768.370 2.680 ;
        RECT 1769.490 2.400 1774.350 2.680 ;
        RECT 1775.470 2.400 1780.330 2.680 ;
        RECT 1781.450 2.400 1785.850 2.680 ;
        RECT 1786.970 2.400 1791.830 2.680 ;
        RECT 1792.950 2.400 1797.810 2.680 ;
        RECT 1798.930 2.400 1803.790 2.680 ;
        RECT 1804.910 2.400 1809.770 2.680 ;
        RECT 1810.890 2.400 1815.290 2.680 ;
        RECT 1816.410 2.400 1821.270 2.680 ;
        RECT 1822.390 2.400 1827.250 2.680 ;
        RECT 1828.370 2.400 1833.230 2.680 ;
        RECT 1834.350 2.400 1839.210 2.680 ;
        RECT 1840.330 2.400 1844.730 2.680 ;
        RECT 1845.850 2.400 1850.710 2.680 ;
        RECT 1851.830 2.400 1856.690 2.680 ;
        RECT 1857.810 2.400 1862.670 2.680 ;
        RECT 1863.790 2.400 1868.650 2.680 ;
        RECT 1869.770 2.400 1874.170 2.680 ;
        RECT 1875.290 2.400 1880.150 2.680 ;
        RECT 1881.270 2.400 1886.130 2.680 ;
        RECT 1887.250 2.400 1892.110 2.680 ;
        RECT 1893.230 2.400 1898.090 2.680 ;
        RECT 1899.210 2.400 1903.610 2.680 ;
        RECT 1904.730 2.400 1909.590 2.680 ;
        RECT 1910.710 2.400 1915.570 2.680 ;
        RECT 1916.690 2.400 1921.550 2.680 ;
        RECT 1922.670 2.400 1927.530 2.680 ;
        RECT 1928.650 2.400 1933.050 2.680 ;
        RECT 1934.170 2.400 1939.030 2.680 ;
        RECT 1940.150 2.400 1945.010 2.680 ;
        RECT 1946.130 2.400 1950.990 2.680 ;
        RECT 1952.110 2.400 1956.970 2.680 ;
        RECT 1958.090 2.400 1962.490 2.680 ;
        RECT 1963.610 2.400 1968.470 2.680 ;
        RECT 1969.590 2.400 1974.450 2.680 ;
        RECT 1975.570 2.400 1980.430 2.680 ;
        RECT 1981.550 2.400 1986.410 2.680 ;
        RECT 1987.530 2.400 1991.930 2.680 ;
        RECT 1993.050 2.400 1997.910 2.680 ;
        RECT 1999.030 2.400 2003.890 2.680 ;
        RECT 2005.010 2.400 2009.870 2.680 ;
        RECT 2010.990 2.400 2015.850 2.680 ;
        RECT 2016.970 2.400 2021.370 2.680 ;
        RECT 2022.490 2.400 2027.350 2.680 ;
        RECT 2028.470 2.400 2033.330 2.680 ;
        RECT 2034.450 2.400 2039.310 2.680 ;
        RECT 2040.430 2.400 2045.290 2.680 ;
        RECT 2046.410 2.400 2050.810 2.680 ;
        RECT 2051.930 2.400 2056.790 2.680 ;
        RECT 2057.910 2.400 2062.770 2.680 ;
        RECT 2063.890 2.400 2068.750 2.680 ;
        RECT 2069.870 2.400 2074.730 2.680 ;
        RECT 2075.850 2.400 2080.250 2.680 ;
        RECT 2081.370 2.400 2086.230 2.680 ;
        RECT 2087.350 2.400 2092.210 2.680 ;
        RECT 2093.330 2.400 2098.190 2.680 ;
        RECT 2099.310 2.400 2104.170 2.680 ;
        RECT 2105.290 2.400 2109.690 2.680 ;
        RECT 2110.810 2.400 2115.670 2.680 ;
        RECT 2116.790 2.400 2121.650 2.680 ;
        RECT 2122.770 2.400 2127.630 2.680 ;
        RECT 2128.750 2.400 2133.610 2.680 ;
        RECT 2134.730 2.400 2139.130 2.680 ;
        RECT 2140.250 2.400 2145.110 2.680 ;
        RECT 2146.230 2.400 2151.090 2.680 ;
        RECT 2152.210 2.400 2157.070 2.680 ;
        RECT 2158.190 2.400 2163.050 2.680 ;
        RECT 2164.170 2.400 2168.570 2.680 ;
        RECT 2169.690 2.400 2174.550 2.680 ;
        RECT 2175.670 2.400 2180.530 2.680 ;
        RECT 2181.650 2.400 2186.510 2.680 ;
        RECT 2187.630 2.400 2192.490 2.680 ;
        RECT 2193.610 2.400 2198.010 2.680 ;
        RECT 2199.130 2.400 2203.990 2.680 ;
        RECT 2205.110 2.400 2209.970 2.680 ;
        RECT 2211.090 2.400 2215.950 2.680 ;
        RECT 2217.070 2.400 2221.470 2.680 ;
        RECT 2222.590 2.400 2227.450 2.680 ;
        RECT 2228.570 2.400 2233.430 2.680 ;
        RECT 2234.550 2.400 2239.410 2.680 ;
        RECT 2240.530 2.400 2245.390 2.680 ;
        RECT 2246.510 2.400 2250.910 2.680 ;
        RECT 2252.030 2.400 2256.890 2.680 ;
        RECT 2258.010 2.400 2262.870 2.680 ;
        RECT 2263.990 2.400 2268.850 2.680 ;
        RECT 2269.970 2.400 2274.830 2.680 ;
        RECT 2275.950 2.400 2280.350 2.680 ;
        RECT 2281.470 2.400 2286.330 2.680 ;
        RECT 2287.450 2.400 2292.310 2.680 ;
        RECT 2293.430 2.400 2298.290 2.680 ;
        RECT 2299.410 2.400 2304.270 2.680 ;
        RECT 2305.390 2.400 2309.790 2.680 ;
        RECT 2310.910 2.400 2315.770 2.680 ;
        RECT 2316.890 2.400 2321.750 2.680 ;
        RECT 2322.870 2.400 2327.730 2.680 ;
        RECT 2328.850 2.400 2333.710 2.680 ;
        RECT 2334.830 2.400 2339.230 2.680 ;
        RECT 2340.350 2.400 2345.210 2.680 ;
        RECT 2346.330 2.400 2351.190 2.680 ;
        RECT 2352.310 2.400 2357.170 2.680 ;
        RECT 2358.290 2.400 2363.150 2.680 ;
        RECT 2364.270 2.400 2368.670 2.680 ;
        RECT 2369.790 2.400 2374.650 2.680 ;
        RECT 2375.770 2.400 2380.630 2.680 ;
        RECT 2381.750 2.400 2386.610 2.680 ;
        RECT 2387.730 2.400 2392.590 2.680 ;
        RECT 2393.710 2.400 2398.110 2.680 ;
        RECT 2399.230 2.400 2404.090 2.680 ;
        RECT 2405.210 2.400 2410.070 2.680 ;
        RECT 2411.190 2.400 2416.050 2.680 ;
        RECT 2417.170 2.400 2422.030 2.680 ;
        RECT 2423.150 2.400 2427.550 2.680 ;
        RECT 2428.670 2.400 2433.530 2.680 ;
        RECT 2434.650 2.400 2439.510 2.680 ;
        RECT 2440.630 2.400 2445.490 2.680 ;
        RECT 2446.610 2.400 2451.470 2.680 ;
        RECT 2452.590 2.400 2456.990 2.680 ;
        RECT 2458.110 2.400 2462.970 2.680 ;
        RECT 2464.090 2.400 2468.950 2.680 ;
        RECT 2470.070 2.400 2474.930 2.680 ;
        RECT 2476.050 2.400 2480.910 2.680 ;
        RECT 2482.030 2.400 2486.430 2.680 ;
        RECT 2487.550 2.400 2492.410 2.680 ;
        RECT 2493.530 2.400 2498.390 2.680 ;
        RECT 2499.510 2.400 2504.370 2.680 ;
        RECT 2505.490 2.400 2510.350 2.680 ;
        RECT 2511.470 2.400 2515.870 2.680 ;
        RECT 2516.990 2.400 2521.850 2.680 ;
        RECT 2522.970 2.400 2527.830 2.680 ;
        RECT 2528.950 2.400 2533.810 2.680 ;
        RECT 2534.930 2.400 2539.790 2.680 ;
        RECT 2540.910 2.400 2545.310 2.680 ;
        RECT 2546.430 2.400 2551.290 2.680 ;
        RECT 2552.410 2.400 2557.270 2.680 ;
        RECT 2558.390 2.400 2563.250 2.680 ;
        RECT 2564.370 2.400 2569.230 2.680 ;
        RECT 2570.350 2.400 2574.750 2.680 ;
        RECT 2575.870 2.400 2580.730 2.680 ;
        RECT 2581.850 2.400 2586.710 2.680 ;
        RECT 2587.830 2.400 2592.690 2.680 ;
        RECT 2593.810 2.400 2598.670 2.680 ;
        RECT 2599.790 2.400 2604.190 2.680 ;
        RECT 2605.310 2.400 2610.170 2.680 ;
        RECT 2611.290 2.400 2616.150 2.680 ;
        RECT 2617.270 2.400 2622.130 2.680 ;
        RECT 2623.250 2.400 2628.110 2.680 ;
        RECT 2629.230 2.400 2633.630 2.680 ;
        RECT 2634.750 2.400 2639.610 2.680 ;
        RECT 2640.730 2.400 2645.590 2.680 ;
        RECT 2646.710 2.400 2651.570 2.680 ;
        RECT 2652.690 2.400 2657.550 2.680 ;
        RECT 2658.670 2.400 2663.070 2.680 ;
        RECT 2664.190 2.400 2669.050 2.680 ;
        RECT 2670.170 2.400 2675.030 2.680 ;
        RECT 2676.150 2.400 2681.010 2.680 ;
        RECT 2682.130 2.400 2686.990 2.680 ;
        RECT 2688.110 2.400 2692.510 2.680 ;
        RECT 2693.630 2.400 2698.490 2.680 ;
        RECT 2699.610 2.400 2704.470 2.680 ;
        RECT 2705.590 2.400 2710.450 2.680 ;
        RECT 2711.570 2.400 2716.430 2.680 ;
        RECT 2717.550 2.400 2721.950 2.680 ;
        RECT 2723.070 2.400 2727.930 2.680 ;
        RECT 2729.050 2.400 2733.910 2.680 ;
        RECT 2735.030 2.400 2739.890 2.680 ;
        RECT 2741.010 2.400 2745.870 2.680 ;
        RECT 2746.990 2.400 2751.390 2.680 ;
        RECT 2752.510 2.400 2757.370 2.680 ;
        RECT 2758.490 2.400 2763.350 2.680 ;
        RECT 2764.470 2.400 2769.330 2.680 ;
        RECT 2770.450 2.400 2775.310 2.680 ;
        RECT 2776.430 2.400 2780.830 2.680 ;
        RECT 2781.950 2.400 2786.810 2.680 ;
        RECT 2787.930 2.400 2792.790 2.680 ;
        RECT 2793.910 2.400 2798.770 2.680 ;
        RECT 2799.890 2.400 2804.750 2.680 ;
        RECT 2805.870 2.400 2810.270 2.680 ;
        RECT 2811.390 2.400 2816.250 2.680 ;
        RECT 2817.370 2.400 2822.230 2.680 ;
        RECT 2823.350 2.400 2828.210 2.680 ;
        RECT 2829.330 2.400 2834.190 2.680 ;
        RECT 2835.310 2.400 2839.710 2.680 ;
        RECT 2840.830 2.400 2845.690 2.680 ;
        RECT 2846.810 2.400 2851.670 2.680 ;
        RECT 2852.790 2.400 2857.650 2.680 ;
        RECT 2858.770 2.400 2863.630 2.680 ;
        RECT 2864.750 2.400 2869.150 2.680 ;
        RECT 2870.270 2.400 2875.130 2.680 ;
        RECT 2876.250 2.400 2881.110 2.680 ;
        RECT 2882.230 2.400 2887.090 2.680 ;
        RECT 2888.210 2.400 2893.070 2.680 ;
        RECT 2894.190 2.400 2898.590 2.680 ;
        RECT 2899.710 2.400 2904.570 2.680 ;
      LAYER met3 ;
        RECT 2.800 3424.500 2917.600 3425.665 ;
        RECT 1.230 3424.460 2917.600 3424.500 ;
        RECT 1.230 3422.460 2917.200 3424.460 ;
        RECT 1.230 3363.260 2917.600 3422.460 ;
        RECT 2.800 3361.260 2917.600 3363.260 ;
        RECT 1.230 3360.540 2917.600 3361.260 ;
        RECT 1.230 3358.540 2917.200 3360.540 ;
        RECT 1.230 3300.700 2917.600 3358.540 ;
        RECT 2.800 3298.700 2917.600 3300.700 ;
        RECT 1.230 3296.620 2917.600 3298.700 ;
        RECT 1.230 3294.620 2917.200 3296.620 ;
        RECT 1.230 3237.460 2917.600 3294.620 ;
        RECT 2.800 3235.460 2917.600 3237.460 ;
        RECT 1.230 3232.700 2917.600 3235.460 ;
        RECT 1.230 3230.700 2917.200 3232.700 ;
        RECT 1.230 3174.900 2917.600 3230.700 ;
        RECT 2.800 3172.900 2917.600 3174.900 ;
        RECT 1.230 3168.780 2917.600 3172.900 ;
        RECT 1.230 3166.780 2917.200 3168.780 ;
        RECT 1.230 3112.340 2917.600 3166.780 ;
        RECT 2.800 3110.340 2917.600 3112.340 ;
        RECT 1.230 3104.860 2917.600 3110.340 ;
        RECT 1.230 3102.860 2917.200 3104.860 ;
        RECT 1.230 3049.100 2917.600 3102.860 ;
        RECT 2.800 3047.100 2917.600 3049.100 ;
        RECT 1.230 3040.940 2917.600 3047.100 ;
        RECT 1.230 3038.940 2917.200 3040.940 ;
        RECT 1.230 2986.540 2917.600 3038.940 ;
        RECT 2.800 2984.540 2917.600 2986.540 ;
        RECT 1.230 2977.020 2917.600 2984.540 ;
        RECT 1.230 2975.020 2917.200 2977.020 ;
        RECT 1.230 2923.300 2917.600 2975.020 ;
        RECT 2.800 2921.300 2917.600 2923.300 ;
        RECT 1.230 2912.420 2917.600 2921.300 ;
        RECT 1.230 2910.420 2917.200 2912.420 ;
        RECT 1.230 2860.740 2917.600 2910.420 ;
        RECT 2.800 2858.740 2917.600 2860.740 ;
        RECT 1.230 2848.500 2917.600 2858.740 ;
        RECT 1.230 2846.500 2917.200 2848.500 ;
        RECT 1.230 2797.500 2917.600 2846.500 ;
        RECT 2.800 2795.500 2917.600 2797.500 ;
        RECT 1.230 2784.580 2917.600 2795.500 ;
        RECT 1.230 2782.580 2917.200 2784.580 ;
        RECT 1.230 2734.940 2917.600 2782.580 ;
        RECT 2.800 2732.940 2917.600 2734.940 ;
        RECT 1.230 2720.660 2917.600 2732.940 ;
        RECT 1.230 2718.660 2917.200 2720.660 ;
        RECT 1.230 2672.380 2917.600 2718.660 ;
        RECT 2.800 2670.380 2917.600 2672.380 ;
        RECT 1.230 2656.740 2917.600 2670.380 ;
        RECT 1.230 2654.740 2917.200 2656.740 ;
        RECT 1.230 2609.140 2917.600 2654.740 ;
        RECT 2.800 2607.140 2917.600 2609.140 ;
        RECT 1.230 2592.820 2917.600 2607.140 ;
        RECT 1.230 2590.820 2917.200 2592.820 ;
        RECT 1.230 2546.580 2917.600 2590.820 ;
        RECT 2.800 2544.580 2917.600 2546.580 ;
        RECT 1.230 2528.900 2917.600 2544.580 ;
        RECT 1.230 2526.900 2917.200 2528.900 ;
        RECT 1.230 2483.340 2917.600 2526.900 ;
        RECT 2.800 2481.340 2917.600 2483.340 ;
        RECT 1.230 2464.980 2917.600 2481.340 ;
        RECT 1.230 2462.980 2917.200 2464.980 ;
        RECT 1.230 2420.780 2917.600 2462.980 ;
        RECT 2.800 2418.780 2917.600 2420.780 ;
        RECT 1.230 2401.060 2917.600 2418.780 ;
        RECT 1.230 2399.060 2917.200 2401.060 ;
        RECT 1.230 2357.540 2917.600 2399.060 ;
        RECT 2.800 2355.540 2917.600 2357.540 ;
        RECT 1.230 2336.460 2917.600 2355.540 ;
        RECT 1.230 2334.460 2917.200 2336.460 ;
        RECT 1.230 2294.980 2917.600 2334.460 ;
        RECT 2.800 2292.980 2917.600 2294.980 ;
        RECT 1.230 2272.540 2917.600 2292.980 ;
        RECT 1.230 2270.540 2917.200 2272.540 ;
        RECT 1.230 2232.420 2917.600 2270.540 ;
        RECT 2.800 2230.420 2917.600 2232.420 ;
        RECT 1.230 2208.620 2917.600 2230.420 ;
        RECT 1.230 2206.620 2917.200 2208.620 ;
        RECT 1.230 2169.180 2917.600 2206.620 ;
        RECT 2.800 2167.180 2917.600 2169.180 ;
        RECT 1.230 2144.700 2917.600 2167.180 ;
        RECT 1.230 2142.700 2917.200 2144.700 ;
        RECT 1.230 2106.620 2917.600 2142.700 ;
        RECT 2.800 2104.620 2917.600 2106.620 ;
        RECT 1.230 2080.780 2917.600 2104.620 ;
        RECT 1.230 2078.780 2917.200 2080.780 ;
        RECT 1.230 2043.380 2917.600 2078.780 ;
        RECT 2.800 2041.380 2917.600 2043.380 ;
        RECT 1.230 2016.860 2917.600 2041.380 ;
        RECT 1.230 2014.860 2917.200 2016.860 ;
        RECT 1.230 1980.820 2917.600 2014.860 ;
        RECT 2.800 1978.820 2917.600 1980.820 ;
        RECT 1.230 1952.940 2917.600 1978.820 ;
        RECT 1.230 1950.940 2917.200 1952.940 ;
        RECT 1.230 1917.580 2917.600 1950.940 ;
        RECT 2.800 1915.580 2917.600 1917.580 ;
        RECT 1.230 1889.020 2917.600 1915.580 ;
        RECT 1.230 1887.020 2917.200 1889.020 ;
        RECT 1.230 1855.020 2917.600 1887.020 ;
        RECT 2.800 1853.020 2917.600 1855.020 ;
        RECT 1.230 1825.100 2917.600 1853.020 ;
        RECT 1.230 1823.100 2917.200 1825.100 ;
        RECT 1.230 1792.460 2917.600 1823.100 ;
        RECT 2.800 1790.460 2917.600 1792.460 ;
        RECT 1.230 1760.500 2917.600 1790.460 ;
        RECT 1.230 1758.500 2917.200 1760.500 ;
        RECT 1.230 1729.220 2917.600 1758.500 ;
        RECT 2.800 1727.220 2917.600 1729.220 ;
        RECT 1.230 1696.580 2917.600 1727.220 ;
        RECT 1.230 1694.580 2917.200 1696.580 ;
        RECT 1.230 1666.660 2917.600 1694.580 ;
        RECT 2.800 1664.660 2917.600 1666.660 ;
        RECT 1.230 1632.660 2917.600 1664.660 ;
        RECT 1.230 1630.660 2917.200 1632.660 ;
        RECT 1.230 1603.420 2917.600 1630.660 ;
        RECT 2.800 1601.420 2917.600 1603.420 ;
        RECT 1.230 1568.740 2917.600 1601.420 ;
        RECT 1.230 1566.740 2917.200 1568.740 ;
        RECT 1.230 1540.860 2917.600 1566.740 ;
        RECT 2.800 1538.860 2917.600 1540.860 ;
        RECT 1.230 1504.820 2917.600 1538.860 ;
        RECT 1.230 1502.820 2917.200 1504.820 ;
        RECT 1.230 1477.620 2917.600 1502.820 ;
        RECT 2.800 1475.620 2917.600 1477.620 ;
        RECT 1.230 1440.900 2917.600 1475.620 ;
        RECT 1.230 1438.900 2917.200 1440.900 ;
        RECT 1.230 1415.060 2917.600 1438.900 ;
        RECT 2.800 1413.060 2917.600 1415.060 ;
        RECT 1.230 1376.980 2917.600 1413.060 ;
        RECT 1.230 1374.980 2917.200 1376.980 ;
        RECT 1.230 1352.500 2917.600 1374.980 ;
        RECT 2.800 1350.500 2917.600 1352.500 ;
        RECT 1.230 1313.060 2917.600 1350.500 ;
        RECT 1.230 1311.060 2917.200 1313.060 ;
        RECT 1.230 1289.260 2917.600 1311.060 ;
        RECT 2.800 1287.260 2917.600 1289.260 ;
        RECT 1.230 1249.140 2917.600 1287.260 ;
        RECT 1.230 1247.140 2917.200 1249.140 ;
        RECT 1.230 1226.700 2917.600 1247.140 ;
        RECT 2.800 1224.700 2917.600 1226.700 ;
        RECT 1.230 1184.540 2917.600 1224.700 ;
        RECT 1.230 1182.540 2917.200 1184.540 ;
        RECT 1.230 1163.460 2917.600 1182.540 ;
        RECT 2.800 1161.460 2917.600 1163.460 ;
        RECT 1.230 1120.620 2917.600 1161.460 ;
        RECT 1.230 1118.620 2917.200 1120.620 ;
        RECT 1.230 1100.900 2917.600 1118.620 ;
        RECT 2.800 1098.900 2917.600 1100.900 ;
        RECT 1.230 1056.700 2917.600 1098.900 ;
        RECT 1.230 1054.700 2917.200 1056.700 ;
        RECT 1.230 1037.660 2917.600 1054.700 ;
        RECT 2.800 1035.660 2917.600 1037.660 ;
        RECT 1.230 992.780 2917.600 1035.660 ;
        RECT 1.230 990.780 2917.200 992.780 ;
        RECT 1.230 975.100 2917.600 990.780 ;
        RECT 2.800 973.100 2917.600 975.100 ;
        RECT 1.230 928.860 2917.600 973.100 ;
        RECT 1.230 926.860 2917.200 928.860 ;
        RECT 1.230 912.540 2917.600 926.860 ;
        RECT 2.800 910.540 2917.600 912.540 ;
        RECT 1.230 864.940 2917.600 910.540 ;
        RECT 1.230 862.940 2917.200 864.940 ;
        RECT 1.230 849.300 2917.600 862.940 ;
        RECT 2.800 847.300 2917.600 849.300 ;
        RECT 1.230 801.020 2917.600 847.300 ;
        RECT 1.230 799.020 2917.200 801.020 ;
        RECT 1.230 786.740 2917.600 799.020 ;
        RECT 2.800 784.740 2917.600 786.740 ;
        RECT 1.230 737.100 2917.600 784.740 ;
        RECT 1.230 735.100 2917.200 737.100 ;
        RECT 1.230 723.500 2917.600 735.100 ;
        RECT 2.800 721.500 2917.600 723.500 ;
        RECT 1.230 673.180 2917.600 721.500 ;
        RECT 1.230 671.180 2917.200 673.180 ;
        RECT 1.230 660.940 2917.600 671.180 ;
        RECT 2.800 658.940 2917.600 660.940 ;
        RECT 1.230 608.580 2917.600 658.940 ;
        RECT 1.230 606.580 2917.200 608.580 ;
        RECT 1.230 597.700 2917.600 606.580 ;
        RECT 2.800 595.700 2917.600 597.700 ;
        RECT 1.230 544.660 2917.600 595.700 ;
        RECT 1.230 542.660 2917.200 544.660 ;
        RECT 1.230 535.140 2917.600 542.660 ;
        RECT 2.800 533.140 2917.600 535.140 ;
        RECT 1.230 480.740 2917.600 533.140 ;
        RECT 1.230 478.740 2917.200 480.740 ;
        RECT 1.230 472.580 2917.600 478.740 ;
        RECT 2.800 470.580 2917.600 472.580 ;
        RECT 1.230 416.820 2917.600 470.580 ;
        RECT 1.230 414.820 2917.200 416.820 ;
        RECT 1.230 409.340 2917.600 414.820 ;
        RECT 2.800 407.340 2917.600 409.340 ;
        RECT 1.230 352.900 2917.600 407.340 ;
        RECT 1.230 350.900 2917.200 352.900 ;
        RECT 1.230 346.780 2917.600 350.900 ;
        RECT 2.800 344.780 2917.600 346.780 ;
        RECT 1.230 288.980 2917.600 344.780 ;
        RECT 1.230 286.980 2917.200 288.980 ;
        RECT 1.230 283.540 2917.600 286.980 ;
        RECT 2.800 281.540 2917.600 283.540 ;
        RECT 1.230 225.060 2917.600 281.540 ;
        RECT 1.230 223.060 2917.200 225.060 ;
        RECT 1.230 220.980 2917.600 223.060 ;
        RECT 2.800 218.980 2917.600 220.980 ;
        RECT 1.230 161.140 2917.600 218.980 ;
        RECT 1.230 159.140 2917.200 161.140 ;
        RECT 1.230 157.740 2917.600 159.140 ;
        RECT 2.800 156.575 2917.600 157.740 ;
      LAYER met4 ;
        RECT 223.855 199.415 225.770 3231.185 ;
        RECT 229.670 199.415 244.370 3231.185 ;
        RECT 248.270 199.415 278.570 3231.185 ;
        RECT 282.470 3200.095 297.170 3231.185 ;
        RECT 301.070 3200.095 315.770 3231.185 ;
        RECT 319.670 3200.095 334.370 3231.185 ;
        RECT 338.270 3200.095 368.570 3231.185 ;
        RECT 372.470 3200.095 387.170 3231.185 ;
        RECT 391.070 3200.095 405.770 3231.185 ;
        RECT 409.670 3200.095 424.370 3231.185 ;
        RECT 428.270 3200.095 458.570 3231.185 ;
        RECT 462.470 3200.095 477.170 3231.185 ;
        RECT 481.070 3200.095 495.770 3231.185 ;
        RECT 499.670 3200.095 514.370 3231.185 ;
        RECT 518.270 3200.095 548.570 3231.185 ;
        RECT 552.470 3200.095 567.170 3231.185 ;
        RECT 571.070 3200.095 585.770 3231.185 ;
        RECT 589.670 3200.095 604.370 3231.185 ;
        RECT 608.270 3200.095 638.570 3231.185 ;
        RECT 282.470 2865.400 638.570 3200.095 ;
        RECT 282.470 2784.600 297.170 2865.400 ;
        RECT 301.070 2784.600 315.770 2865.400 ;
        RECT 319.670 2784.600 334.370 2865.400 ;
        RECT 338.270 2784.600 368.570 2865.400 ;
        RECT 372.470 2784.600 387.170 2865.400 ;
        RECT 391.070 2784.600 405.770 2865.400 ;
        RECT 409.670 2784.600 424.370 2865.400 ;
        RECT 428.270 2784.600 458.570 2865.400 ;
        RECT 462.470 2784.600 477.170 2865.400 ;
        RECT 481.070 2784.600 495.770 2865.400 ;
        RECT 499.670 2784.600 514.370 2865.400 ;
        RECT 518.270 2784.600 548.570 2865.400 ;
        RECT 552.470 2784.600 567.170 2865.400 ;
        RECT 571.070 2784.600 585.770 2865.400 ;
        RECT 589.670 2784.600 604.370 2865.400 ;
        RECT 608.270 2784.600 638.570 2865.400 ;
        RECT 642.470 2784.600 657.170 3231.185 ;
        RECT 661.070 2784.600 675.770 3231.185 ;
        RECT 679.670 3200.095 694.370 3231.185 ;
        RECT 698.270 3200.095 728.570 3231.185 ;
        RECT 732.470 3200.095 747.170 3231.185 ;
        RECT 751.070 3200.095 765.770 3231.185 ;
        RECT 769.670 3200.095 784.370 3231.185 ;
        RECT 788.270 3200.095 818.570 3231.185 ;
        RECT 822.470 3200.095 837.170 3231.185 ;
        RECT 841.070 3200.095 855.770 3231.185 ;
        RECT 859.670 3200.095 874.370 3231.185 ;
        RECT 878.270 3200.095 908.570 3231.185 ;
        RECT 912.470 3200.095 927.170 3231.185 ;
        RECT 931.070 3200.095 945.770 3231.185 ;
        RECT 949.670 3200.095 964.370 3231.185 ;
        RECT 968.270 3200.095 998.570 3231.185 ;
        RECT 1002.470 3200.095 1017.170 3231.185 ;
        RECT 679.670 2865.400 1017.170 3200.095 ;
        RECT 679.670 2784.600 694.370 2865.400 ;
        RECT 698.270 2784.600 728.570 2865.400 ;
        RECT 732.470 2784.600 747.170 2865.400 ;
        RECT 751.070 2784.600 765.770 2865.400 ;
        RECT 769.670 2784.600 784.370 2865.400 ;
        RECT 788.270 2784.600 818.570 2865.400 ;
        RECT 822.470 2784.600 837.170 2865.400 ;
        RECT 841.070 2784.600 855.770 2865.400 ;
        RECT 859.670 2784.600 874.370 2865.400 ;
        RECT 878.270 2784.600 908.570 2865.400 ;
        RECT 912.470 2784.600 927.170 2865.400 ;
        RECT 931.070 2784.600 945.770 2865.400 ;
        RECT 949.670 2784.600 964.370 2865.400 ;
        RECT 968.270 2784.600 998.570 2865.400 ;
        RECT 1002.470 2784.600 1017.170 2865.400 ;
        RECT 1021.070 2784.600 1035.770 3231.185 ;
        RECT 1039.670 2784.600 1054.370 3231.185 ;
        RECT 1058.270 3200.095 1088.570 3231.185 ;
        RECT 1092.470 3200.095 1107.170 3231.185 ;
        RECT 1111.070 3200.095 1125.770 3231.185 ;
        RECT 1129.670 3200.095 1144.370 3231.185 ;
        RECT 1148.270 3200.095 1178.570 3231.185 ;
        RECT 1182.470 3200.095 1197.170 3231.185 ;
        RECT 1201.070 3200.095 1215.770 3231.185 ;
        RECT 1219.670 3200.095 1234.370 3231.185 ;
        RECT 1238.270 3200.095 1268.570 3231.185 ;
        RECT 1272.470 3200.095 1287.170 3231.185 ;
        RECT 1291.070 3200.095 1305.770 3231.185 ;
        RECT 1309.670 3200.095 1324.370 3231.185 ;
        RECT 1328.270 3200.095 1358.570 3231.185 ;
        RECT 1362.470 3200.095 1377.170 3231.185 ;
        RECT 1381.070 3200.095 1395.770 3231.185 ;
        RECT 1399.670 3200.095 1414.370 3231.185 ;
        RECT 1418.270 3200.095 1448.570 3231.185 ;
        RECT 1058.270 2865.400 1448.570 3200.095 ;
        RECT 1058.270 2784.600 1088.570 2865.400 ;
        RECT 1092.470 2784.600 1107.170 2865.400 ;
        RECT 1111.070 2784.600 1125.770 2865.400 ;
        RECT 1129.670 2784.600 1144.370 2865.400 ;
        RECT 1148.270 2784.600 1178.570 2865.400 ;
        RECT 1182.470 2784.600 1197.170 2865.400 ;
        RECT 1201.070 2784.600 1215.770 2865.400 ;
        RECT 1219.670 2784.600 1234.370 2865.400 ;
        RECT 1238.270 2784.600 1268.570 2865.400 ;
        RECT 1272.470 2784.600 1287.170 2865.400 ;
        RECT 1291.070 2784.600 1305.770 2865.400 ;
        RECT 1309.670 2784.600 1324.370 2865.400 ;
        RECT 1328.270 2784.600 1358.570 2865.400 ;
        RECT 1362.470 2784.600 1377.170 2865.400 ;
        RECT 1381.070 2784.600 1395.770 2865.400 ;
        RECT 1399.670 2784.600 1414.370 2865.400 ;
        RECT 1418.270 2784.600 1448.570 2865.400 ;
        RECT 1452.470 2784.600 1467.170 3231.185 ;
        RECT 1471.070 2784.600 1485.770 3231.185 ;
        RECT 1489.670 2784.600 1504.370 3231.185 ;
        RECT 1508.270 2784.600 1538.570 3231.185 ;
        RECT 282.470 2465.400 1538.570 2784.600 ;
        RECT 282.470 2301.140 297.170 2465.400 ;
        RECT 301.070 2301.140 315.770 2465.400 ;
        RECT 319.670 2301.140 334.370 2465.400 ;
        RECT 338.270 2301.140 368.570 2465.400 ;
        RECT 372.470 2301.140 387.170 2465.400 ;
        RECT 391.070 2301.140 405.770 2465.400 ;
        RECT 409.670 2301.140 424.370 2465.400 ;
        RECT 428.270 2301.140 458.570 2465.400 ;
        RECT 462.470 2301.140 477.170 2465.400 ;
        RECT 481.070 2301.140 495.770 2465.400 ;
        RECT 499.670 2301.140 514.370 2465.400 ;
        RECT 518.270 2301.140 548.570 2465.400 ;
        RECT 552.470 2301.140 567.170 2465.400 ;
        RECT 571.070 2301.140 585.770 2465.400 ;
        RECT 589.670 2301.140 604.370 2465.400 ;
        RECT 608.270 2301.140 638.570 2465.400 ;
        RECT 642.470 2301.140 657.170 2465.400 ;
        RECT 661.070 2301.140 675.770 2465.400 ;
        RECT 679.670 2301.140 694.370 2465.400 ;
        RECT 698.270 2301.140 728.570 2465.400 ;
        RECT 732.470 2301.140 747.170 2465.400 ;
        RECT 751.070 2301.140 765.770 2465.400 ;
        RECT 769.670 2301.140 784.370 2465.400 ;
        RECT 788.270 2301.140 818.570 2465.400 ;
        RECT 822.470 2301.140 837.170 2465.400 ;
        RECT 841.070 2301.140 855.770 2465.400 ;
        RECT 859.670 2301.140 874.370 2465.400 ;
        RECT 878.270 2301.140 908.570 2465.400 ;
        RECT 912.470 2301.140 927.170 2465.400 ;
        RECT 931.070 2301.140 945.770 2465.400 ;
        RECT 949.670 2301.140 964.370 2465.400 ;
        RECT 968.270 2301.140 998.570 2465.400 ;
        RECT 282.470 1865.400 998.570 2301.140 ;
        RECT 282.470 1751.140 297.170 1865.400 ;
        RECT 301.070 1751.140 315.770 1865.400 ;
        RECT 319.670 1751.140 334.370 1865.400 ;
        RECT 338.270 1751.140 368.570 1865.400 ;
        RECT 372.470 1751.140 387.170 1865.400 ;
        RECT 391.070 1751.140 405.770 1865.400 ;
        RECT 409.670 1751.140 424.370 1865.400 ;
        RECT 428.270 1751.140 458.570 1865.400 ;
        RECT 462.470 1751.140 477.170 1865.400 ;
        RECT 481.070 1751.140 495.770 1865.400 ;
        RECT 499.670 1751.140 514.370 1865.400 ;
        RECT 518.270 1751.140 548.570 1865.400 ;
        RECT 552.470 1751.140 567.170 1865.400 ;
        RECT 571.070 1751.140 585.770 1865.400 ;
        RECT 589.670 1751.140 604.370 1865.400 ;
        RECT 608.270 1751.140 638.570 1865.400 ;
        RECT 642.470 1751.140 657.170 1865.400 ;
        RECT 661.070 1751.140 675.770 1865.400 ;
        RECT 679.670 1751.140 694.370 1865.400 ;
        RECT 698.270 1751.140 728.570 1865.400 ;
        RECT 732.470 1751.140 747.170 1865.400 ;
        RECT 751.070 1751.140 765.770 1865.400 ;
        RECT 769.670 1751.140 784.370 1865.400 ;
        RECT 788.270 1751.140 818.570 1865.400 ;
        RECT 822.470 1751.140 837.170 1865.400 ;
        RECT 841.070 1751.140 855.770 1865.400 ;
        RECT 859.670 1751.140 874.370 1865.400 ;
        RECT 878.270 1751.140 908.570 1865.400 ;
        RECT 912.470 1751.140 927.170 1865.400 ;
        RECT 931.070 1751.140 945.770 1865.400 ;
        RECT 949.670 1751.140 964.370 1865.400 ;
        RECT 968.270 1751.140 998.570 1865.400 ;
        RECT 282.470 1315.400 998.570 1751.140 ;
        RECT 282.470 1201.140 297.170 1315.400 ;
        RECT 301.070 1201.140 315.770 1315.400 ;
        RECT 319.670 1201.140 334.370 1315.400 ;
        RECT 338.270 1201.140 368.570 1315.400 ;
        RECT 372.470 1201.140 387.170 1315.400 ;
        RECT 391.070 1201.140 405.770 1315.400 ;
        RECT 409.670 1201.140 424.370 1315.400 ;
        RECT 428.270 1201.140 458.570 1315.400 ;
        RECT 462.470 1201.140 477.170 1315.400 ;
        RECT 481.070 1201.140 495.770 1315.400 ;
        RECT 499.670 1201.140 514.370 1315.400 ;
        RECT 518.270 1201.140 548.570 1315.400 ;
        RECT 552.470 1201.140 567.170 1315.400 ;
        RECT 571.070 1201.140 585.770 1315.400 ;
        RECT 589.670 1201.140 604.370 1315.400 ;
        RECT 608.270 1201.140 638.570 1315.400 ;
        RECT 642.470 1201.140 657.170 1315.400 ;
        RECT 661.070 1201.140 675.770 1315.400 ;
        RECT 679.670 1201.140 694.370 1315.400 ;
        RECT 698.270 1201.140 728.570 1315.400 ;
        RECT 732.470 1201.140 747.170 1315.400 ;
        RECT 751.070 1201.140 765.770 1315.400 ;
        RECT 769.670 1201.140 784.370 1315.400 ;
        RECT 788.270 1201.140 818.570 1315.400 ;
        RECT 822.470 1201.140 837.170 1315.400 ;
        RECT 841.070 1201.140 855.770 1315.400 ;
        RECT 859.670 1201.140 874.370 1315.400 ;
        RECT 878.270 1201.140 908.570 1315.400 ;
        RECT 912.470 1201.140 927.170 1315.400 ;
        RECT 931.070 1201.140 945.770 1315.400 ;
        RECT 949.670 1201.140 964.370 1315.400 ;
        RECT 968.270 1201.140 998.570 1315.400 ;
        RECT 282.470 765.400 998.570 1201.140 ;
        RECT 282.470 651.140 297.170 765.400 ;
        RECT 301.070 651.140 315.770 765.400 ;
        RECT 319.670 651.140 334.370 765.400 ;
        RECT 338.270 651.140 368.570 765.400 ;
        RECT 372.470 651.140 387.170 765.400 ;
        RECT 391.070 651.140 405.770 765.400 ;
        RECT 409.670 651.140 424.370 765.400 ;
        RECT 428.270 651.140 458.570 765.400 ;
        RECT 462.470 651.140 477.170 765.400 ;
        RECT 481.070 651.140 495.770 765.400 ;
        RECT 499.670 651.140 514.370 765.400 ;
        RECT 518.270 651.140 548.570 765.400 ;
        RECT 552.470 651.140 567.170 765.400 ;
        RECT 571.070 651.140 585.770 765.400 ;
        RECT 589.670 651.140 604.370 765.400 ;
        RECT 608.270 651.140 638.570 765.400 ;
        RECT 642.470 651.140 657.170 765.400 ;
        RECT 661.070 651.140 675.770 765.400 ;
        RECT 679.670 651.140 694.370 765.400 ;
        RECT 698.270 651.140 728.570 765.400 ;
        RECT 732.470 651.140 747.170 765.400 ;
        RECT 751.070 651.140 765.770 765.400 ;
        RECT 769.670 651.140 784.370 765.400 ;
        RECT 788.270 651.140 818.570 765.400 ;
        RECT 822.470 651.140 837.170 765.400 ;
        RECT 841.070 651.140 855.770 765.400 ;
        RECT 859.670 651.140 874.370 765.400 ;
        RECT 878.270 651.140 908.570 765.400 ;
        RECT 912.470 651.140 927.170 765.400 ;
        RECT 931.070 651.140 945.770 765.400 ;
        RECT 949.670 651.140 964.370 765.400 ;
        RECT 968.270 651.140 998.570 765.400 ;
        RECT 282.470 215.400 998.570 651.140 ;
        RECT 282.470 199.415 297.170 215.400 ;
        RECT 301.070 199.415 315.770 215.400 ;
        RECT 319.670 199.415 334.370 215.400 ;
        RECT 338.270 199.415 368.570 215.400 ;
        RECT 372.470 199.415 387.170 215.400 ;
        RECT 391.070 199.415 405.770 215.400 ;
        RECT 409.670 199.415 424.370 215.400 ;
        RECT 428.270 199.415 458.570 215.400 ;
        RECT 462.470 199.415 477.170 215.400 ;
        RECT 481.070 199.415 495.770 215.400 ;
        RECT 499.670 199.415 514.370 215.400 ;
        RECT 518.270 199.415 548.570 215.400 ;
        RECT 552.470 199.415 567.170 215.400 ;
        RECT 571.070 199.415 585.770 215.400 ;
        RECT 589.670 199.415 604.370 215.400 ;
        RECT 608.270 199.415 638.570 215.400 ;
        RECT 642.470 199.415 657.170 215.400 ;
        RECT 661.070 199.415 675.770 215.400 ;
        RECT 679.670 199.415 694.370 215.400 ;
        RECT 698.270 199.415 728.570 215.400 ;
        RECT 732.470 199.415 747.170 215.400 ;
        RECT 751.070 199.415 765.770 215.400 ;
        RECT 769.670 199.415 784.370 215.400 ;
        RECT 788.270 199.415 818.570 215.400 ;
        RECT 822.470 199.415 837.170 215.400 ;
        RECT 841.070 199.415 855.770 215.400 ;
        RECT 859.670 199.415 874.370 215.400 ;
        RECT 878.270 199.415 908.570 215.400 ;
        RECT 912.470 199.415 927.170 215.400 ;
        RECT 931.070 199.415 945.770 215.400 ;
        RECT 949.670 199.415 964.370 215.400 ;
        RECT 968.270 199.415 998.570 215.400 ;
        RECT 1002.470 199.415 1017.170 2465.400 ;
        RECT 1021.070 199.415 1035.770 2465.400 ;
        RECT 1039.670 199.415 1054.370 2465.400 ;
        RECT 1058.270 2301.140 1088.570 2465.400 ;
        RECT 1092.470 2301.140 1107.170 2465.400 ;
        RECT 1111.070 2301.140 1125.770 2465.400 ;
        RECT 1129.670 2301.140 1144.370 2465.400 ;
        RECT 1148.270 2301.140 1178.570 2465.400 ;
        RECT 1182.470 2301.140 1197.170 2465.400 ;
        RECT 1201.070 2301.140 1215.770 2465.400 ;
        RECT 1219.670 2301.140 1234.370 2465.400 ;
        RECT 1238.270 2301.140 1268.570 2465.400 ;
        RECT 1272.470 2301.140 1287.170 2465.400 ;
        RECT 1291.070 2301.140 1305.770 2465.400 ;
        RECT 1309.670 2301.140 1324.370 2465.400 ;
        RECT 1328.270 2301.140 1358.570 2465.400 ;
        RECT 1362.470 2301.140 1377.170 2465.400 ;
        RECT 1381.070 2301.140 1395.770 2465.400 ;
        RECT 1399.670 2301.140 1414.370 2465.400 ;
        RECT 1418.270 2301.140 1448.570 2465.400 ;
        RECT 1452.470 2301.140 1467.170 2465.400 ;
        RECT 1471.070 2301.140 1485.770 2465.400 ;
        RECT 1489.670 2301.140 1504.370 2465.400 ;
        RECT 1508.270 2301.140 1538.570 2465.400 ;
        RECT 1542.470 2301.140 1557.170 3231.185 ;
        RECT 1561.070 2301.140 1575.770 3231.185 ;
        RECT 1579.670 2665.400 2168.570 3231.185 ;
        RECT 1579.670 2301.140 1594.370 2665.400 ;
        RECT 1598.270 2301.140 1628.570 2665.400 ;
        RECT 1632.470 2301.140 1647.170 2665.400 ;
        RECT 1651.070 2301.140 1665.770 2665.400 ;
        RECT 1669.670 2301.140 1684.370 2665.400 ;
        RECT 1688.270 2301.140 1718.570 2665.400 ;
        RECT 1722.470 2301.140 1737.170 2665.400 ;
        RECT 1741.070 2301.140 1755.770 2665.400 ;
        RECT 1759.670 2301.140 1774.370 2665.400 ;
        RECT 1778.270 2301.140 1808.570 2665.400 ;
        RECT 1058.270 1865.400 1808.570 2301.140 ;
        RECT 1058.270 1751.140 1088.570 1865.400 ;
        RECT 1092.470 1751.140 1107.170 1865.400 ;
        RECT 1111.070 1751.140 1125.770 1865.400 ;
        RECT 1129.670 1751.140 1144.370 1865.400 ;
        RECT 1148.270 1751.140 1178.570 1865.400 ;
        RECT 1182.470 1751.140 1197.170 1865.400 ;
        RECT 1201.070 1751.140 1215.770 1865.400 ;
        RECT 1219.670 1751.140 1234.370 1865.400 ;
        RECT 1238.270 1751.140 1268.570 1865.400 ;
        RECT 1272.470 1751.140 1287.170 1865.400 ;
        RECT 1291.070 1751.140 1305.770 1865.400 ;
        RECT 1309.670 1751.140 1324.370 1865.400 ;
        RECT 1328.270 1751.140 1358.570 1865.400 ;
        RECT 1362.470 1751.140 1377.170 1865.400 ;
        RECT 1381.070 1751.140 1395.770 1865.400 ;
        RECT 1399.670 1751.140 1414.370 1865.400 ;
        RECT 1418.270 1751.140 1448.570 1865.400 ;
        RECT 1452.470 1751.140 1467.170 1865.400 ;
        RECT 1471.070 1751.140 1485.770 1865.400 ;
        RECT 1489.670 1751.140 1504.370 1865.400 ;
        RECT 1508.270 1751.140 1538.570 1865.400 ;
        RECT 1542.470 1751.140 1557.170 1865.400 ;
        RECT 1561.070 1751.140 1575.770 1865.400 ;
        RECT 1579.670 1751.140 1594.370 1865.400 ;
        RECT 1598.270 1751.140 1628.570 1865.400 ;
        RECT 1632.470 1751.140 1647.170 1865.400 ;
        RECT 1651.070 1751.140 1665.770 1865.400 ;
        RECT 1669.670 1751.140 1684.370 1865.400 ;
        RECT 1688.270 1751.140 1718.570 1865.400 ;
        RECT 1722.470 1751.140 1737.170 1865.400 ;
        RECT 1741.070 1751.140 1755.770 1865.400 ;
        RECT 1759.670 1751.140 1774.370 1865.400 ;
        RECT 1778.270 1751.140 1808.570 1865.400 ;
        RECT 1058.270 1315.400 1808.570 1751.140 ;
        RECT 1058.270 1201.140 1088.570 1315.400 ;
        RECT 1092.470 1201.140 1107.170 1315.400 ;
        RECT 1111.070 1201.140 1125.770 1315.400 ;
        RECT 1129.670 1201.140 1144.370 1315.400 ;
        RECT 1148.270 1201.140 1178.570 1315.400 ;
        RECT 1182.470 1201.140 1197.170 1315.400 ;
        RECT 1201.070 1201.140 1215.770 1315.400 ;
        RECT 1219.670 1201.140 1234.370 1315.400 ;
        RECT 1238.270 1201.140 1268.570 1315.400 ;
        RECT 1272.470 1201.140 1287.170 1315.400 ;
        RECT 1291.070 1201.140 1305.770 1315.400 ;
        RECT 1309.670 1201.140 1324.370 1315.400 ;
        RECT 1328.270 1201.140 1358.570 1315.400 ;
        RECT 1362.470 1201.140 1377.170 1315.400 ;
        RECT 1381.070 1201.140 1395.770 1315.400 ;
        RECT 1399.670 1201.140 1414.370 1315.400 ;
        RECT 1418.270 1201.140 1448.570 1315.400 ;
        RECT 1452.470 1201.140 1467.170 1315.400 ;
        RECT 1471.070 1201.140 1485.770 1315.400 ;
        RECT 1489.670 1201.140 1504.370 1315.400 ;
        RECT 1508.270 1201.140 1538.570 1315.400 ;
        RECT 1542.470 1201.140 1557.170 1315.400 ;
        RECT 1561.070 1201.140 1575.770 1315.400 ;
        RECT 1579.670 1201.140 1594.370 1315.400 ;
        RECT 1598.270 1201.140 1628.570 1315.400 ;
        RECT 1632.470 1201.140 1647.170 1315.400 ;
        RECT 1651.070 1201.140 1665.770 1315.400 ;
        RECT 1669.670 1201.140 1684.370 1315.400 ;
        RECT 1688.270 1201.140 1718.570 1315.400 ;
        RECT 1722.470 1201.140 1737.170 1315.400 ;
        RECT 1741.070 1201.140 1755.770 1315.400 ;
        RECT 1759.670 1201.140 1774.370 1315.400 ;
        RECT 1778.270 1201.140 1808.570 1315.400 ;
        RECT 1058.270 765.400 1808.570 1201.140 ;
        RECT 1058.270 651.140 1088.570 765.400 ;
        RECT 1092.470 651.140 1107.170 765.400 ;
        RECT 1111.070 651.140 1125.770 765.400 ;
        RECT 1129.670 651.140 1144.370 765.400 ;
        RECT 1148.270 651.140 1178.570 765.400 ;
        RECT 1182.470 651.140 1197.170 765.400 ;
        RECT 1201.070 651.140 1215.770 765.400 ;
        RECT 1219.670 651.140 1234.370 765.400 ;
        RECT 1238.270 651.140 1268.570 765.400 ;
        RECT 1272.470 651.140 1287.170 765.400 ;
        RECT 1291.070 651.140 1305.770 765.400 ;
        RECT 1309.670 651.140 1324.370 765.400 ;
        RECT 1328.270 651.140 1358.570 765.400 ;
        RECT 1362.470 651.140 1377.170 765.400 ;
        RECT 1381.070 651.140 1395.770 765.400 ;
        RECT 1399.670 651.140 1414.370 765.400 ;
        RECT 1418.270 651.140 1448.570 765.400 ;
        RECT 1452.470 651.140 1467.170 765.400 ;
        RECT 1471.070 651.140 1485.770 765.400 ;
        RECT 1489.670 651.140 1504.370 765.400 ;
        RECT 1508.270 651.140 1538.570 765.400 ;
        RECT 1542.470 651.140 1557.170 765.400 ;
        RECT 1561.070 651.140 1575.770 765.400 ;
        RECT 1579.670 651.140 1594.370 765.400 ;
        RECT 1598.270 651.140 1628.570 765.400 ;
        RECT 1632.470 651.140 1647.170 765.400 ;
        RECT 1651.070 651.140 1665.770 765.400 ;
        RECT 1669.670 651.140 1684.370 765.400 ;
        RECT 1688.270 651.140 1718.570 765.400 ;
        RECT 1722.470 651.140 1737.170 765.400 ;
        RECT 1741.070 651.140 1755.770 765.400 ;
        RECT 1759.670 651.140 1774.370 765.400 ;
        RECT 1778.270 651.140 1808.570 765.400 ;
        RECT 1058.270 215.400 1808.570 651.140 ;
        RECT 1058.270 199.415 1088.570 215.400 ;
        RECT 1092.470 199.415 1107.170 215.400 ;
        RECT 1111.070 199.415 1125.770 215.400 ;
        RECT 1129.670 199.415 1144.370 215.400 ;
        RECT 1148.270 199.415 1178.570 215.400 ;
        RECT 1182.470 199.415 1197.170 215.400 ;
        RECT 1201.070 199.415 1215.770 215.400 ;
        RECT 1219.670 199.415 1234.370 215.400 ;
        RECT 1238.270 199.415 1268.570 215.400 ;
        RECT 1272.470 199.415 1287.170 215.400 ;
        RECT 1291.070 199.415 1305.770 215.400 ;
        RECT 1309.670 199.415 1324.370 215.400 ;
        RECT 1328.270 199.415 1358.570 215.400 ;
        RECT 1362.470 199.415 1377.170 215.400 ;
        RECT 1381.070 199.415 1395.770 215.400 ;
        RECT 1399.670 199.415 1414.370 215.400 ;
        RECT 1418.270 199.415 1448.570 215.400 ;
        RECT 1452.470 199.415 1467.170 215.400 ;
        RECT 1471.070 199.415 1485.770 215.400 ;
        RECT 1489.670 199.415 1504.370 215.400 ;
        RECT 1508.270 199.415 1538.570 215.400 ;
        RECT 1542.470 199.415 1557.170 215.400 ;
        RECT 1561.070 199.415 1575.770 215.400 ;
        RECT 1579.670 199.415 1594.370 215.400 ;
        RECT 1598.270 199.415 1628.570 215.400 ;
        RECT 1632.470 199.415 1647.170 215.400 ;
        RECT 1651.070 199.415 1665.770 215.400 ;
        RECT 1669.670 199.415 1684.370 215.400 ;
        RECT 1688.270 199.415 1718.570 215.400 ;
        RECT 1722.470 199.415 1737.170 215.400 ;
        RECT 1741.070 199.415 1755.770 215.400 ;
        RECT 1759.670 199.415 1774.370 215.400 ;
        RECT 1778.270 199.415 1808.570 215.400 ;
        RECT 1812.470 199.415 1827.170 2665.400 ;
        RECT 1831.070 199.415 1845.770 2665.400 ;
        RECT 1849.670 199.415 1864.370 2665.400 ;
        RECT 1868.270 2301.140 1898.570 2665.400 ;
        RECT 1902.470 2301.140 1917.170 2665.400 ;
        RECT 1921.070 2301.140 1935.770 2665.400 ;
        RECT 1939.670 2301.140 1954.370 2665.400 ;
        RECT 1958.270 2301.140 1988.570 2665.400 ;
        RECT 1992.470 2301.140 2007.170 2665.400 ;
        RECT 2011.070 2301.140 2025.770 2665.400 ;
        RECT 2029.670 2301.140 2044.370 2665.400 ;
        RECT 2048.270 2301.140 2078.570 2665.400 ;
        RECT 2082.470 2301.140 2097.170 2665.400 ;
        RECT 2101.070 2301.140 2115.770 2665.400 ;
        RECT 2119.670 2301.140 2134.370 2665.400 ;
        RECT 2138.270 2301.140 2168.570 2665.400 ;
        RECT 2172.470 2301.140 2187.170 3231.185 ;
        RECT 2191.070 2301.140 2205.770 3231.185 ;
        RECT 2209.670 2301.140 2224.370 3231.185 ;
        RECT 2228.270 2301.140 2258.570 3231.185 ;
        RECT 2262.470 2301.140 2277.170 3231.185 ;
        RECT 2281.070 3184.600 2295.770 3231.185 ;
        RECT 2299.670 3184.600 2314.370 3231.185 ;
        RECT 2318.270 3184.600 2348.570 3231.185 ;
        RECT 2352.470 3184.600 2367.170 3231.185 ;
        RECT 2371.070 3184.600 2385.770 3231.185 ;
        RECT 2389.670 3184.600 2404.370 3231.185 ;
        RECT 2408.270 3184.600 2438.570 3231.185 ;
        RECT 2442.470 3184.600 2457.170 3231.185 ;
        RECT 2461.070 3184.600 2475.770 3231.185 ;
        RECT 2479.670 3184.600 2494.370 3231.185 ;
        RECT 2498.270 3184.600 2528.570 3231.185 ;
        RECT 2532.470 3184.600 2547.170 3231.185 ;
        RECT 2551.070 3184.600 2565.770 3231.185 ;
        RECT 2281.070 2915.400 2565.770 3184.600 ;
        RECT 2281.070 2301.140 2295.770 2915.400 ;
        RECT 2299.670 2301.140 2314.370 2915.400 ;
        RECT 2318.270 2301.140 2348.570 2915.400 ;
        RECT 2352.470 2301.140 2367.170 2915.400 ;
        RECT 2371.070 2301.140 2385.770 2915.400 ;
        RECT 2389.670 2301.140 2404.370 2915.400 ;
        RECT 2408.270 2301.140 2438.570 2915.400 ;
        RECT 2442.470 2301.140 2457.170 2915.400 ;
        RECT 2461.070 2301.140 2475.770 2915.400 ;
        RECT 2479.670 2301.140 2494.370 2915.400 ;
        RECT 2498.270 2301.140 2528.570 2915.400 ;
        RECT 2532.470 2301.140 2547.170 2915.400 ;
        RECT 2551.070 2301.140 2565.770 2915.400 ;
        RECT 2569.670 2301.140 2582.480 3231.185 ;
        RECT 1868.270 1865.400 2582.480 2301.140 ;
        RECT 1868.270 1751.140 1898.570 1865.400 ;
        RECT 1902.470 1751.140 1917.170 1865.400 ;
        RECT 1921.070 1751.140 1935.770 1865.400 ;
        RECT 1939.670 1751.140 1954.370 1865.400 ;
        RECT 1958.270 1751.140 1988.570 1865.400 ;
        RECT 1992.470 1751.140 2007.170 1865.400 ;
        RECT 2011.070 1751.140 2025.770 1865.400 ;
        RECT 2029.670 1751.140 2044.370 1865.400 ;
        RECT 2048.270 1751.140 2078.570 1865.400 ;
        RECT 2082.470 1751.140 2097.170 1865.400 ;
        RECT 2101.070 1751.140 2115.770 1865.400 ;
        RECT 2119.670 1751.140 2134.370 1865.400 ;
        RECT 2138.270 1751.140 2168.570 1865.400 ;
        RECT 2172.470 1751.140 2187.170 1865.400 ;
        RECT 2191.070 1751.140 2205.770 1865.400 ;
        RECT 2209.670 1751.140 2224.370 1865.400 ;
        RECT 2228.270 1751.140 2258.570 1865.400 ;
        RECT 2262.470 1751.140 2277.170 1865.400 ;
        RECT 2281.070 1751.140 2295.770 1865.400 ;
        RECT 2299.670 1751.140 2314.370 1865.400 ;
        RECT 2318.270 1751.140 2348.570 1865.400 ;
        RECT 2352.470 1751.140 2367.170 1865.400 ;
        RECT 2371.070 1751.140 2385.770 1865.400 ;
        RECT 2389.670 1751.140 2404.370 1865.400 ;
        RECT 2408.270 1751.140 2438.570 1865.400 ;
        RECT 2442.470 1751.140 2457.170 1865.400 ;
        RECT 2461.070 1751.140 2475.770 1865.400 ;
        RECT 2479.670 1751.140 2494.370 1865.400 ;
        RECT 2498.270 1751.140 2528.570 1865.400 ;
        RECT 2532.470 1751.140 2547.170 1865.400 ;
        RECT 2551.070 1751.140 2565.770 1865.400 ;
        RECT 2569.670 1751.140 2582.480 1865.400 ;
        RECT 1868.270 1315.400 2582.480 1751.140 ;
        RECT 1868.270 1201.140 1898.570 1315.400 ;
        RECT 1902.470 1201.140 1917.170 1315.400 ;
        RECT 1921.070 1201.140 1935.770 1315.400 ;
        RECT 1939.670 1201.140 1954.370 1315.400 ;
        RECT 1958.270 1201.140 1988.570 1315.400 ;
        RECT 1992.470 1201.140 2007.170 1315.400 ;
        RECT 2011.070 1201.140 2025.770 1315.400 ;
        RECT 2029.670 1201.140 2044.370 1315.400 ;
        RECT 2048.270 1201.140 2078.570 1315.400 ;
        RECT 2082.470 1201.140 2097.170 1315.400 ;
        RECT 2101.070 1201.140 2115.770 1315.400 ;
        RECT 2119.670 1201.140 2134.370 1315.400 ;
        RECT 2138.270 1201.140 2168.570 1315.400 ;
        RECT 2172.470 1201.140 2187.170 1315.400 ;
        RECT 2191.070 1201.140 2205.770 1315.400 ;
        RECT 2209.670 1201.140 2224.370 1315.400 ;
        RECT 2228.270 1201.140 2258.570 1315.400 ;
        RECT 2262.470 1201.140 2277.170 1315.400 ;
        RECT 2281.070 1201.140 2295.770 1315.400 ;
        RECT 2299.670 1201.140 2314.370 1315.400 ;
        RECT 2318.270 1201.140 2348.570 1315.400 ;
        RECT 2352.470 1201.140 2367.170 1315.400 ;
        RECT 2371.070 1201.140 2385.770 1315.400 ;
        RECT 2389.670 1201.140 2404.370 1315.400 ;
        RECT 2408.270 1201.140 2438.570 1315.400 ;
        RECT 2442.470 1201.140 2457.170 1315.400 ;
        RECT 2461.070 1201.140 2475.770 1315.400 ;
        RECT 2479.670 1201.140 2494.370 1315.400 ;
        RECT 2498.270 1201.140 2528.570 1315.400 ;
        RECT 2532.470 1201.140 2547.170 1315.400 ;
        RECT 2551.070 1201.140 2565.770 1315.400 ;
        RECT 2569.670 1201.140 2582.480 1315.400 ;
        RECT 1868.270 765.400 2582.480 1201.140 ;
        RECT 1868.270 651.140 1898.570 765.400 ;
        RECT 1902.470 651.140 1917.170 765.400 ;
        RECT 1921.070 651.140 1935.770 765.400 ;
        RECT 1939.670 651.140 1954.370 765.400 ;
        RECT 1958.270 651.140 1988.570 765.400 ;
        RECT 1992.470 651.140 2007.170 765.400 ;
        RECT 2011.070 651.140 2025.770 765.400 ;
        RECT 2029.670 651.140 2044.370 765.400 ;
        RECT 2048.270 651.140 2078.570 765.400 ;
        RECT 2082.470 651.140 2097.170 765.400 ;
        RECT 2101.070 651.140 2115.770 765.400 ;
        RECT 2119.670 651.140 2134.370 765.400 ;
        RECT 2138.270 651.140 2168.570 765.400 ;
        RECT 2172.470 651.140 2187.170 765.400 ;
        RECT 2191.070 651.140 2205.770 765.400 ;
        RECT 2209.670 651.140 2224.370 765.400 ;
        RECT 2228.270 651.140 2258.570 765.400 ;
        RECT 2262.470 651.140 2277.170 765.400 ;
        RECT 2281.070 651.140 2295.770 765.400 ;
        RECT 2299.670 651.140 2314.370 765.400 ;
        RECT 2318.270 651.140 2348.570 765.400 ;
        RECT 2352.470 651.140 2367.170 765.400 ;
        RECT 2371.070 651.140 2385.770 765.400 ;
        RECT 2389.670 651.140 2404.370 765.400 ;
        RECT 2408.270 651.140 2438.570 765.400 ;
        RECT 2442.470 651.140 2457.170 765.400 ;
        RECT 2461.070 651.140 2475.770 765.400 ;
        RECT 2479.670 651.140 2494.370 765.400 ;
        RECT 2498.270 651.140 2528.570 765.400 ;
        RECT 2532.470 651.140 2547.170 765.400 ;
        RECT 2551.070 651.140 2565.770 765.400 ;
        RECT 2569.670 651.140 2582.480 765.400 ;
        RECT 1868.270 215.400 2582.480 651.140 ;
        RECT 1868.270 199.415 1898.570 215.400 ;
        RECT 1902.470 199.415 1917.170 215.400 ;
        RECT 1921.070 199.415 1935.770 215.400 ;
        RECT 1939.670 199.415 1954.370 215.400 ;
        RECT 1958.270 199.415 1988.570 215.400 ;
        RECT 1992.470 199.415 2007.170 215.400 ;
        RECT 2011.070 199.415 2025.770 215.400 ;
        RECT 2029.670 199.415 2044.370 215.400 ;
        RECT 2048.270 199.415 2078.570 215.400 ;
        RECT 2082.470 199.415 2097.170 215.400 ;
        RECT 2101.070 199.415 2115.770 215.400 ;
        RECT 2119.670 199.415 2134.370 215.400 ;
        RECT 2138.270 199.415 2168.570 215.400 ;
        RECT 2172.470 199.415 2187.170 215.400 ;
        RECT 2191.070 199.415 2205.770 215.400 ;
        RECT 2209.670 199.415 2224.370 215.400 ;
        RECT 2228.270 199.415 2258.570 215.400 ;
        RECT 2262.470 199.415 2277.170 215.400 ;
        RECT 2281.070 199.415 2295.770 215.400 ;
        RECT 2299.670 199.415 2314.370 215.400 ;
        RECT 2318.270 199.415 2348.570 215.400 ;
        RECT 2352.470 199.415 2367.170 215.400 ;
        RECT 2371.070 199.415 2385.770 215.400 ;
        RECT 2389.670 199.415 2404.370 215.400 ;
        RECT 2408.270 199.415 2438.570 215.400 ;
        RECT 2442.470 199.415 2457.170 215.400 ;
        RECT 2461.070 199.415 2475.770 215.400 ;
        RECT 2479.670 199.415 2494.370 215.400 ;
        RECT 2498.270 199.415 2528.570 215.400 ;
        RECT 2532.470 199.415 2547.170 215.400 ;
        RECT 2551.070 199.415 2565.770 215.400 ;
        RECT 2569.670 199.415 2582.480 215.400 ;
  END
END user_project_wrapper
END LIBRARY

