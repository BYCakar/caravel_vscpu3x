* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_sram_2kbyte_1rw1r_32x512_8 abstract view
.subckt sky130_sram_2kbyte_1rw1r_32x512_8 din0[0] din0[1] din0[2] din0[3] din0[4]
+ din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr1[0]
+ addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] addr1[8] csb0 csb1
+ web0 clk0 clk1 wmask0[0] wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[30] dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4]
+ dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13]
+ dout1[14] dout1[15] dout1[16] dout1[17] dout1[18] dout1[19] dout1[20] dout1[21]
+ dout1[22] dout1[23] dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29]
+ dout1[30] dout1[31] vccd1 vssd1
.ends

* Black-box entry subcircuit for VerySimpleCPU_core abstract view
.subckt VerySimpleCPU_core clk done mem_ctrl_addr[0] mem_ctrl_addr[10] mem_ctrl_addr[11]
+ mem_ctrl_addr[12] mem_ctrl_addr[13] mem_ctrl_addr[1] mem_ctrl_addr[2] mem_ctrl_addr[3]
+ mem_ctrl_addr[4] mem_ctrl_addr[5] mem_ctrl_addr[6] mem_ctrl_addr[7] mem_ctrl_addr[8]
+ mem_ctrl_addr[9] mem_ctrl_in[0] mem_ctrl_in[10] mem_ctrl_in[11] mem_ctrl_in[12]
+ mem_ctrl_in[13] mem_ctrl_in[14] mem_ctrl_in[15] mem_ctrl_in[16] mem_ctrl_in[17]
+ mem_ctrl_in[18] mem_ctrl_in[19] mem_ctrl_in[1] mem_ctrl_in[20] mem_ctrl_in[21] mem_ctrl_in[22]
+ mem_ctrl_in[23] mem_ctrl_in[24] mem_ctrl_in[25] mem_ctrl_in[26] mem_ctrl_in[27]
+ mem_ctrl_in[28] mem_ctrl_in[29] mem_ctrl_in[2] mem_ctrl_in[30] mem_ctrl_in[31] mem_ctrl_in[3]
+ mem_ctrl_in[4] mem_ctrl_in[5] mem_ctrl_in[6] mem_ctrl_in[7] mem_ctrl_in[8] mem_ctrl_in[9]
+ mem_ctrl_out[0] mem_ctrl_out[10] mem_ctrl_out[11] mem_ctrl_out[12] mem_ctrl_out[13]
+ mem_ctrl_out[14] mem_ctrl_out[15] mem_ctrl_out[16] mem_ctrl_out[17] mem_ctrl_out[18]
+ mem_ctrl_out[19] mem_ctrl_out[1] mem_ctrl_out[20] mem_ctrl_out[21] mem_ctrl_out[22]
+ mem_ctrl_out[23] mem_ctrl_out[24] mem_ctrl_out[25] mem_ctrl_out[26] mem_ctrl_out[27]
+ mem_ctrl_out[28] mem_ctrl_out[29] mem_ctrl_out[2] mem_ctrl_out[30] mem_ctrl_out[31]
+ mem_ctrl_out[3] mem_ctrl_out[4] mem_ctrl_out[5] mem_ctrl_out[6] mem_ctrl_out[7]
+ mem_ctrl_out[8] mem_ctrl_out[9] mem_ctrl_req mem_ctrl_vld mem_ctrl_we rst vccd1
+ vssd1
.ends

* Black-box entry subcircuit for main_memory abstract view
.subckt main_memory addra[0] addra[1] addra[2] addra[3] addra[4] addra[5] clk dina[0]
+ dina[10] dina[11] dina[12] dina[13] dina[14] dina[15] dina[16] dina[17] dina[18]
+ dina[19] dina[1] dina[20] dina[21] dina[22] dina[23] dina[24] dina[25] dina[26]
+ dina[27] dina[28] dina[29] dina[2] dina[30] dina[31] dina[3] dina[4] dina[5] dina[6]
+ dina[7] dina[8] dina[9] douta[0] douta[10] douta[11] douta[12] douta[13] douta[14]
+ douta[15] douta[16] douta[17] douta[18] douta[19] douta[1] douta[20] douta[21] douta[22]
+ douta[23] douta[24] douta[25] douta[26] douta[27] douta[28] douta[29] douta[2] douta[30]
+ douta[31] douta[3] douta[4] douta[5] douta[6] douta[7] douta[8] douta[9] gpio_in[0]
+ gpio_in[10] gpio_in[1] gpio_in[2] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7]
+ gpio_in[8] gpio_in[9] gpio_out[0] gpio_out[10] gpio_out[1] gpio_out[2] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] vccd1 vssd1
+ wea
.ends

* Black-box entry subcircuit for uart abstract view
.subckt uart clk r_data[0] r_data[1] r_data[2] r_data[3] r_data[4] r_data[5] r_data[6]
+ r_data[7] rd_uart reset rx rx_empty rx_fifo_flush_enable tx tx_full vccd1 vssd1
+ w_data[0] w_data[1] w_data[2] w_data[3] w_data[4] w_data[5] w_data[6] w_data[7]
+ wr_uart
.ends

* Black-box entry subcircuit for main_controller abstract view
.subckt main_controller agent_1_mem_ctrl_addr[0] agent_1_mem_ctrl_addr[10] agent_1_mem_ctrl_addr[11]
+ agent_1_mem_ctrl_addr[12] agent_1_mem_ctrl_addr[13] agent_1_mem_ctrl_addr[1] agent_1_mem_ctrl_addr[2]
+ agent_1_mem_ctrl_addr[3] agent_1_mem_ctrl_addr[4] agent_1_mem_ctrl_addr[5] agent_1_mem_ctrl_addr[6]
+ agent_1_mem_ctrl_addr[7] agent_1_mem_ctrl_addr[8] agent_1_mem_ctrl_addr[9] agent_1_mem_ctrl_in[0]
+ agent_1_mem_ctrl_in[10] agent_1_mem_ctrl_in[11] agent_1_mem_ctrl_in[12] agent_1_mem_ctrl_in[13]
+ agent_1_mem_ctrl_in[14] agent_1_mem_ctrl_in[15] agent_1_mem_ctrl_in[16] agent_1_mem_ctrl_in[17]
+ agent_1_mem_ctrl_in[18] agent_1_mem_ctrl_in[19] agent_1_mem_ctrl_in[1] agent_1_mem_ctrl_in[20]
+ agent_1_mem_ctrl_in[21] agent_1_mem_ctrl_in[22] agent_1_mem_ctrl_in[23] agent_1_mem_ctrl_in[24]
+ agent_1_mem_ctrl_in[25] agent_1_mem_ctrl_in[26] agent_1_mem_ctrl_in[27] agent_1_mem_ctrl_in[28]
+ agent_1_mem_ctrl_in[29] agent_1_mem_ctrl_in[2] agent_1_mem_ctrl_in[30] agent_1_mem_ctrl_in[31]
+ agent_1_mem_ctrl_in[3] agent_1_mem_ctrl_in[4] agent_1_mem_ctrl_in[5] agent_1_mem_ctrl_in[6]
+ agent_1_mem_ctrl_in[7] agent_1_mem_ctrl_in[8] agent_1_mem_ctrl_in[9] agent_1_mem_ctrl_out[0]
+ agent_1_mem_ctrl_out[10] agent_1_mem_ctrl_out[11] agent_1_mem_ctrl_out[12] agent_1_mem_ctrl_out[13]
+ agent_1_mem_ctrl_out[14] agent_1_mem_ctrl_out[15] agent_1_mem_ctrl_out[16] agent_1_mem_ctrl_out[17]
+ agent_1_mem_ctrl_out[18] agent_1_mem_ctrl_out[19] agent_1_mem_ctrl_out[1] agent_1_mem_ctrl_out[20]
+ agent_1_mem_ctrl_out[21] agent_1_mem_ctrl_out[22] agent_1_mem_ctrl_out[23] agent_1_mem_ctrl_out[24]
+ agent_1_mem_ctrl_out[25] agent_1_mem_ctrl_out[26] agent_1_mem_ctrl_out[27] agent_1_mem_ctrl_out[28]
+ agent_1_mem_ctrl_out[29] agent_1_mem_ctrl_out[2] agent_1_mem_ctrl_out[30] agent_1_mem_ctrl_out[31]
+ agent_1_mem_ctrl_out[3] agent_1_mem_ctrl_out[4] agent_1_mem_ctrl_out[5] agent_1_mem_ctrl_out[6]
+ agent_1_mem_ctrl_out[7] agent_1_mem_ctrl_out[8] agent_1_mem_ctrl_out[9] agent_1_mem_ctrl_req
+ agent_1_mem_ctrl_vld agent_1_mem_ctrl_we agent_1_sram0_csb0 agent_1_sram0_dout0[0]
+ agent_1_sram0_dout0[10] agent_1_sram0_dout0[11] agent_1_sram0_dout0[12] agent_1_sram0_dout0[13]
+ agent_1_sram0_dout0[14] agent_1_sram0_dout0[15] agent_1_sram0_dout0[16] agent_1_sram0_dout0[17]
+ agent_1_sram0_dout0[18] agent_1_sram0_dout0[19] agent_1_sram0_dout0[1] agent_1_sram0_dout0[20]
+ agent_1_sram0_dout0[21] agent_1_sram0_dout0[22] agent_1_sram0_dout0[23] agent_1_sram0_dout0[24]
+ agent_1_sram0_dout0[25] agent_1_sram0_dout0[26] agent_1_sram0_dout0[27] agent_1_sram0_dout0[28]
+ agent_1_sram0_dout0[29] agent_1_sram0_dout0[2] agent_1_sram0_dout0[30] agent_1_sram0_dout0[31]
+ agent_1_sram0_dout0[3] agent_1_sram0_dout0[4] agent_1_sram0_dout0[5] agent_1_sram0_dout0[6]
+ agent_1_sram0_dout0[7] agent_1_sram0_dout0[8] agent_1_sram0_dout0[9] agent_1_sram0_web0
+ agent_1_sram1_csb0 agent_1_sram1_dout0[0] agent_1_sram1_dout0[10] agent_1_sram1_dout0[11]
+ agent_1_sram1_dout0[12] agent_1_sram1_dout0[13] agent_1_sram1_dout0[14] agent_1_sram1_dout0[15]
+ agent_1_sram1_dout0[16] agent_1_sram1_dout0[17] agent_1_sram1_dout0[18] agent_1_sram1_dout0[19]
+ agent_1_sram1_dout0[1] agent_1_sram1_dout0[20] agent_1_sram1_dout0[21] agent_1_sram1_dout0[22]
+ agent_1_sram1_dout0[23] agent_1_sram1_dout0[24] agent_1_sram1_dout0[25] agent_1_sram1_dout0[26]
+ agent_1_sram1_dout0[27] agent_1_sram1_dout0[28] agent_1_sram1_dout0[29] agent_1_sram1_dout0[2]
+ agent_1_sram1_dout0[30] agent_1_sram1_dout0[31] agent_1_sram1_dout0[3] agent_1_sram1_dout0[4]
+ agent_1_sram1_dout0[5] agent_1_sram1_dout0[6] agent_1_sram1_dout0[7] agent_1_sram1_dout0[8]
+ agent_1_sram1_dout0[9] agent_1_sram1_web0 agent_1_sram2_csb0 agent_1_sram2_dout0[0]
+ agent_1_sram2_dout0[10] agent_1_sram2_dout0[11] agent_1_sram2_dout0[12] agent_1_sram2_dout0[13]
+ agent_1_sram2_dout0[14] agent_1_sram2_dout0[15] agent_1_sram2_dout0[16] agent_1_sram2_dout0[17]
+ agent_1_sram2_dout0[18] agent_1_sram2_dout0[19] agent_1_sram2_dout0[1] agent_1_sram2_dout0[20]
+ agent_1_sram2_dout0[21] agent_1_sram2_dout0[22] agent_1_sram2_dout0[23] agent_1_sram2_dout0[24]
+ agent_1_sram2_dout0[25] agent_1_sram2_dout0[26] agent_1_sram2_dout0[27] agent_1_sram2_dout0[28]
+ agent_1_sram2_dout0[29] agent_1_sram2_dout0[2] agent_1_sram2_dout0[30] agent_1_sram2_dout0[31]
+ agent_1_sram2_dout0[3] agent_1_sram2_dout0[4] agent_1_sram2_dout0[5] agent_1_sram2_dout0[6]
+ agent_1_sram2_dout0[7] agent_1_sram2_dout0[8] agent_1_sram2_dout0[9] agent_1_sram2_web0
+ agent_1_sram_comm_addr0[0] agent_1_sram_comm_addr0[1] agent_1_sram_comm_addr0[2]
+ agent_1_sram_comm_addr0[3] agent_1_sram_comm_addr0[4] agent_1_sram_comm_addr0[5]
+ agent_1_sram_comm_addr0[6] agent_1_sram_comm_addr0[7] agent_1_sram_comm_addr0[8]
+ agent_1_sram_comm_din0[0] agent_1_sram_comm_din0[10] agent_1_sram_comm_din0[11]
+ agent_1_sram_comm_din0[12] agent_1_sram_comm_din0[13] agent_1_sram_comm_din0[14]
+ agent_1_sram_comm_din0[15] agent_1_sram_comm_din0[16] agent_1_sram_comm_din0[17]
+ agent_1_sram_comm_din0[18] agent_1_sram_comm_din0[19] agent_1_sram_comm_din0[1]
+ agent_1_sram_comm_din0[20] agent_1_sram_comm_din0[21] agent_1_sram_comm_din0[22]
+ agent_1_sram_comm_din0[23] agent_1_sram_comm_din0[24] agent_1_sram_comm_din0[25]
+ agent_1_sram_comm_din0[26] agent_1_sram_comm_din0[27] agent_1_sram_comm_din0[28]
+ agent_1_sram_comm_din0[29] agent_1_sram_comm_din0[2] agent_1_sram_comm_din0[30]
+ agent_1_sram_comm_din0[31] agent_1_sram_comm_din0[3] agent_1_sram_comm_din0[4] agent_1_sram_comm_din0[5]
+ agent_1_sram_comm_din0[6] agent_1_sram_comm_din0[7] agent_1_sram_comm_din0[8] agent_1_sram_comm_din0[9]
+ clk cm_mem_ctrl_addr[0] cm_mem_ctrl_addr[10] cm_mem_ctrl_addr[11] cm_mem_ctrl_addr[12]
+ cm_mem_ctrl_addr[13] cm_mem_ctrl_addr[1] cm_mem_ctrl_addr[2] cm_mem_ctrl_addr[3]
+ cm_mem_ctrl_addr[4] cm_mem_ctrl_addr[5] cm_mem_ctrl_addr[6] cm_mem_ctrl_addr[7]
+ cm_mem_ctrl_addr[8] cm_mem_ctrl_addr[9] cm_mem_ctrl_in[0] cm_mem_ctrl_in[10] cm_mem_ctrl_in[11]
+ cm_mem_ctrl_in[12] cm_mem_ctrl_in[13] cm_mem_ctrl_in[14] cm_mem_ctrl_in[15] cm_mem_ctrl_in[16]
+ cm_mem_ctrl_in[17] cm_mem_ctrl_in[18] cm_mem_ctrl_in[19] cm_mem_ctrl_in[1] cm_mem_ctrl_in[20]
+ cm_mem_ctrl_in[21] cm_mem_ctrl_in[22] cm_mem_ctrl_in[23] cm_mem_ctrl_in[24] cm_mem_ctrl_in[25]
+ cm_mem_ctrl_in[26] cm_mem_ctrl_in[27] cm_mem_ctrl_in[28] cm_mem_ctrl_in[29] cm_mem_ctrl_in[2]
+ cm_mem_ctrl_in[30] cm_mem_ctrl_in[31] cm_mem_ctrl_in[3] cm_mem_ctrl_in[4] cm_mem_ctrl_in[5]
+ cm_mem_ctrl_in[6] cm_mem_ctrl_in[7] cm_mem_ctrl_in[8] cm_mem_ctrl_in[9] cm_mem_ctrl_out[0]
+ cm_mem_ctrl_out[10] cm_mem_ctrl_out[11] cm_mem_ctrl_out[12] cm_mem_ctrl_out[13]
+ cm_mem_ctrl_out[14] cm_mem_ctrl_out[15] cm_mem_ctrl_out[16] cm_mem_ctrl_out[17]
+ cm_mem_ctrl_out[18] cm_mem_ctrl_out[19] cm_mem_ctrl_out[1] cm_mem_ctrl_out[20] cm_mem_ctrl_out[21]
+ cm_mem_ctrl_out[22] cm_mem_ctrl_out[23] cm_mem_ctrl_out[24] cm_mem_ctrl_out[25]
+ cm_mem_ctrl_out[26] cm_mem_ctrl_out[27] cm_mem_ctrl_out[28] cm_mem_ctrl_out[29]
+ cm_mem_ctrl_out[2] cm_mem_ctrl_out[30] cm_mem_ctrl_out[31] cm_mem_ctrl_out[3] cm_mem_ctrl_out[4]
+ cm_mem_ctrl_out[5] cm_mem_ctrl_out[6] cm_mem_ctrl_out[7] cm_mem_ctrl_out[8] cm_mem_ctrl_out[9]
+ cm_mem_ctrl_req cm_mem_ctrl_vld cm_mem_ctrl_we cm_sram0_csb0 cm_sram0_dout0[0] cm_sram0_dout0[10]
+ cm_sram0_dout0[11] cm_sram0_dout0[12] cm_sram0_dout0[13] cm_sram0_dout0[14] cm_sram0_dout0[15]
+ cm_sram0_dout0[16] cm_sram0_dout0[17] cm_sram0_dout0[18] cm_sram0_dout0[19] cm_sram0_dout0[1]
+ cm_sram0_dout0[20] cm_sram0_dout0[21] cm_sram0_dout0[22] cm_sram0_dout0[23] cm_sram0_dout0[24]
+ cm_sram0_dout0[25] cm_sram0_dout0[26] cm_sram0_dout0[27] cm_sram0_dout0[28] cm_sram0_dout0[29]
+ cm_sram0_dout0[2] cm_sram0_dout0[30] cm_sram0_dout0[31] cm_sram0_dout0[3] cm_sram0_dout0[4]
+ cm_sram0_dout0[5] cm_sram0_dout0[6] cm_sram0_dout0[7] cm_sram0_dout0[8] cm_sram0_dout0[9]
+ cm_sram0_web0 cm_sram1_csb0 cm_sram1_dout0[0] cm_sram1_dout0[10] cm_sram1_dout0[11]
+ cm_sram1_dout0[12] cm_sram1_dout0[13] cm_sram1_dout0[14] cm_sram1_dout0[15] cm_sram1_dout0[16]
+ cm_sram1_dout0[17] cm_sram1_dout0[18] cm_sram1_dout0[19] cm_sram1_dout0[1] cm_sram1_dout0[20]
+ cm_sram1_dout0[21] cm_sram1_dout0[22] cm_sram1_dout0[23] cm_sram1_dout0[24] cm_sram1_dout0[25]
+ cm_sram1_dout0[26] cm_sram1_dout0[27] cm_sram1_dout0[28] cm_sram1_dout0[29] cm_sram1_dout0[2]
+ cm_sram1_dout0[30] cm_sram1_dout0[31] cm_sram1_dout0[3] cm_sram1_dout0[4] cm_sram1_dout0[5]
+ cm_sram1_dout0[6] cm_sram1_dout0[7] cm_sram1_dout0[8] cm_sram1_dout0[9] cm_sram1_web0
+ cm_sram2_csb0 cm_sram2_dout0[0] cm_sram2_dout0[10] cm_sram2_dout0[11] cm_sram2_dout0[12]
+ cm_sram2_dout0[13] cm_sram2_dout0[14] cm_sram2_dout0[15] cm_sram2_dout0[16] cm_sram2_dout0[17]
+ cm_sram2_dout0[18] cm_sram2_dout0[19] cm_sram2_dout0[1] cm_sram2_dout0[20] cm_sram2_dout0[21]
+ cm_sram2_dout0[22] cm_sram2_dout0[23] cm_sram2_dout0[24] cm_sram2_dout0[25] cm_sram2_dout0[26]
+ cm_sram2_dout0[27] cm_sram2_dout0[28] cm_sram2_dout0[29] cm_sram2_dout0[2] cm_sram2_dout0[30]
+ cm_sram2_dout0[31] cm_sram2_dout0[3] cm_sram2_dout0[4] cm_sram2_dout0[5] cm_sram2_dout0[6]
+ cm_sram2_dout0[7] cm_sram2_dout0[8] cm_sram2_dout0[9] cm_sram2_web0 cm_sram3_csb0
+ cm_sram3_dout0[0] cm_sram3_dout0[10] cm_sram3_dout0[11] cm_sram3_dout0[12] cm_sram3_dout0[13]
+ cm_sram3_dout0[14] cm_sram3_dout0[15] cm_sram3_dout0[16] cm_sram3_dout0[17] cm_sram3_dout0[18]
+ cm_sram3_dout0[19] cm_sram3_dout0[1] cm_sram3_dout0[20] cm_sram3_dout0[21] cm_sram3_dout0[22]
+ cm_sram3_dout0[23] cm_sram3_dout0[24] cm_sram3_dout0[25] cm_sram3_dout0[26] cm_sram3_dout0[27]
+ cm_sram3_dout0[28] cm_sram3_dout0[29] cm_sram3_dout0[2] cm_sram3_dout0[30] cm_sram3_dout0[31]
+ cm_sram3_dout0[3] cm_sram3_dout0[4] cm_sram3_dout0[5] cm_sram3_dout0[6] cm_sram3_dout0[7]
+ cm_sram3_dout0[8] cm_sram3_dout0[9] cm_sram3_web0 cm_sram_comm_addr0[0] cm_sram_comm_addr0[1]
+ cm_sram_comm_addr0[2] cm_sram_comm_addr0[3] cm_sram_comm_addr0[4] cm_sram_comm_addr0[5]
+ cm_sram_comm_addr0[6] cm_sram_comm_addr0[7] cm_sram_comm_addr0[8] cm_sram_comm_din0[0]
+ cm_sram_comm_din0[10] cm_sram_comm_din0[11] cm_sram_comm_din0[12] cm_sram_comm_din0[13]
+ cm_sram_comm_din0[14] cm_sram_comm_din0[15] cm_sram_comm_din0[16] cm_sram_comm_din0[17]
+ cm_sram_comm_din0[18] cm_sram_comm_din0[19] cm_sram_comm_din0[1] cm_sram_comm_din0[20]
+ cm_sram_comm_din0[21] cm_sram_comm_din0[22] cm_sram_comm_din0[23] cm_sram_comm_din0[24]
+ cm_sram_comm_din0[25] cm_sram_comm_din0[26] cm_sram_comm_din0[27] cm_sram_comm_din0[28]
+ cm_sram_comm_din0[29] cm_sram_comm_din0[2] cm_sram_comm_din0[30] cm_sram_comm_din0[31]
+ cm_sram_comm_din0[3] cm_sram_comm_din0[4] cm_sram_comm_din0[5] cm_sram_comm_din0[6]
+ cm_sram_comm_din0[7] cm_sram_comm_din0[8] cm_sram_comm_din0[9] ct_mem_ctrl_addr[0]
+ ct_mem_ctrl_addr[10] ct_mem_ctrl_addr[11] ct_mem_ctrl_addr[12] ct_mem_ctrl_addr[13]
+ ct_mem_ctrl_addr[1] ct_mem_ctrl_addr[2] ct_mem_ctrl_addr[3] ct_mem_ctrl_addr[4]
+ ct_mem_ctrl_addr[5] ct_mem_ctrl_addr[6] ct_mem_ctrl_addr[7] ct_mem_ctrl_addr[8]
+ ct_mem_ctrl_addr[9] ct_mem_ctrl_in[0] ct_mem_ctrl_in[10] ct_mem_ctrl_in[11] ct_mem_ctrl_in[12]
+ ct_mem_ctrl_in[13] ct_mem_ctrl_in[14] ct_mem_ctrl_in[15] ct_mem_ctrl_in[16] ct_mem_ctrl_in[17]
+ ct_mem_ctrl_in[18] ct_mem_ctrl_in[19] ct_mem_ctrl_in[1] ct_mem_ctrl_in[20] ct_mem_ctrl_in[21]
+ ct_mem_ctrl_in[22] ct_mem_ctrl_in[23] ct_mem_ctrl_in[24] ct_mem_ctrl_in[25] ct_mem_ctrl_in[26]
+ ct_mem_ctrl_in[27] ct_mem_ctrl_in[28] ct_mem_ctrl_in[29] ct_mem_ctrl_in[2] ct_mem_ctrl_in[30]
+ ct_mem_ctrl_in[31] ct_mem_ctrl_in[3] ct_mem_ctrl_in[4] ct_mem_ctrl_in[5] ct_mem_ctrl_in[6]
+ ct_mem_ctrl_in[7] ct_mem_ctrl_in[8] ct_mem_ctrl_in[9] ct_mem_ctrl_out[0] ct_mem_ctrl_out[10]
+ ct_mem_ctrl_out[11] ct_mem_ctrl_out[12] ct_mem_ctrl_out[13] ct_mem_ctrl_out[14]
+ ct_mem_ctrl_out[15] ct_mem_ctrl_out[16] ct_mem_ctrl_out[17] ct_mem_ctrl_out[18]
+ ct_mem_ctrl_out[19] ct_mem_ctrl_out[1] ct_mem_ctrl_out[20] ct_mem_ctrl_out[21] ct_mem_ctrl_out[22]
+ ct_mem_ctrl_out[23] ct_mem_ctrl_out[24] ct_mem_ctrl_out[25] ct_mem_ctrl_out[26]
+ ct_mem_ctrl_out[27] ct_mem_ctrl_out[28] ct_mem_ctrl_out[29] ct_mem_ctrl_out[2] ct_mem_ctrl_out[30]
+ ct_mem_ctrl_out[31] ct_mem_ctrl_out[3] ct_mem_ctrl_out[4] ct_mem_ctrl_out[5] ct_mem_ctrl_out[6]
+ ct_mem_ctrl_out[7] ct_mem_ctrl_out[8] ct_mem_ctrl_out[9] ct_mem_ctrl_req ct_mem_ctrl_vld
+ ct_mem_ctrl_we ct_sram0_csb0 ct_sram0_dout0[0] ct_sram0_dout0[10] ct_sram0_dout0[11]
+ ct_sram0_dout0[12] ct_sram0_dout0[13] ct_sram0_dout0[14] ct_sram0_dout0[15] ct_sram0_dout0[16]
+ ct_sram0_dout0[17] ct_sram0_dout0[18] ct_sram0_dout0[19] ct_sram0_dout0[1] ct_sram0_dout0[20]
+ ct_sram0_dout0[21] ct_sram0_dout0[22] ct_sram0_dout0[23] ct_sram0_dout0[24] ct_sram0_dout0[25]
+ ct_sram0_dout0[26] ct_sram0_dout0[27] ct_sram0_dout0[28] ct_sram0_dout0[29] ct_sram0_dout0[2]
+ ct_sram0_dout0[30] ct_sram0_dout0[31] ct_sram0_dout0[3] ct_sram0_dout0[4] ct_sram0_dout0[5]
+ ct_sram0_dout0[6] ct_sram0_dout0[7] ct_sram0_dout0[8] ct_sram0_dout0[9] ct_sram0_web0
+ ct_sram1_csb0 ct_sram1_dout0[0] ct_sram1_dout0[10] ct_sram1_dout0[11] ct_sram1_dout0[12]
+ ct_sram1_dout0[13] ct_sram1_dout0[14] ct_sram1_dout0[15] ct_sram1_dout0[16] ct_sram1_dout0[17]
+ ct_sram1_dout0[18] ct_sram1_dout0[19] ct_sram1_dout0[1] ct_sram1_dout0[20] ct_sram1_dout0[21]
+ ct_sram1_dout0[22] ct_sram1_dout0[23] ct_sram1_dout0[24] ct_sram1_dout0[25] ct_sram1_dout0[26]
+ ct_sram1_dout0[27] ct_sram1_dout0[28] ct_sram1_dout0[29] ct_sram1_dout0[2] ct_sram1_dout0[30]
+ ct_sram1_dout0[31] ct_sram1_dout0[3] ct_sram1_dout0[4] ct_sram1_dout0[5] ct_sram1_dout0[6]
+ ct_sram1_dout0[7] ct_sram1_dout0[8] ct_sram1_dout0[9] ct_sram1_web0 ct_sram2_csb0
+ ct_sram2_dout0[0] ct_sram2_dout0[10] ct_sram2_dout0[11] ct_sram2_dout0[12] ct_sram2_dout0[13]
+ ct_sram2_dout0[14] ct_sram2_dout0[15] ct_sram2_dout0[16] ct_sram2_dout0[17] ct_sram2_dout0[18]
+ ct_sram2_dout0[19] ct_sram2_dout0[1] ct_sram2_dout0[20] ct_sram2_dout0[21] ct_sram2_dout0[22]
+ ct_sram2_dout0[23] ct_sram2_dout0[24] ct_sram2_dout0[25] ct_sram2_dout0[26] ct_sram2_dout0[27]
+ ct_sram2_dout0[28] ct_sram2_dout0[29] ct_sram2_dout0[2] ct_sram2_dout0[30] ct_sram2_dout0[31]
+ ct_sram2_dout0[3] ct_sram2_dout0[4] ct_sram2_dout0[5] ct_sram2_dout0[6] ct_sram2_dout0[7]
+ ct_sram2_dout0[8] ct_sram2_dout0[9] ct_sram2_web0 ct_sram3_csb0 ct_sram3_dout0[0]
+ ct_sram3_dout0[10] ct_sram3_dout0[11] ct_sram3_dout0[12] ct_sram3_dout0[13] ct_sram3_dout0[14]
+ ct_sram3_dout0[15] ct_sram3_dout0[16] ct_sram3_dout0[17] ct_sram3_dout0[18] ct_sram3_dout0[19]
+ ct_sram3_dout0[1] ct_sram3_dout0[20] ct_sram3_dout0[21] ct_sram3_dout0[22] ct_sram3_dout0[23]
+ ct_sram3_dout0[24] ct_sram3_dout0[25] ct_sram3_dout0[26] ct_sram3_dout0[27] ct_sram3_dout0[28]
+ ct_sram3_dout0[29] ct_sram3_dout0[2] ct_sram3_dout0[30] ct_sram3_dout0[31] ct_sram3_dout0[3]
+ ct_sram3_dout0[4] ct_sram3_dout0[5] ct_sram3_dout0[6] ct_sram3_dout0[7] ct_sram3_dout0[8]
+ ct_sram3_dout0[9] ct_sram3_web0 ct_sram4_csb0 ct_sram4_dout0[0] ct_sram4_dout0[10]
+ ct_sram4_dout0[11] ct_sram4_dout0[12] ct_sram4_dout0[13] ct_sram4_dout0[14] ct_sram4_dout0[15]
+ ct_sram4_dout0[16] ct_sram4_dout0[17] ct_sram4_dout0[18] ct_sram4_dout0[19] ct_sram4_dout0[1]
+ ct_sram4_dout0[20] ct_sram4_dout0[21] ct_sram4_dout0[22] ct_sram4_dout0[23] ct_sram4_dout0[24]
+ ct_sram4_dout0[25] ct_sram4_dout0[26] ct_sram4_dout0[27] ct_sram4_dout0[28] ct_sram4_dout0[29]
+ ct_sram4_dout0[2] ct_sram4_dout0[30] ct_sram4_dout0[31] ct_sram4_dout0[3] ct_sram4_dout0[4]
+ ct_sram4_dout0[5] ct_sram4_dout0[6] ct_sram4_dout0[7] ct_sram4_dout0[8] ct_sram4_dout0[9]
+ ct_sram4_web0 ct_sram_comm_addr0[0] ct_sram_comm_addr0[1] ct_sram_comm_addr0[2]
+ ct_sram_comm_addr0[3] ct_sram_comm_addr0[4] ct_sram_comm_addr0[5] ct_sram_comm_addr0[6]
+ ct_sram_comm_addr0[7] ct_sram_comm_addr0[8] ct_sram_comm_din0[0] ct_sram_comm_din0[10]
+ ct_sram_comm_din0[11] ct_sram_comm_din0[12] ct_sram_comm_din0[13] ct_sram_comm_din0[14]
+ ct_sram_comm_din0[15] ct_sram_comm_din0[16] ct_sram_comm_din0[17] ct_sram_comm_din0[18]
+ ct_sram_comm_din0[19] ct_sram_comm_din0[1] ct_sram_comm_din0[20] ct_sram_comm_din0[21]
+ ct_sram_comm_din0[22] ct_sram_comm_din0[23] ct_sram_comm_din0[24] ct_sram_comm_din0[25]
+ ct_sram_comm_din0[26] ct_sram_comm_din0[27] ct_sram_comm_din0[28] ct_sram_comm_din0[29]
+ ct_sram_comm_din0[2] ct_sram_comm_din0[30] ct_sram_comm_din0[31] ct_sram_comm_din0[3]
+ ct_sram_comm_din0[4] ct_sram_comm_din0[5] ct_sram_comm_din0[6] ct_sram_comm_din0[7]
+ ct_sram_comm_din0[8] ct_sram_comm_din0[9] main_mem_addr[0] main_mem_addr[1] main_mem_addr[2]
+ main_mem_addr[3] main_mem_addr[4] main_mem_addr[5] main_mem_in[0] main_mem_in[10]
+ main_mem_in[11] main_mem_in[12] main_mem_in[13] main_mem_in[14] main_mem_in[15]
+ main_mem_in[16] main_mem_in[17] main_mem_in[18] main_mem_in[19] main_mem_in[1] main_mem_in[20]
+ main_mem_in[21] main_mem_in[22] main_mem_in[23] main_mem_in[24] main_mem_in[25]
+ main_mem_in[26] main_mem_in[27] main_mem_in[28] main_mem_in[29] main_mem_in[2] main_mem_in[30]
+ main_mem_in[31] main_mem_in[3] main_mem_in[4] main_mem_in[5] main_mem_in[6] main_mem_in[7]
+ main_mem_in[8] main_mem_in[9] main_mem_out[0] main_mem_out[10] main_mem_out[11]
+ main_mem_out[12] main_mem_out[13] main_mem_out[14] main_mem_out[15] main_mem_out[16]
+ main_mem_out[17] main_mem_out[18] main_mem_out[19] main_mem_out[1] main_mem_out[20]
+ main_mem_out[21] main_mem_out[22] main_mem_out[23] main_mem_out[24] main_mem_out[25]
+ main_mem_out[26] main_mem_out[27] main_mem_out[28] main_mem_out[29] main_mem_out[2]
+ main_mem_out[30] main_mem_out[31] main_mem_out[3] main_mem_out[4] main_mem_out[5]
+ main_mem_out[6] main_mem_out[7] main_mem_out[8] main_mem_out[9] main_mem_we program_sel[0]
+ program_sel[1] r_data[0] r_data[1] r_data[2] r_data[3] r_data[4] r_data[5] r_data[6]
+ r_data[7] rd_uart rst rst_asserted rx_empty rx_fifo_flush_enable sram_const_addr1[0]
+ sram_const_addr1[1] sram_const_addr1[2] sram_const_addr1[3] sram_const_addr1[4]
+ sram_const_addr1[5] sram_const_addr1[6] sram_const_addr1[7] sram_const_addr1[8]
+ sram_const_csb1 sram_const_wmask0[0] sram_const_wmask0[1] sram_const_wmask0[2] sram_const_wmask0[3]
+ tx_full vccd1 vssd1 w_data[0] w_data[1] w_data[2] w_data[3] w_data[4] w_data[5]
+ w_data[6] w_data[7] wr_uart
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xcodemaker_sram2k_inst1 codemaker_sram2k_inst3/din0[0] codemaker_sram2k_inst3/din0[1]
+ codemaker_sram2k_inst3/din0[2] codemaker_sram2k_inst3/din0[3] codemaker_sram2k_inst3/din0[4]
+ codemaker_sram2k_inst3/din0[5] codemaker_sram2k_inst3/din0[6] codemaker_sram2k_inst3/din0[7]
+ codemaker_sram2k_inst3/din0[8] codemaker_sram2k_inst3/din0[9] codemaker_sram2k_inst3/din0[10]
+ codemaker_sram2k_inst3/din0[11] codemaker_sram2k_inst3/din0[12] codemaker_sram2k_inst3/din0[13]
+ codemaker_sram2k_inst3/din0[14] codemaker_sram2k_inst3/din0[15] codemaker_sram2k_inst3/din0[16]
+ codemaker_sram2k_inst3/din0[17] codemaker_sram2k_inst3/din0[18] codemaker_sram2k_inst3/din0[19]
+ codemaker_sram2k_inst3/din0[20] codemaker_sram2k_inst3/din0[21] codemaker_sram2k_inst3/din0[22]
+ codemaker_sram2k_inst3/din0[23] codemaker_sram2k_inst3/din0[24] codemaker_sram2k_inst3/din0[25]
+ codemaker_sram2k_inst3/din0[26] codemaker_sram2k_inst3/din0[27] codemaker_sram2k_inst3/din0[28]
+ codemaker_sram2k_inst3/din0[29] codemaker_sram2k_inst3/din0[30] codemaker_sram2k_inst3/din0[31]
+ codemaker_sram2k_inst3/addr0[0] codemaker_sram2k_inst3/addr0[1] codemaker_sram2k_inst3/addr0[2]
+ codemaker_sram2k_inst3/addr0[3] codemaker_sram2k_inst3/addr0[4] codemaker_sram2k_inst3/addr0[5]
+ codemaker_sram2k_inst3/addr0[6] codemaker_sram2k_inst3/addr0[7] codemaker_sram2k_inst3/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] codemaker_sram2k_inst1/csb0 agent_1_sram2k_inst2/csb1 codemaker_sram2k_inst1/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] codemaker_sram2k_inst1/dout0[0]
+ codemaker_sram2k_inst1/dout0[1] codemaker_sram2k_inst1/dout0[2] codemaker_sram2k_inst1/dout0[3]
+ codemaker_sram2k_inst1/dout0[4] codemaker_sram2k_inst1/dout0[5] codemaker_sram2k_inst1/dout0[6]
+ codemaker_sram2k_inst1/dout0[7] codemaker_sram2k_inst1/dout0[8] codemaker_sram2k_inst1/dout0[9]
+ codemaker_sram2k_inst1/dout0[10] codemaker_sram2k_inst1/dout0[11] codemaker_sram2k_inst1/dout0[12]
+ codemaker_sram2k_inst1/dout0[13] codemaker_sram2k_inst1/dout0[14] codemaker_sram2k_inst1/dout0[15]
+ codemaker_sram2k_inst1/dout0[16] codemaker_sram2k_inst1/dout0[17] codemaker_sram2k_inst1/dout0[18]
+ codemaker_sram2k_inst1/dout0[19] codemaker_sram2k_inst1/dout0[20] codemaker_sram2k_inst1/dout0[21]
+ codemaker_sram2k_inst1/dout0[22] codemaker_sram2k_inst1/dout0[23] codemaker_sram2k_inst1/dout0[24]
+ codemaker_sram2k_inst1/dout0[25] codemaker_sram2k_inst1/dout0[26] codemaker_sram2k_inst1/dout0[27]
+ codemaker_sram2k_inst1/dout0[28] codemaker_sram2k_inst1/dout0[29] codemaker_sram2k_inst1/dout0[30]
+ codemaker_sram2k_inst1/dout0[31] codemaker_sram2k_inst1/dout1[0] codemaker_sram2k_inst1/dout1[1]
+ codemaker_sram2k_inst1/dout1[2] codemaker_sram2k_inst1/dout1[3] codemaker_sram2k_inst1/dout1[4]
+ codemaker_sram2k_inst1/dout1[5] codemaker_sram2k_inst1/dout1[6] codemaker_sram2k_inst1/dout1[7]
+ codemaker_sram2k_inst1/dout1[8] codemaker_sram2k_inst1/dout1[9] codemaker_sram2k_inst1/dout1[10]
+ codemaker_sram2k_inst1/dout1[11] codemaker_sram2k_inst1/dout1[12] codemaker_sram2k_inst1/dout1[13]
+ codemaker_sram2k_inst1/dout1[14] codemaker_sram2k_inst1/dout1[15] codemaker_sram2k_inst1/dout1[16]
+ codemaker_sram2k_inst1/dout1[17] codemaker_sram2k_inst1/dout1[18] codemaker_sram2k_inst1/dout1[19]
+ codemaker_sram2k_inst1/dout1[20] codemaker_sram2k_inst1/dout1[21] codemaker_sram2k_inst1/dout1[22]
+ codemaker_sram2k_inst1/dout1[23] codemaker_sram2k_inst1/dout1[24] codemaker_sram2k_inst1/dout1[25]
+ codemaker_sram2k_inst1/dout1[26] codemaker_sram2k_inst1/dout1[27] codemaker_sram2k_inst1/dout1[28]
+ codemaker_sram2k_inst1/dout1[29] codemaker_sram2k_inst1/dout1[30] codemaker_sram2k_inst1/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xcodemaker_sram2k_inst0 codemaker_sram2k_inst3/din0[0] codemaker_sram2k_inst3/din0[1]
+ codemaker_sram2k_inst3/din0[2] codemaker_sram2k_inst3/din0[3] codemaker_sram2k_inst3/din0[4]
+ codemaker_sram2k_inst3/din0[5] codemaker_sram2k_inst3/din0[6] codemaker_sram2k_inst3/din0[7]
+ codemaker_sram2k_inst3/din0[8] codemaker_sram2k_inst3/din0[9] codemaker_sram2k_inst3/din0[10]
+ codemaker_sram2k_inst3/din0[11] codemaker_sram2k_inst3/din0[12] codemaker_sram2k_inst3/din0[13]
+ codemaker_sram2k_inst3/din0[14] codemaker_sram2k_inst3/din0[15] codemaker_sram2k_inst3/din0[16]
+ codemaker_sram2k_inst3/din0[17] codemaker_sram2k_inst3/din0[18] codemaker_sram2k_inst3/din0[19]
+ codemaker_sram2k_inst3/din0[20] codemaker_sram2k_inst3/din0[21] codemaker_sram2k_inst3/din0[22]
+ codemaker_sram2k_inst3/din0[23] codemaker_sram2k_inst3/din0[24] codemaker_sram2k_inst3/din0[25]
+ codemaker_sram2k_inst3/din0[26] codemaker_sram2k_inst3/din0[27] codemaker_sram2k_inst3/din0[28]
+ codemaker_sram2k_inst3/din0[29] codemaker_sram2k_inst3/din0[30] codemaker_sram2k_inst3/din0[31]
+ codemaker_sram2k_inst3/addr0[0] codemaker_sram2k_inst3/addr0[1] codemaker_sram2k_inst3/addr0[2]
+ codemaker_sram2k_inst3/addr0[3] codemaker_sram2k_inst3/addr0[4] codemaker_sram2k_inst3/addr0[5]
+ codemaker_sram2k_inst3/addr0[6] codemaker_sram2k_inst3/addr0[7] codemaker_sram2k_inst3/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] codemaker_sram2k_inst0/csb0 agent_1_sram2k_inst2/csb1 codemaker_sram2k_inst0/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] codemaker_sram2k_inst0/dout0[0]
+ codemaker_sram2k_inst0/dout0[1] codemaker_sram2k_inst0/dout0[2] codemaker_sram2k_inst0/dout0[3]
+ codemaker_sram2k_inst0/dout0[4] codemaker_sram2k_inst0/dout0[5] codemaker_sram2k_inst0/dout0[6]
+ codemaker_sram2k_inst0/dout0[7] codemaker_sram2k_inst0/dout0[8] codemaker_sram2k_inst0/dout0[9]
+ codemaker_sram2k_inst0/dout0[10] codemaker_sram2k_inst0/dout0[11] codemaker_sram2k_inst0/dout0[12]
+ codemaker_sram2k_inst0/dout0[13] codemaker_sram2k_inst0/dout0[14] codemaker_sram2k_inst0/dout0[15]
+ codemaker_sram2k_inst0/dout0[16] codemaker_sram2k_inst0/dout0[17] codemaker_sram2k_inst0/dout0[18]
+ codemaker_sram2k_inst0/dout0[19] codemaker_sram2k_inst0/dout0[20] codemaker_sram2k_inst0/dout0[21]
+ codemaker_sram2k_inst0/dout0[22] codemaker_sram2k_inst0/dout0[23] codemaker_sram2k_inst0/dout0[24]
+ codemaker_sram2k_inst0/dout0[25] codemaker_sram2k_inst0/dout0[26] codemaker_sram2k_inst0/dout0[27]
+ codemaker_sram2k_inst0/dout0[28] codemaker_sram2k_inst0/dout0[29] codemaker_sram2k_inst0/dout0[30]
+ codemaker_sram2k_inst0/dout0[31] codemaker_sram2k_inst0/dout1[0] codemaker_sram2k_inst0/dout1[1]
+ codemaker_sram2k_inst0/dout1[2] codemaker_sram2k_inst0/dout1[3] codemaker_sram2k_inst0/dout1[4]
+ codemaker_sram2k_inst0/dout1[5] codemaker_sram2k_inst0/dout1[6] codemaker_sram2k_inst0/dout1[7]
+ codemaker_sram2k_inst0/dout1[8] codemaker_sram2k_inst0/dout1[9] codemaker_sram2k_inst0/dout1[10]
+ codemaker_sram2k_inst0/dout1[11] codemaker_sram2k_inst0/dout1[12] codemaker_sram2k_inst0/dout1[13]
+ codemaker_sram2k_inst0/dout1[14] codemaker_sram2k_inst0/dout1[15] codemaker_sram2k_inst0/dout1[16]
+ codemaker_sram2k_inst0/dout1[17] codemaker_sram2k_inst0/dout1[18] codemaker_sram2k_inst0/dout1[19]
+ codemaker_sram2k_inst0/dout1[20] codemaker_sram2k_inst0/dout1[21] codemaker_sram2k_inst0/dout1[22]
+ codemaker_sram2k_inst0/dout1[23] codemaker_sram2k_inst0/dout1[24] codemaker_sram2k_inst0/dout1[25]
+ codemaker_sram2k_inst0/dout1[26] codemaker_sram2k_inst0/dout1[27] codemaker_sram2k_inst0/dout1[28]
+ codemaker_sram2k_inst0/dout1[29] codemaker_sram2k_inst0/dout1[30] codemaker_sram2k_inst0/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xcontrol_tower_sram2k_inst0 control_tower_sram2k_inst4/din0[0] control_tower_sram2k_inst4/din0[1]
+ control_tower_sram2k_inst4/din0[2] control_tower_sram2k_inst4/din0[3] control_tower_sram2k_inst4/din0[4]
+ control_tower_sram2k_inst4/din0[5] control_tower_sram2k_inst4/din0[6] control_tower_sram2k_inst4/din0[7]
+ control_tower_sram2k_inst4/din0[8] control_tower_sram2k_inst4/din0[9] control_tower_sram2k_inst4/din0[10]
+ control_tower_sram2k_inst4/din0[11] control_tower_sram2k_inst4/din0[12] control_tower_sram2k_inst4/din0[13]
+ control_tower_sram2k_inst4/din0[14] control_tower_sram2k_inst4/din0[15] control_tower_sram2k_inst4/din0[16]
+ control_tower_sram2k_inst4/din0[17] control_tower_sram2k_inst4/din0[18] control_tower_sram2k_inst4/din0[19]
+ control_tower_sram2k_inst4/din0[20] control_tower_sram2k_inst4/din0[21] control_tower_sram2k_inst4/din0[22]
+ control_tower_sram2k_inst4/din0[23] control_tower_sram2k_inst4/din0[24] control_tower_sram2k_inst4/din0[25]
+ control_tower_sram2k_inst4/din0[26] control_tower_sram2k_inst4/din0[27] control_tower_sram2k_inst4/din0[28]
+ control_tower_sram2k_inst4/din0[29] control_tower_sram2k_inst4/din0[30] control_tower_sram2k_inst4/din0[31]
+ control_tower_sram2k_inst4/addr0[0] control_tower_sram2k_inst4/addr0[1] control_tower_sram2k_inst4/addr0[2]
+ control_tower_sram2k_inst4/addr0[3] control_tower_sram2k_inst4/addr0[4] control_tower_sram2k_inst4/addr0[5]
+ control_tower_sram2k_inst4/addr0[6] control_tower_sram2k_inst4/addr0[7] control_tower_sram2k_inst4/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] control_tower_sram2k_inst0/csb0 agent_1_sram2k_inst2/csb1 control_tower_sram2k_inst0/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] control_tower_sram2k_inst0/dout0[0]
+ control_tower_sram2k_inst0/dout0[1] control_tower_sram2k_inst0/dout0[2] control_tower_sram2k_inst0/dout0[3]
+ control_tower_sram2k_inst0/dout0[4] control_tower_sram2k_inst0/dout0[5] control_tower_sram2k_inst0/dout0[6]
+ control_tower_sram2k_inst0/dout0[7] control_tower_sram2k_inst0/dout0[8] control_tower_sram2k_inst0/dout0[9]
+ control_tower_sram2k_inst0/dout0[10] control_tower_sram2k_inst0/dout0[11] control_tower_sram2k_inst0/dout0[12]
+ control_tower_sram2k_inst0/dout0[13] control_tower_sram2k_inst0/dout0[14] control_tower_sram2k_inst0/dout0[15]
+ control_tower_sram2k_inst0/dout0[16] control_tower_sram2k_inst0/dout0[17] control_tower_sram2k_inst0/dout0[18]
+ control_tower_sram2k_inst0/dout0[19] control_tower_sram2k_inst0/dout0[20] control_tower_sram2k_inst0/dout0[21]
+ control_tower_sram2k_inst0/dout0[22] control_tower_sram2k_inst0/dout0[23] control_tower_sram2k_inst0/dout0[24]
+ control_tower_sram2k_inst0/dout0[25] control_tower_sram2k_inst0/dout0[26] control_tower_sram2k_inst0/dout0[27]
+ control_tower_sram2k_inst0/dout0[28] control_tower_sram2k_inst0/dout0[29] control_tower_sram2k_inst0/dout0[30]
+ control_tower_sram2k_inst0/dout0[31] control_tower_sram2k_inst0/dout1[0] control_tower_sram2k_inst0/dout1[1]
+ control_tower_sram2k_inst0/dout1[2] control_tower_sram2k_inst0/dout1[3] control_tower_sram2k_inst0/dout1[4]
+ control_tower_sram2k_inst0/dout1[5] control_tower_sram2k_inst0/dout1[6] control_tower_sram2k_inst0/dout1[7]
+ control_tower_sram2k_inst0/dout1[8] control_tower_sram2k_inst0/dout1[9] control_tower_sram2k_inst0/dout1[10]
+ control_tower_sram2k_inst0/dout1[11] control_tower_sram2k_inst0/dout1[12] control_tower_sram2k_inst0/dout1[13]
+ control_tower_sram2k_inst0/dout1[14] control_tower_sram2k_inst0/dout1[15] control_tower_sram2k_inst0/dout1[16]
+ control_tower_sram2k_inst0/dout1[17] control_tower_sram2k_inst0/dout1[18] control_tower_sram2k_inst0/dout1[19]
+ control_tower_sram2k_inst0/dout1[20] control_tower_sram2k_inst0/dout1[21] control_tower_sram2k_inst0/dout1[22]
+ control_tower_sram2k_inst0/dout1[23] control_tower_sram2k_inst0/dout1[24] control_tower_sram2k_inst0/dout1[25]
+ control_tower_sram2k_inst0/dout1[26] control_tower_sram2k_inst0/dout1[27] control_tower_sram2k_inst0/dout1[28]
+ control_tower_sram2k_inst0/dout1[29] control_tower_sram2k_inst0/dout1[30] control_tower_sram2k_inst0/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xcodemaker_sram2k_inst2 codemaker_sram2k_inst3/din0[0] codemaker_sram2k_inst3/din0[1]
+ codemaker_sram2k_inst3/din0[2] codemaker_sram2k_inst3/din0[3] codemaker_sram2k_inst3/din0[4]
+ codemaker_sram2k_inst3/din0[5] codemaker_sram2k_inst3/din0[6] codemaker_sram2k_inst3/din0[7]
+ codemaker_sram2k_inst3/din0[8] codemaker_sram2k_inst3/din0[9] codemaker_sram2k_inst3/din0[10]
+ codemaker_sram2k_inst3/din0[11] codemaker_sram2k_inst3/din0[12] codemaker_sram2k_inst3/din0[13]
+ codemaker_sram2k_inst3/din0[14] codemaker_sram2k_inst3/din0[15] codemaker_sram2k_inst3/din0[16]
+ codemaker_sram2k_inst3/din0[17] codemaker_sram2k_inst3/din0[18] codemaker_sram2k_inst3/din0[19]
+ codemaker_sram2k_inst3/din0[20] codemaker_sram2k_inst3/din0[21] codemaker_sram2k_inst3/din0[22]
+ codemaker_sram2k_inst3/din0[23] codemaker_sram2k_inst3/din0[24] codemaker_sram2k_inst3/din0[25]
+ codemaker_sram2k_inst3/din0[26] codemaker_sram2k_inst3/din0[27] codemaker_sram2k_inst3/din0[28]
+ codemaker_sram2k_inst3/din0[29] codemaker_sram2k_inst3/din0[30] codemaker_sram2k_inst3/din0[31]
+ codemaker_sram2k_inst3/addr0[0] codemaker_sram2k_inst3/addr0[1] codemaker_sram2k_inst3/addr0[2]
+ codemaker_sram2k_inst3/addr0[3] codemaker_sram2k_inst3/addr0[4] codemaker_sram2k_inst3/addr0[5]
+ codemaker_sram2k_inst3/addr0[6] codemaker_sram2k_inst3/addr0[7] codemaker_sram2k_inst3/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] codemaker_sram2k_inst2/csb0 agent_1_sram2k_inst2/csb1 codemaker_sram2k_inst2/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] codemaker_sram2k_inst2/dout0[0]
+ codemaker_sram2k_inst2/dout0[1] codemaker_sram2k_inst2/dout0[2] codemaker_sram2k_inst2/dout0[3]
+ codemaker_sram2k_inst2/dout0[4] codemaker_sram2k_inst2/dout0[5] codemaker_sram2k_inst2/dout0[6]
+ codemaker_sram2k_inst2/dout0[7] codemaker_sram2k_inst2/dout0[8] codemaker_sram2k_inst2/dout0[9]
+ codemaker_sram2k_inst2/dout0[10] codemaker_sram2k_inst2/dout0[11] codemaker_sram2k_inst2/dout0[12]
+ codemaker_sram2k_inst2/dout0[13] codemaker_sram2k_inst2/dout0[14] codemaker_sram2k_inst2/dout0[15]
+ codemaker_sram2k_inst2/dout0[16] codemaker_sram2k_inst2/dout0[17] codemaker_sram2k_inst2/dout0[18]
+ codemaker_sram2k_inst2/dout0[19] codemaker_sram2k_inst2/dout0[20] codemaker_sram2k_inst2/dout0[21]
+ codemaker_sram2k_inst2/dout0[22] codemaker_sram2k_inst2/dout0[23] codemaker_sram2k_inst2/dout0[24]
+ codemaker_sram2k_inst2/dout0[25] codemaker_sram2k_inst2/dout0[26] codemaker_sram2k_inst2/dout0[27]
+ codemaker_sram2k_inst2/dout0[28] codemaker_sram2k_inst2/dout0[29] codemaker_sram2k_inst2/dout0[30]
+ codemaker_sram2k_inst2/dout0[31] codemaker_sram2k_inst2/dout1[0] codemaker_sram2k_inst2/dout1[1]
+ codemaker_sram2k_inst2/dout1[2] codemaker_sram2k_inst2/dout1[3] codemaker_sram2k_inst2/dout1[4]
+ codemaker_sram2k_inst2/dout1[5] codemaker_sram2k_inst2/dout1[6] codemaker_sram2k_inst2/dout1[7]
+ codemaker_sram2k_inst2/dout1[8] codemaker_sram2k_inst2/dout1[9] codemaker_sram2k_inst2/dout1[10]
+ codemaker_sram2k_inst2/dout1[11] codemaker_sram2k_inst2/dout1[12] codemaker_sram2k_inst2/dout1[13]
+ codemaker_sram2k_inst2/dout1[14] codemaker_sram2k_inst2/dout1[15] codemaker_sram2k_inst2/dout1[16]
+ codemaker_sram2k_inst2/dout1[17] codemaker_sram2k_inst2/dout1[18] codemaker_sram2k_inst2/dout1[19]
+ codemaker_sram2k_inst2/dout1[20] codemaker_sram2k_inst2/dout1[21] codemaker_sram2k_inst2/dout1[22]
+ codemaker_sram2k_inst2/dout1[23] codemaker_sram2k_inst2/dout1[24] codemaker_sram2k_inst2/dout1[25]
+ codemaker_sram2k_inst2/dout1[26] codemaker_sram2k_inst2/dout1[27] codemaker_sram2k_inst2/dout1[28]
+ codemaker_sram2k_inst2/dout1[29] codemaker_sram2k_inst2/dout1[30] codemaker_sram2k_inst2/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xcodemaker_sram2k_inst3 codemaker_sram2k_inst3/din0[0] codemaker_sram2k_inst3/din0[1]
+ codemaker_sram2k_inst3/din0[2] codemaker_sram2k_inst3/din0[3] codemaker_sram2k_inst3/din0[4]
+ codemaker_sram2k_inst3/din0[5] codemaker_sram2k_inst3/din0[6] codemaker_sram2k_inst3/din0[7]
+ codemaker_sram2k_inst3/din0[8] codemaker_sram2k_inst3/din0[9] codemaker_sram2k_inst3/din0[10]
+ codemaker_sram2k_inst3/din0[11] codemaker_sram2k_inst3/din0[12] codemaker_sram2k_inst3/din0[13]
+ codemaker_sram2k_inst3/din0[14] codemaker_sram2k_inst3/din0[15] codemaker_sram2k_inst3/din0[16]
+ codemaker_sram2k_inst3/din0[17] codemaker_sram2k_inst3/din0[18] codemaker_sram2k_inst3/din0[19]
+ codemaker_sram2k_inst3/din0[20] codemaker_sram2k_inst3/din0[21] codemaker_sram2k_inst3/din0[22]
+ codemaker_sram2k_inst3/din0[23] codemaker_sram2k_inst3/din0[24] codemaker_sram2k_inst3/din0[25]
+ codemaker_sram2k_inst3/din0[26] codemaker_sram2k_inst3/din0[27] codemaker_sram2k_inst3/din0[28]
+ codemaker_sram2k_inst3/din0[29] codemaker_sram2k_inst3/din0[30] codemaker_sram2k_inst3/din0[31]
+ codemaker_sram2k_inst3/addr0[0] codemaker_sram2k_inst3/addr0[1] codemaker_sram2k_inst3/addr0[2]
+ codemaker_sram2k_inst3/addr0[3] codemaker_sram2k_inst3/addr0[4] codemaker_sram2k_inst3/addr0[5]
+ codemaker_sram2k_inst3/addr0[6] codemaker_sram2k_inst3/addr0[7] codemaker_sram2k_inst3/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] codemaker_sram2k_inst3/csb0 agent_1_sram2k_inst2/csb1 codemaker_sram2k_inst3/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] codemaker_sram2k_inst3/dout0[0]
+ codemaker_sram2k_inst3/dout0[1] codemaker_sram2k_inst3/dout0[2] codemaker_sram2k_inst3/dout0[3]
+ codemaker_sram2k_inst3/dout0[4] codemaker_sram2k_inst3/dout0[5] codemaker_sram2k_inst3/dout0[6]
+ codemaker_sram2k_inst3/dout0[7] codemaker_sram2k_inst3/dout0[8] codemaker_sram2k_inst3/dout0[9]
+ codemaker_sram2k_inst3/dout0[10] codemaker_sram2k_inst3/dout0[11] codemaker_sram2k_inst3/dout0[12]
+ codemaker_sram2k_inst3/dout0[13] codemaker_sram2k_inst3/dout0[14] codemaker_sram2k_inst3/dout0[15]
+ codemaker_sram2k_inst3/dout0[16] codemaker_sram2k_inst3/dout0[17] codemaker_sram2k_inst3/dout0[18]
+ codemaker_sram2k_inst3/dout0[19] codemaker_sram2k_inst3/dout0[20] codemaker_sram2k_inst3/dout0[21]
+ codemaker_sram2k_inst3/dout0[22] codemaker_sram2k_inst3/dout0[23] codemaker_sram2k_inst3/dout0[24]
+ codemaker_sram2k_inst3/dout0[25] codemaker_sram2k_inst3/dout0[26] codemaker_sram2k_inst3/dout0[27]
+ codemaker_sram2k_inst3/dout0[28] codemaker_sram2k_inst3/dout0[29] codemaker_sram2k_inst3/dout0[30]
+ codemaker_sram2k_inst3/dout0[31] codemaker_sram2k_inst3/dout1[0] codemaker_sram2k_inst3/dout1[1]
+ codemaker_sram2k_inst3/dout1[2] codemaker_sram2k_inst3/dout1[3] codemaker_sram2k_inst3/dout1[4]
+ codemaker_sram2k_inst3/dout1[5] codemaker_sram2k_inst3/dout1[6] codemaker_sram2k_inst3/dout1[7]
+ codemaker_sram2k_inst3/dout1[8] codemaker_sram2k_inst3/dout1[9] codemaker_sram2k_inst3/dout1[10]
+ codemaker_sram2k_inst3/dout1[11] codemaker_sram2k_inst3/dout1[12] codemaker_sram2k_inst3/dout1[13]
+ codemaker_sram2k_inst3/dout1[14] codemaker_sram2k_inst3/dout1[15] codemaker_sram2k_inst3/dout1[16]
+ codemaker_sram2k_inst3/dout1[17] codemaker_sram2k_inst3/dout1[18] codemaker_sram2k_inst3/dout1[19]
+ codemaker_sram2k_inst3/dout1[20] codemaker_sram2k_inst3/dout1[21] codemaker_sram2k_inst3/dout1[22]
+ codemaker_sram2k_inst3/dout1[23] codemaker_sram2k_inst3/dout1[24] codemaker_sram2k_inst3/dout1[25]
+ codemaker_sram2k_inst3/dout1[26] codemaker_sram2k_inst3/dout1[27] codemaker_sram2k_inst3/dout1[28]
+ codemaker_sram2k_inst3/dout1[29] codemaker_sram2k_inst3/dout1[30] codemaker_sram2k_inst3/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xcontrol_tower_sram2k_inst1 control_tower_sram2k_inst4/din0[0] control_tower_sram2k_inst4/din0[1]
+ control_tower_sram2k_inst4/din0[2] control_tower_sram2k_inst4/din0[3] control_tower_sram2k_inst4/din0[4]
+ control_tower_sram2k_inst4/din0[5] control_tower_sram2k_inst4/din0[6] control_tower_sram2k_inst4/din0[7]
+ control_tower_sram2k_inst4/din0[8] control_tower_sram2k_inst4/din0[9] control_tower_sram2k_inst4/din0[10]
+ control_tower_sram2k_inst4/din0[11] control_tower_sram2k_inst4/din0[12] control_tower_sram2k_inst4/din0[13]
+ control_tower_sram2k_inst4/din0[14] control_tower_sram2k_inst4/din0[15] control_tower_sram2k_inst4/din0[16]
+ control_tower_sram2k_inst4/din0[17] control_tower_sram2k_inst4/din0[18] control_tower_sram2k_inst4/din0[19]
+ control_tower_sram2k_inst4/din0[20] control_tower_sram2k_inst4/din0[21] control_tower_sram2k_inst4/din0[22]
+ control_tower_sram2k_inst4/din0[23] control_tower_sram2k_inst4/din0[24] control_tower_sram2k_inst4/din0[25]
+ control_tower_sram2k_inst4/din0[26] control_tower_sram2k_inst4/din0[27] control_tower_sram2k_inst4/din0[28]
+ control_tower_sram2k_inst4/din0[29] control_tower_sram2k_inst4/din0[30] control_tower_sram2k_inst4/din0[31]
+ control_tower_sram2k_inst4/addr0[0] control_tower_sram2k_inst4/addr0[1] control_tower_sram2k_inst4/addr0[2]
+ control_tower_sram2k_inst4/addr0[3] control_tower_sram2k_inst4/addr0[4] control_tower_sram2k_inst4/addr0[5]
+ control_tower_sram2k_inst4/addr0[6] control_tower_sram2k_inst4/addr0[7] control_tower_sram2k_inst4/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] control_tower_sram2k_inst1/csb0 agent_1_sram2k_inst2/csb1 control_tower_sram2k_inst1/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] control_tower_sram2k_inst1/dout0[0]
+ control_tower_sram2k_inst1/dout0[1] control_tower_sram2k_inst1/dout0[2] control_tower_sram2k_inst1/dout0[3]
+ control_tower_sram2k_inst1/dout0[4] control_tower_sram2k_inst1/dout0[5] control_tower_sram2k_inst1/dout0[6]
+ control_tower_sram2k_inst1/dout0[7] control_tower_sram2k_inst1/dout0[8] control_tower_sram2k_inst1/dout0[9]
+ control_tower_sram2k_inst1/dout0[10] control_tower_sram2k_inst1/dout0[11] control_tower_sram2k_inst1/dout0[12]
+ control_tower_sram2k_inst1/dout0[13] control_tower_sram2k_inst1/dout0[14] control_tower_sram2k_inst1/dout0[15]
+ control_tower_sram2k_inst1/dout0[16] control_tower_sram2k_inst1/dout0[17] control_tower_sram2k_inst1/dout0[18]
+ control_tower_sram2k_inst1/dout0[19] control_tower_sram2k_inst1/dout0[20] control_tower_sram2k_inst1/dout0[21]
+ control_tower_sram2k_inst1/dout0[22] control_tower_sram2k_inst1/dout0[23] control_tower_sram2k_inst1/dout0[24]
+ control_tower_sram2k_inst1/dout0[25] control_tower_sram2k_inst1/dout0[26] control_tower_sram2k_inst1/dout0[27]
+ control_tower_sram2k_inst1/dout0[28] control_tower_sram2k_inst1/dout0[29] control_tower_sram2k_inst1/dout0[30]
+ control_tower_sram2k_inst1/dout0[31] control_tower_sram2k_inst1/dout1[0] control_tower_sram2k_inst1/dout1[1]
+ control_tower_sram2k_inst1/dout1[2] control_tower_sram2k_inst1/dout1[3] control_tower_sram2k_inst1/dout1[4]
+ control_tower_sram2k_inst1/dout1[5] control_tower_sram2k_inst1/dout1[6] control_tower_sram2k_inst1/dout1[7]
+ control_tower_sram2k_inst1/dout1[8] control_tower_sram2k_inst1/dout1[9] control_tower_sram2k_inst1/dout1[10]
+ control_tower_sram2k_inst1/dout1[11] control_tower_sram2k_inst1/dout1[12] control_tower_sram2k_inst1/dout1[13]
+ control_tower_sram2k_inst1/dout1[14] control_tower_sram2k_inst1/dout1[15] control_tower_sram2k_inst1/dout1[16]
+ control_tower_sram2k_inst1/dout1[17] control_tower_sram2k_inst1/dout1[18] control_tower_sram2k_inst1/dout1[19]
+ control_tower_sram2k_inst1/dout1[20] control_tower_sram2k_inst1/dout1[21] control_tower_sram2k_inst1/dout1[22]
+ control_tower_sram2k_inst1/dout1[23] control_tower_sram2k_inst1/dout1[24] control_tower_sram2k_inst1/dout1[25]
+ control_tower_sram2k_inst1/dout1[26] control_tower_sram2k_inst1/dout1[27] control_tower_sram2k_inst1/dout1[28]
+ control_tower_sram2k_inst1/dout1[29] control_tower_sram2k_inst1/dout1[30] control_tower_sram2k_inst1/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xcontrol_tower_sram2k_inst2 control_tower_sram2k_inst4/din0[0] control_tower_sram2k_inst4/din0[1]
+ control_tower_sram2k_inst4/din0[2] control_tower_sram2k_inst4/din0[3] control_tower_sram2k_inst4/din0[4]
+ control_tower_sram2k_inst4/din0[5] control_tower_sram2k_inst4/din0[6] control_tower_sram2k_inst4/din0[7]
+ control_tower_sram2k_inst4/din0[8] control_tower_sram2k_inst4/din0[9] control_tower_sram2k_inst4/din0[10]
+ control_tower_sram2k_inst4/din0[11] control_tower_sram2k_inst4/din0[12] control_tower_sram2k_inst4/din0[13]
+ control_tower_sram2k_inst4/din0[14] control_tower_sram2k_inst4/din0[15] control_tower_sram2k_inst4/din0[16]
+ control_tower_sram2k_inst4/din0[17] control_tower_sram2k_inst4/din0[18] control_tower_sram2k_inst4/din0[19]
+ control_tower_sram2k_inst4/din0[20] control_tower_sram2k_inst4/din0[21] control_tower_sram2k_inst4/din0[22]
+ control_tower_sram2k_inst4/din0[23] control_tower_sram2k_inst4/din0[24] control_tower_sram2k_inst4/din0[25]
+ control_tower_sram2k_inst4/din0[26] control_tower_sram2k_inst4/din0[27] control_tower_sram2k_inst4/din0[28]
+ control_tower_sram2k_inst4/din0[29] control_tower_sram2k_inst4/din0[30] control_tower_sram2k_inst4/din0[31]
+ control_tower_sram2k_inst4/addr0[0] control_tower_sram2k_inst4/addr0[1] control_tower_sram2k_inst4/addr0[2]
+ control_tower_sram2k_inst4/addr0[3] control_tower_sram2k_inst4/addr0[4] control_tower_sram2k_inst4/addr0[5]
+ control_tower_sram2k_inst4/addr0[6] control_tower_sram2k_inst4/addr0[7] control_tower_sram2k_inst4/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] control_tower_sram2k_inst2/csb0 agent_1_sram2k_inst2/csb1 control_tower_sram2k_inst2/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] control_tower_sram2k_inst2/dout0[0]
+ control_tower_sram2k_inst2/dout0[1] control_tower_sram2k_inst2/dout0[2] control_tower_sram2k_inst2/dout0[3]
+ control_tower_sram2k_inst2/dout0[4] control_tower_sram2k_inst2/dout0[5] control_tower_sram2k_inst2/dout0[6]
+ control_tower_sram2k_inst2/dout0[7] control_tower_sram2k_inst2/dout0[8] control_tower_sram2k_inst2/dout0[9]
+ control_tower_sram2k_inst2/dout0[10] control_tower_sram2k_inst2/dout0[11] control_tower_sram2k_inst2/dout0[12]
+ control_tower_sram2k_inst2/dout0[13] control_tower_sram2k_inst2/dout0[14] control_tower_sram2k_inst2/dout0[15]
+ control_tower_sram2k_inst2/dout0[16] control_tower_sram2k_inst2/dout0[17] control_tower_sram2k_inst2/dout0[18]
+ control_tower_sram2k_inst2/dout0[19] control_tower_sram2k_inst2/dout0[20] control_tower_sram2k_inst2/dout0[21]
+ control_tower_sram2k_inst2/dout0[22] control_tower_sram2k_inst2/dout0[23] control_tower_sram2k_inst2/dout0[24]
+ control_tower_sram2k_inst2/dout0[25] control_tower_sram2k_inst2/dout0[26] control_tower_sram2k_inst2/dout0[27]
+ control_tower_sram2k_inst2/dout0[28] control_tower_sram2k_inst2/dout0[29] control_tower_sram2k_inst2/dout0[30]
+ control_tower_sram2k_inst2/dout0[31] control_tower_sram2k_inst2/dout1[0] control_tower_sram2k_inst2/dout1[1]
+ control_tower_sram2k_inst2/dout1[2] control_tower_sram2k_inst2/dout1[3] control_tower_sram2k_inst2/dout1[4]
+ control_tower_sram2k_inst2/dout1[5] control_tower_sram2k_inst2/dout1[6] control_tower_sram2k_inst2/dout1[7]
+ control_tower_sram2k_inst2/dout1[8] control_tower_sram2k_inst2/dout1[9] control_tower_sram2k_inst2/dout1[10]
+ control_tower_sram2k_inst2/dout1[11] control_tower_sram2k_inst2/dout1[12] control_tower_sram2k_inst2/dout1[13]
+ control_tower_sram2k_inst2/dout1[14] control_tower_sram2k_inst2/dout1[15] control_tower_sram2k_inst2/dout1[16]
+ control_tower_sram2k_inst2/dout1[17] control_tower_sram2k_inst2/dout1[18] control_tower_sram2k_inst2/dout1[19]
+ control_tower_sram2k_inst2/dout1[20] control_tower_sram2k_inst2/dout1[21] control_tower_sram2k_inst2/dout1[22]
+ control_tower_sram2k_inst2/dout1[23] control_tower_sram2k_inst2/dout1[24] control_tower_sram2k_inst2/dout1[25]
+ control_tower_sram2k_inst2/dout1[26] control_tower_sram2k_inst2/dout1[27] control_tower_sram2k_inst2/dout1[28]
+ control_tower_sram2k_inst2/dout1[29] control_tower_sram2k_inst2/dout1[30] control_tower_sram2k_inst2/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xcontrol_tower_sram2k_inst3 control_tower_sram2k_inst4/din0[0] control_tower_sram2k_inst4/din0[1]
+ control_tower_sram2k_inst4/din0[2] control_tower_sram2k_inst4/din0[3] control_tower_sram2k_inst4/din0[4]
+ control_tower_sram2k_inst4/din0[5] control_tower_sram2k_inst4/din0[6] control_tower_sram2k_inst4/din0[7]
+ control_tower_sram2k_inst4/din0[8] control_tower_sram2k_inst4/din0[9] control_tower_sram2k_inst4/din0[10]
+ control_tower_sram2k_inst4/din0[11] control_tower_sram2k_inst4/din0[12] control_tower_sram2k_inst4/din0[13]
+ control_tower_sram2k_inst4/din0[14] control_tower_sram2k_inst4/din0[15] control_tower_sram2k_inst4/din0[16]
+ control_tower_sram2k_inst4/din0[17] control_tower_sram2k_inst4/din0[18] control_tower_sram2k_inst4/din0[19]
+ control_tower_sram2k_inst4/din0[20] control_tower_sram2k_inst4/din0[21] control_tower_sram2k_inst4/din0[22]
+ control_tower_sram2k_inst4/din0[23] control_tower_sram2k_inst4/din0[24] control_tower_sram2k_inst4/din0[25]
+ control_tower_sram2k_inst4/din0[26] control_tower_sram2k_inst4/din0[27] control_tower_sram2k_inst4/din0[28]
+ control_tower_sram2k_inst4/din0[29] control_tower_sram2k_inst4/din0[30] control_tower_sram2k_inst4/din0[31]
+ control_tower_sram2k_inst4/addr0[0] control_tower_sram2k_inst4/addr0[1] control_tower_sram2k_inst4/addr0[2]
+ control_tower_sram2k_inst4/addr0[3] control_tower_sram2k_inst4/addr0[4] control_tower_sram2k_inst4/addr0[5]
+ control_tower_sram2k_inst4/addr0[6] control_tower_sram2k_inst4/addr0[7] control_tower_sram2k_inst4/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] control_tower_sram2k_inst3/csb0 agent_1_sram2k_inst2/csb1 control_tower_sram2k_inst3/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] control_tower_sram2k_inst3/dout0[0]
+ control_tower_sram2k_inst3/dout0[1] control_tower_sram2k_inst3/dout0[2] control_tower_sram2k_inst3/dout0[3]
+ control_tower_sram2k_inst3/dout0[4] control_tower_sram2k_inst3/dout0[5] control_tower_sram2k_inst3/dout0[6]
+ control_tower_sram2k_inst3/dout0[7] control_tower_sram2k_inst3/dout0[8] control_tower_sram2k_inst3/dout0[9]
+ control_tower_sram2k_inst3/dout0[10] control_tower_sram2k_inst3/dout0[11] control_tower_sram2k_inst3/dout0[12]
+ control_tower_sram2k_inst3/dout0[13] control_tower_sram2k_inst3/dout0[14] control_tower_sram2k_inst3/dout0[15]
+ control_tower_sram2k_inst3/dout0[16] control_tower_sram2k_inst3/dout0[17] control_tower_sram2k_inst3/dout0[18]
+ control_tower_sram2k_inst3/dout0[19] control_tower_sram2k_inst3/dout0[20] control_tower_sram2k_inst3/dout0[21]
+ control_tower_sram2k_inst3/dout0[22] control_tower_sram2k_inst3/dout0[23] control_tower_sram2k_inst3/dout0[24]
+ control_tower_sram2k_inst3/dout0[25] control_tower_sram2k_inst3/dout0[26] control_tower_sram2k_inst3/dout0[27]
+ control_tower_sram2k_inst3/dout0[28] control_tower_sram2k_inst3/dout0[29] control_tower_sram2k_inst3/dout0[30]
+ control_tower_sram2k_inst3/dout0[31] control_tower_sram2k_inst3/dout1[0] control_tower_sram2k_inst3/dout1[1]
+ control_tower_sram2k_inst3/dout1[2] control_tower_sram2k_inst3/dout1[3] control_tower_sram2k_inst3/dout1[4]
+ control_tower_sram2k_inst3/dout1[5] control_tower_sram2k_inst3/dout1[6] control_tower_sram2k_inst3/dout1[7]
+ control_tower_sram2k_inst3/dout1[8] control_tower_sram2k_inst3/dout1[9] control_tower_sram2k_inst3/dout1[10]
+ control_tower_sram2k_inst3/dout1[11] control_tower_sram2k_inst3/dout1[12] control_tower_sram2k_inst3/dout1[13]
+ control_tower_sram2k_inst3/dout1[14] control_tower_sram2k_inst3/dout1[15] control_tower_sram2k_inst3/dout1[16]
+ control_tower_sram2k_inst3/dout1[17] control_tower_sram2k_inst3/dout1[18] control_tower_sram2k_inst3/dout1[19]
+ control_tower_sram2k_inst3/dout1[20] control_tower_sram2k_inst3/dout1[21] control_tower_sram2k_inst3/dout1[22]
+ control_tower_sram2k_inst3/dout1[23] control_tower_sram2k_inst3/dout1[24] control_tower_sram2k_inst3/dout1[25]
+ control_tower_sram2k_inst3/dout1[26] control_tower_sram2k_inst3/dout1[27] control_tower_sram2k_inst3/dout1[28]
+ control_tower_sram2k_inst3/dout1[29] control_tower_sram2k_inst3/dout1[30] control_tower_sram2k_inst3/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xcontrol_tower_sram2k_inst4 control_tower_sram2k_inst4/din0[0] control_tower_sram2k_inst4/din0[1]
+ control_tower_sram2k_inst4/din0[2] control_tower_sram2k_inst4/din0[3] control_tower_sram2k_inst4/din0[4]
+ control_tower_sram2k_inst4/din0[5] control_tower_sram2k_inst4/din0[6] control_tower_sram2k_inst4/din0[7]
+ control_tower_sram2k_inst4/din0[8] control_tower_sram2k_inst4/din0[9] control_tower_sram2k_inst4/din0[10]
+ control_tower_sram2k_inst4/din0[11] control_tower_sram2k_inst4/din0[12] control_tower_sram2k_inst4/din0[13]
+ control_tower_sram2k_inst4/din0[14] control_tower_sram2k_inst4/din0[15] control_tower_sram2k_inst4/din0[16]
+ control_tower_sram2k_inst4/din0[17] control_tower_sram2k_inst4/din0[18] control_tower_sram2k_inst4/din0[19]
+ control_tower_sram2k_inst4/din0[20] control_tower_sram2k_inst4/din0[21] control_tower_sram2k_inst4/din0[22]
+ control_tower_sram2k_inst4/din0[23] control_tower_sram2k_inst4/din0[24] control_tower_sram2k_inst4/din0[25]
+ control_tower_sram2k_inst4/din0[26] control_tower_sram2k_inst4/din0[27] control_tower_sram2k_inst4/din0[28]
+ control_tower_sram2k_inst4/din0[29] control_tower_sram2k_inst4/din0[30] control_tower_sram2k_inst4/din0[31]
+ control_tower_sram2k_inst4/addr0[0] control_tower_sram2k_inst4/addr0[1] control_tower_sram2k_inst4/addr0[2]
+ control_tower_sram2k_inst4/addr0[3] control_tower_sram2k_inst4/addr0[4] control_tower_sram2k_inst4/addr0[5]
+ control_tower_sram2k_inst4/addr0[6] control_tower_sram2k_inst4/addr0[7] control_tower_sram2k_inst4/addr0[8]
+ io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] control_tower_sram2k_inst4/csb0 agent_1_sram2k_inst2/csb1 control_tower_sram2k_inst4/web0
+ wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1]
+ agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3] control_tower_sram2k_inst4/dout0[0]
+ control_tower_sram2k_inst4/dout0[1] control_tower_sram2k_inst4/dout0[2] control_tower_sram2k_inst4/dout0[3]
+ control_tower_sram2k_inst4/dout0[4] control_tower_sram2k_inst4/dout0[5] control_tower_sram2k_inst4/dout0[6]
+ control_tower_sram2k_inst4/dout0[7] control_tower_sram2k_inst4/dout0[8] control_tower_sram2k_inst4/dout0[9]
+ control_tower_sram2k_inst4/dout0[10] control_tower_sram2k_inst4/dout0[11] control_tower_sram2k_inst4/dout0[12]
+ control_tower_sram2k_inst4/dout0[13] control_tower_sram2k_inst4/dout0[14] control_tower_sram2k_inst4/dout0[15]
+ control_tower_sram2k_inst4/dout0[16] control_tower_sram2k_inst4/dout0[17] control_tower_sram2k_inst4/dout0[18]
+ control_tower_sram2k_inst4/dout0[19] control_tower_sram2k_inst4/dout0[20] control_tower_sram2k_inst4/dout0[21]
+ control_tower_sram2k_inst4/dout0[22] control_tower_sram2k_inst4/dout0[23] control_tower_sram2k_inst4/dout0[24]
+ control_tower_sram2k_inst4/dout0[25] control_tower_sram2k_inst4/dout0[26] control_tower_sram2k_inst4/dout0[27]
+ control_tower_sram2k_inst4/dout0[28] control_tower_sram2k_inst4/dout0[29] control_tower_sram2k_inst4/dout0[30]
+ control_tower_sram2k_inst4/dout0[31] control_tower_sram2k_inst4/dout1[0] control_tower_sram2k_inst4/dout1[1]
+ control_tower_sram2k_inst4/dout1[2] control_tower_sram2k_inst4/dout1[3] control_tower_sram2k_inst4/dout1[4]
+ control_tower_sram2k_inst4/dout1[5] control_tower_sram2k_inst4/dout1[6] control_tower_sram2k_inst4/dout1[7]
+ control_tower_sram2k_inst4/dout1[8] control_tower_sram2k_inst4/dout1[9] control_tower_sram2k_inst4/dout1[10]
+ control_tower_sram2k_inst4/dout1[11] control_tower_sram2k_inst4/dout1[12] control_tower_sram2k_inst4/dout1[13]
+ control_tower_sram2k_inst4/dout1[14] control_tower_sram2k_inst4/dout1[15] control_tower_sram2k_inst4/dout1[16]
+ control_tower_sram2k_inst4/dout1[17] control_tower_sram2k_inst4/dout1[18] control_tower_sram2k_inst4/dout1[19]
+ control_tower_sram2k_inst4/dout1[20] control_tower_sram2k_inst4/dout1[21] control_tower_sram2k_inst4/dout1[22]
+ control_tower_sram2k_inst4/dout1[23] control_tower_sram2k_inst4/dout1[24] control_tower_sram2k_inst4/dout1[25]
+ control_tower_sram2k_inst4/dout1[26] control_tower_sram2k_inst4/dout1[27] control_tower_sram2k_inst4/dout1[28]
+ control_tower_sram2k_inst4/dout1[29] control_tower_sram2k_inst4/dout1[30] control_tower_sram2k_inst4/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xinst_codemaker wb_clk_i io_out[13] inst_codemaker/mem_ctrl_addr[0] inst_codemaker/mem_ctrl_addr[10]
+ inst_codemaker/mem_ctrl_addr[11] inst_codemaker/mem_ctrl_addr[12] inst_codemaker/mem_ctrl_addr[13]
+ inst_codemaker/mem_ctrl_addr[1] inst_codemaker/mem_ctrl_addr[2] inst_codemaker/mem_ctrl_addr[3]
+ inst_codemaker/mem_ctrl_addr[4] inst_codemaker/mem_ctrl_addr[5] inst_codemaker/mem_ctrl_addr[6]
+ inst_codemaker/mem_ctrl_addr[7] inst_codemaker/mem_ctrl_addr[8] inst_codemaker/mem_ctrl_addr[9]
+ inst_codemaker/mem_ctrl_in[0] inst_codemaker/mem_ctrl_in[10] inst_codemaker/mem_ctrl_in[11]
+ inst_codemaker/mem_ctrl_in[12] inst_codemaker/mem_ctrl_in[13] inst_codemaker/mem_ctrl_in[14]
+ inst_codemaker/mem_ctrl_in[15] inst_codemaker/mem_ctrl_in[16] inst_codemaker/mem_ctrl_in[17]
+ inst_codemaker/mem_ctrl_in[18] inst_codemaker/mem_ctrl_in[19] inst_codemaker/mem_ctrl_in[1]
+ inst_codemaker/mem_ctrl_in[20] inst_codemaker/mem_ctrl_in[21] inst_codemaker/mem_ctrl_in[22]
+ inst_codemaker/mem_ctrl_in[23] inst_codemaker/mem_ctrl_in[24] inst_codemaker/mem_ctrl_in[25]
+ inst_codemaker/mem_ctrl_in[26] inst_codemaker/mem_ctrl_in[27] inst_codemaker/mem_ctrl_in[28]
+ inst_codemaker/mem_ctrl_in[29] inst_codemaker/mem_ctrl_in[2] inst_codemaker/mem_ctrl_in[30]
+ inst_codemaker/mem_ctrl_in[31] inst_codemaker/mem_ctrl_in[3] inst_codemaker/mem_ctrl_in[4]
+ inst_codemaker/mem_ctrl_in[5] inst_codemaker/mem_ctrl_in[6] inst_codemaker/mem_ctrl_in[7]
+ inst_codemaker/mem_ctrl_in[8] inst_codemaker/mem_ctrl_in[9] inst_codemaker/mem_ctrl_out[0]
+ inst_codemaker/mem_ctrl_out[10] inst_codemaker/mem_ctrl_out[11] inst_codemaker/mem_ctrl_out[12]
+ inst_codemaker/mem_ctrl_out[13] inst_codemaker/mem_ctrl_out[14] inst_codemaker/mem_ctrl_out[15]
+ inst_codemaker/mem_ctrl_out[16] inst_codemaker/mem_ctrl_out[17] inst_codemaker/mem_ctrl_out[18]
+ inst_codemaker/mem_ctrl_out[19] inst_codemaker/mem_ctrl_out[1] inst_codemaker/mem_ctrl_out[20]
+ inst_codemaker/mem_ctrl_out[21] inst_codemaker/mem_ctrl_out[22] inst_codemaker/mem_ctrl_out[23]
+ inst_codemaker/mem_ctrl_out[24] inst_codemaker/mem_ctrl_out[25] inst_codemaker/mem_ctrl_out[26]
+ inst_codemaker/mem_ctrl_out[27] inst_codemaker/mem_ctrl_out[28] inst_codemaker/mem_ctrl_out[29]
+ inst_codemaker/mem_ctrl_out[2] inst_codemaker/mem_ctrl_out[30] inst_codemaker/mem_ctrl_out[31]
+ inst_codemaker/mem_ctrl_out[3] inst_codemaker/mem_ctrl_out[4] inst_codemaker/mem_ctrl_out[5]
+ inst_codemaker/mem_ctrl_out[6] inst_codemaker/mem_ctrl_out[7] inst_codemaker/mem_ctrl_out[8]
+ inst_codemaker/mem_ctrl_out[9] inst_codemaker/mem_ctrl_req inst_codemaker/mem_ctrl_vld
+ inst_codemaker/mem_ctrl_we inst_uart/reset vccd1 vssd1 VerySimpleCPU_core
Xinst_agent_1 wb_clk_i io_out[15] inst_agent_1/mem_ctrl_addr[0] inst_agent_1/mem_ctrl_addr[10]
+ inst_agent_1/mem_ctrl_addr[11] inst_agent_1/mem_ctrl_addr[12] inst_agent_1/mem_ctrl_addr[13]
+ inst_agent_1/mem_ctrl_addr[1] inst_agent_1/mem_ctrl_addr[2] inst_agent_1/mem_ctrl_addr[3]
+ inst_agent_1/mem_ctrl_addr[4] inst_agent_1/mem_ctrl_addr[5] inst_agent_1/mem_ctrl_addr[6]
+ inst_agent_1/mem_ctrl_addr[7] inst_agent_1/mem_ctrl_addr[8] inst_agent_1/mem_ctrl_addr[9]
+ inst_agent_1/mem_ctrl_in[0] inst_agent_1/mem_ctrl_in[10] inst_agent_1/mem_ctrl_in[11]
+ inst_agent_1/mem_ctrl_in[12] inst_agent_1/mem_ctrl_in[13] inst_agent_1/mem_ctrl_in[14]
+ inst_agent_1/mem_ctrl_in[15] inst_agent_1/mem_ctrl_in[16] inst_agent_1/mem_ctrl_in[17]
+ inst_agent_1/mem_ctrl_in[18] inst_agent_1/mem_ctrl_in[19] inst_agent_1/mem_ctrl_in[1]
+ inst_agent_1/mem_ctrl_in[20] inst_agent_1/mem_ctrl_in[21] inst_agent_1/mem_ctrl_in[22]
+ inst_agent_1/mem_ctrl_in[23] inst_agent_1/mem_ctrl_in[24] inst_agent_1/mem_ctrl_in[25]
+ inst_agent_1/mem_ctrl_in[26] inst_agent_1/mem_ctrl_in[27] inst_agent_1/mem_ctrl_in[28]
+ inst_agent_1/mem_ctrl_in[29] inst_agent_1/mem_ctrl_in[2] inst_agent_1/mem_ctrl_in[30]
+ inst_agent_1/mem_ctrl_in[31] inst_agent_1/mem_ctrl_in[3] inst_agent_1/mem_ctrl_in[4]
+ inst_agent_1/mem_ctrl_in[5] inst_agent_1/mem_ctrl_in[6] inst_agent_1/mem_ctrl_in[7]
+ inst_agent_1/mem_ctrl_in[8] inst_agent_1/mem_ctrl_in[9] inst_agent_1/mem_ctrl_out[0]
+ inst_agent_1/mem_ctrl_out[10] inst_agent_1/mem_ctrl_out[11] inst_agent_1/mem_ctrl_out[12]
+ inst_agent_1/mem_ctrl_out[13] inst_agent_1/mem_ctrl_out[14] inst_agent_1/mem_ctrl_out[15]
+ inst_agent_1/mem_ctrl_out[16] inst_agent_1/mem_ctrl_out[17] inst_agent_1/mem_ctrl_out[18]
+ inst_agent_1/mem_ctrl_out[19] inst_agent_1/mem_ctrl_out[1] inst_agent_1/mem_ctrl_out[20]
+ inst_agent_1/mem_ctrl_out[21] inst_agent_1/mem_ctrl_out[22] inst_agent_1/mem_ctrl_out[23]
+ inst_agent_1/mem_ctrl_out[24] inst_agent_1/mem_ctrl_out[25] inst_agent_1/mem_ctrl_out[26]
+ inst_agent_1/mem_ctrl_out[27] inst_agent_1/mem_ctrl_out[28] inst_agent_1/mem_ctrl_out[29]
+ inst_agent_1/mem_ctrl_out[2] inst_agent_1/mem_ctrl_out[30] inst_agent_1/mem_ctrl_out[31]
+ inst_agent_1/mem_ctrl_out[3] inst_agent_1/mem_ctrl_out[4] inst_agent_1/mem_ctrl_out[5]
+ inst_agent_1/mem_ctrl_out[6] inst_agent_1/mem_ctrl_out[7] inst_agent_1/mem_ctrl_out[8]
+ inst_agent_1/mem_ctrl_out[9] inst_agent_1/mem_ctrl_req inst_agent_1/mem_ctrl_vld
+ inst_agent_1/mem_ctrl_we inst_uart/reset vccd1 vssd1 VerySimpleCPU_core
Xagent_1_sram2k_inst0 agent_1_sram2k_inst2/din0[0] agent_1_sram2k_inst2/din0[1] agent_1_sram2k_inst2/din0[2]
+ agent_1_sram2k_inst2/din0[3] agent_1_sram2k_inst2/din0[4] agent_1_sram2k_inst2/din0[5]
+ agent_1_sram2k_inst2/din0[6] agent_1_sram2k_inst2/din0[7] agent_1_sram2k_inst2/din0[8]
+ agent_1_sram2k_inst2/din0[9] agent_1_sram2k_inst2/din0[10] agent_1_sram2k_inst2/din0[11]
+ agent_1_sram2k_inst2/din0[12] agent_1_sram2k_inst2/din0[13] agent_1_sram2k_inst2/din0[14]
+ agent_1_sram2k_inst2/din0[15] agent_1_sram2k_inst2/din0[16] agent_1_sram2k_inst2/din0[17]
+ agent_1_sram2k_inst2/din0[18] agent_1_sram2k_inst2/din0[19] agent_1_sram2k_inst2/din0[20]
+ agent_1_sram2k_inst2/din0[21] agent_1_sram2k_inst2/din0[22] agent_1_sram2k_inst2/din0[23]
+ agent_1_sram2k_inst2/din0[24] agent_1_sram2k_inst2/din0[25] agent_1_sram2k_inst2/din0[26]
+ agent_1_sram2k_inst2/din0[27] agent_1_sram2k_inst2/din0[28] agent_1_sram2k_inst2/din0[29]
+ agent_1_sram2k_inst2/din0[30] agent_1_sram2k_inst2/din0[31] agent_1_sram2k_inst2/addr0[0]
+ agent_1_sram2k_inst2/addr0[1] agent_1_sram2k_inst2/addr0[2] agent_1_sram2k_inst2/addr0[3]
+ agent_1_sram2k_inst2/addr0[4] agent_1_sram2k_inst2/addr0[5] agent_1_sram2k_inst2/addr0[6]
+ agent_1_sram2k_inst2/addr0[7] agent_1_sram2k_inst2/addr0[8] io_oeb[0] io_oeb[1]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] agent_1_sram2k_inst0/csb0
+ agent_1_sram2k_inst2/csb1 agent_1_sram2k_inst0/web0 wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0]
+ agent_1_sram2k_inst2/wmask0[1] agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3]
+ agent_1_sram2k_inst0/dout0[0] agent_1_sram2k_inst0/dout0[1] agent_1_sram2k_inst0/dout0[2]
+ agent_1_sram2k_inst0/dout0[3] agent_1_sram2k_inst0/dout0[4] agent_1_sram2k_inst0/dout0[5]
+ agent_1_sram2k_inst0/dout0[6] agent_1_sram2k_inst0/dout0[7] agent_1_sram2k_inst0/dout0[8]
+ agent_1_sram2k_inst0/dout0[9] agent_1_sram2k_inst0/dout0[10] agent_1_sram2k_inst0/dout0[11]
+ agent_1_sram2k_inst0/dout0[12] agent_1_sram2k_inst0/dout0[13] agent_1_sram2k_inst0/dout0[14]
+ agent_1_sram2k_inst0/dout0[15] agent_1_sram2k_inst0/dout0[16] agent_1_sram2k_inst0/dout0[17]
+ agent_1_sram2k_inst0/dout0[18] agent_1_sram2k_inst0/dout0[19] agent_1_sram2k_inst0/dout0[20]
+ agent_1_sram2k_inst0/dout0[21] agent_1_sram2k_inst0/dout0[22] agent_1_sram2k_inst0/dout0[23]
+ agent_1_sram2k_inst0/dout0[24] agent_1_sram2k_inst0/dout0[25] agent_1_sram2k_inst0/dout0[26]
+ agent_1_sram2k_inst0/dout0[27] agent_1_sram2k_inst0/dout0[28] agent_1_sram2k_inst0/dout0[29]
+ agent_1_sram2k_inst0/dout0[30] agent_1_sram2k_inst0/dout0[31] agent_1_sram2k_inst0/dout1[0]
+ agent_1_sram2k_inst0/dout1[1] agent_1_sram2k_inst0/dout1[2] agent_1_sram2k_inst0/dout1[3]
+ agent_1_sram2k_inst0/dout1[4] agent_1_sram2k_inst0/dout1[5] agent_1_sram2k_inst0/dout1[6]
+ agent_1_sram2k_inst0/dout1[7] agent_1_sram2k_inst0/dout1[8] agent_1_sram2k_inst0/dout1[9]
+ agent_1_sram2k_inst0/dout1[10] agent_1_sram2k_inst0/dout1[11] agent_1_sram2k_inst0/dout1[12]
+ agent_1_sram2k_inst0/dout1[13] agent_1_sram2k_inst0/dout1[14] agent_1_sram2k_inst0/dout1[15]
+ agent_1_sram2k_inst0/dout1[16] agent_1_sram2k_inst0/dout1[17] agent_1_sram2k_inst0/dout1[18]
+ agent_1_sram2k_inst0/dout1[19] agent_1_sram2k_inst0/dout1[20] agent_1_sram2k_inst0/dout1[21]
+ agent_1_sram2k_inst0/dout1[22] agent_1_sram2k_inst0/dout1[23] agent_1_sram2k_inst0/dout1[24]
+ agent_1_sram2k_inst0/dout1[25] agent_1_sram2k_inst0/dout1[26] agent_1_sram2k_inst0/dout1[27]
+ agent_1_sram2k_inst0/dout1[28] agent_1_sram2k_inst0/dout1[29] agent_1_sram2k_inst0/dout1[30]
+ agent_1_sram2k_inst0/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xagent_1_sram2k_inst2 agent_1_sram2k_inst2/din0[0] agent_1_sram2k_inst2/din0[1] agent_1_sram2k_inst2/din0[2]
+ agent_1_sram2k_inst2/din0[3] agent_1_sram2k_inst2/din0[4] agent_1_sram2k_inst2/din0[5]
+ agent_1_sram2k_inst2/din0[6] agent_1_sram2k_inst2/din0[7] agent_1_sram2k_inst2/din0[8]
+ agent_1_sram2k_inst2/din0[9] agent_1_sram2k_inst2/din0[10] agent_1_sram2k_inst2/din0[11]
+ agent_1_sram2k_inst2/din0[12] agent_1_sram2k_inst2/din0[13] agent_1_sram2k_inst2/din0[14]
+ agent_1_sram2k_inst2/din0[15] agent_1_sram2k_inst2/din0[16] agent_1_sram2k_inst2/din0[17]
+ agent_1_sram2k_inst2/din0[18] agent_1_sram2k_inst2/din0[19] agent_1_sram2k_inst2/din0[20]
+ agent_1_sram2k_inst2/din0[21] agent_1_sram2k_inst2/din0[22] agent_1_sram2k_inst2/din0[23]
+ agent_1_sram2k_inst2/din0[24] agent_1_sram2k_inst2/din0[25] agent_1_sram2k_inst2/din0[26]
+ agent_1_sram2k_inst2/din0[27] agent_1_sram2k_inst2/din0[28] agent_1_sram2k_inst2/din0[29]
+ agent_1_sram2k_inst2/din0[30] agent_1_sram2k_inst2/din0[31] agent_1_sram2k_inst2/addr0[0]
+ agent_1_sram2k_inst2/addr0[1] agent_1_sram2k_inst2/addr0[2] agent_1_sram2k_inst2/addr0[3]
+ agent_1_sram2k_inst2/addr0[4] agent_1_sram2k_inst2/addr0[5] agent_1_sram2k_inst2/addr0[6]
+ agent_1_sram2k_inst2/addr0[7] agent_1_sram2k_inst2/addr0[8] io_oeb[0] io_oeb[1]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] agent_1_sram2k_inst2/csb0
+ agent_1_sram2k_inst2/csb1 agent_1_sram2k_inst2/web0 wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0]
+ agent_1_sram2k_inst2/wmask0[1] agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3]
+ agent_1_sram2k_inst2/dout0[0] agent_1_sram2k_inst2/dout0[1] agent_1_sram2k_inst2/dout0[2]
+ agent_1_sram2k_inst2/dout0[3] agent_1_sram2k_inst2/dout0[4] agent_1_sram2k_inst2/dout0[5]
+ agent_1_sram2k_inst2/dout0[6] agent_1_sram2k_inst2/dout0[7] agent_1_sram2k_inst2/dout0[8]
+ agent_1_sram2k_inst2/dout0[9] agent_1_sram2k_inst2/dout0[10] agent_1_sram2k_inst2/dout0[11]
+ agent_1_sram2k_inst2/dout0[12] agent_1_sram2k_inst2/dout0[13] agent_1_sram2k_inst2/dout0[14]
+ agent_1_sram2k_inst2/dout0[15] agent_1_sram2k_inst2/dout0[16] agent_1_sram2k_inst2/dout0[17]
+ agent_1_sram2k_inst2/dout0[18] agent_1_sram2k_inst2/dout0[19] agent_1_sram2k_inst2/dout0[20]
+ agent_1_sram2k_inst2/dout0[21] agent_1_sram2k_inst2/dout0[22] agent_1_sram2k_inst2/dout0[23]
+ agent_1_sram2k_inst2/dout0[24] agent_1_sram2k_inst2/dout0[25] agent_1_sram2k_inst2/dout0[26]
+ agent_1_sram2k_inst2/dout0[27] agent_1_sram2k_inst2/dout0[28] agent_1_sram2k_inst2/dout0[29]
+ agent_1_sram2k_inst2/dout0[30] agent_1_sram2k_inst2/dout0[31] agent_1_sram2k_inst2/dout1[0]
+ agent_1_sram2k_inst2/dout1[1] agent_1_sram2k_inst2/dout1[2] agent_1_sram2k_inst2/dout1[3]
+ agent_1_sram2k_inst2/dout1[4] agent_1_sram2k_inst2/dout1[5] agent_1_sram2k_inst2/dout1[6]
+ agent_1_sram2k_inst2/dout1[7] agent_1_sram2k_inst2/dout1[8] agent_1_sram2k_inst2/dout1[9]
+ agent_1_sram2k_inst2/dout1[10] agent_1_sram2k_inst2/dout1[11] agent_1_sram2k_inst2/dout1[12]
+ agent_1_sram2k_inst2/dout1[13] agent_1_sram2k_inst2/dout1[14] agent_1_sram2k_inst2/dout1[15]
+ agent_1_sram2k_inst2/dout1[16] agent_1_sram2k_inst2/dout1[17] agent_1_sram2k_inst2/dout1[18]
+ agent_1_sram2k_inst2/dout1[19] agent_1_sram2k_inst2/dout1[20] agent_1_sram2k_inst2/dout1[21]
+ agent_1_sram2k_inst2/dout1[22] agent_1_sram2k_inst2/dout1[23] agent_1_sram2k_inst2/dout1[24]
+ agent_1_sram2k_inst2/dout1[25] agent_1_sram2k_inst2/dout1[26] agent_1_sram2k_inst2/dout1[27]
+ agent_1_sram2k_inst2/dout1[28] agent_1_sram2k_inst2/dout1[29] agent_1_sram2k_inst2/dout1[30]
+ agent_1_sram2k_inst2/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xagent_1_sram2k_inst1 agent_1_sram2k_inst2/din0[0] agent_1_sram2k_inst2/din0[1] agent_1_sram2k_inst2/din0[2]
+ agent_1_sram2k_inst2/din0[3] agent_1_sram2k_inst2/din0[4] agent_1_sram2k_inst2/din0[5]
+ agent_1_sram2k_inst2/din0[6] agent_1_sram2k_inst2/din0[7] agent_1_sram2k_inst2/din0[8]
+ agent_1_sram2k_inst2/din0[9] agent_1_sram2k_inst2/din0[10] agent_1_sram2k_inst2/din0[11]
+ agent_1_sram2k_inst2/din0[12] agent_1_sram2k_inst2/din0[13] agent_1_sram2k_inst2/din0[14]
+ agent_1_sram2k_inst2/din0[15] agent_1_sram2k_inst2/din0[16] agent_1_sram2k_inst2/din0[17]
+ agent_1_sram2k_inst2/din0[18] agent_1_sram2k_inst2/din0[19] agent_1_sram2k_inst2/din0[20]
+ agent_1_sram2k_inst2/din0[21] agent_1_sram2k_inst2/din0[22] agent_1_sram2k_inst2/din0[23]
+ agent_1_sram2k_inst2/din0[24] agent_1_sram2k_inst2/din0[25] agent_1_sram2k_inst2/din0[26]
+ agent_1_sram2k_inst2/din0[27] agent_1_sram2k_inst2/din0[28] agent_1_sram2k_inst2/din0[29]
+ agent_1_sram2k_inst2/din0[30] agent_1_sram2k_inst2/din0[31] agent_1_sram2k_inst2/addr0[0]
+ agent_1_sram2k_inst2/addr0[1] agent_1_sram2k_inst2/addr0[2] agent_1_sram2k_inst2/addr0[3]
+ agent_1_sram2k_inst2/addr0[4] agent_1_sram2k_inst2/addr0[5] agent_1_sram2k_inst2/addr0[6]
+ agent_1_sram2k_inst2/addr0[7] agent_1_sram2k_inst2/addr0[8] io_oeb[0] io_oeb[1]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] agent_1_sram2k_inst1/csb0
+ agent_1_sram2k_inst2/csb1 agent_1_sram2k_inst1/web0 wb_clk_i wb_clk_i agent_1_sram2k_inst2/wmask0[0]
+ agent_1_sram2k_inst2/wmask0[1] agent_1_sram2k_inst2/wmask0[2] agent_1_sram2k_inst2/wmask0[3]
+ agent_1_sram2k_inst1/dout0[0] agent_1_sram2k_inst1/dout0[1] agent_1_sram2k_inst1/dout0[2]
+ agent_1_sram2k_inst1/dout0[3] agent_1_sram2k_inst1/dout0[4] agent_1_sram2k_inst1/dout0[5]
+ agent_1_sram2k_inst1/dout0[6] agent_1_sram2k_inst1/dout0[7] agent_1_sram2k_inst1/dout0[8]
+ agent_1_sram2k_inst1/dout0[9] agent_1_sram2k_inst1/dout0[10] agent_1_sram2k_inst1/dout0[11]
+ agent_1_sram2k_inst1/dout0[12] agent_1_sram2k_inst1/dout0[13] agent_1_sram2k_inst1/dout0[14]
+ agent_1_sram2k_inst1/dout0[15] agent_1_sram2k_inst1/dout0[16] agent_1_sram2k_inst1/dout0[17]
+ agent_1_sram2k_inst1/dout0[18] agent_1_sram2k_inst1/dout0[19] agent_1_sram2k_inst1/dout0[20]
+ agent_1_sram2k_inst1/dout0[21] agent_1_sram2k_inst1/dout0[22] agent_1_sram2k_inst1/dout0[23]
+ agent_1_sram2k_inst1/dout0[24] agent_1_sram2k_inst1/dout0[25] agent_1_sram2k_inst1/dout0[26]
+ agent_1_sram2k_inst1/dout0[27] agent_1_sram2k_inst1/dout0[28] agent_1_sram2k_inst1/dout0[29]
+ agent_1_sram2k_inst1/dout0[30] agent_1_sram2k_inst1/dout0[31] agent_1_sram2k_inst1/dout1[0]
+ agent_1_sram2k_inst1/dout1[1] agent_1_sram2k_inst1/dout1[2] agent_1_sram2k_inst1/dout1[3]
+ agent_1_sram2k_inst1/dout1[4] agent_1_sram2k_inst1/dout1[5] agent_1_sram2k_inst1/dout1[6]
+ agent_1_sram2k_inst1/dout1[7] agent_1_sram2k_inst1/dout1[8] agent_1_sram2k_inst1/dout1[9]
+ agent_1_sram2k_inst1/dout1[10] agent_1_sram2k_inst1/dout1[11] agent_1_sram2k_inst1/dout1[12]
+ agent_1_sram2k_inst1/dout1[13] agent_1_sram2k_inst1/dout1[14] agent_1_sram2k_inst1/dout1[15]
+ agent_1_sram2k_inst1/dout1[16] agent_1_sram2k_inst1/dout1[17] agent_1_sram2k_inst1/dout1[18]
+ agent_1_sram2k_inst1/dout1[19] agent_1_sram2k_inst1/dout1[20] agent_1_sram2k_inst1/dout1[21]
+ agent_1_sram2k_inst1/dout1[22] agent_1_sram2k_inst1/dout1[23] agent_1_sram2k_inst1/dout1[24]
+ agent_1_sram2k_inst1/dout1[25] agent_1_sram2k_inst1/dout1[26] agent_1_sram2k_inst1/dout1[27]
+ agent_1_sram2k_inst1/dout1[28] agent_1_sram2k_inst1/dout1[29] agent_1_sram2k_inst1/dout1[30]
+ agent_1_sram2k_inst1/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xinst_control_tower wb_clk_i io_out[14] inst_control_tower/mem_ctrl_addr[0] inst_control_tower/mem_ctrl_addr[10]
+ inst_control_tower/mem_ctrl_addr[11] inst_control_tower/mem_ctrl_addr[12] inst_control_tower/mem_ctrl_addr[13]
+ inst_control_tower/mem_ctrl_addr[1] inst_control_tower/mem_ctrl_addr[2] inst_control_tower/mem_ctrl_addr[3]
+ inst_control_tower/mem_ctrl_addr[4] inst_control_tower/mem_ctrl_addr[5] inst_control_tower/mem_ctrl_addr[6]
+ inst_control_tower/mem_ctrl_addr[7] inst_control_tower/mem_ctrl_addr[8] inst_control_tower/mem_ctrl_addr[9]
+ inst_control_tower/mem_ctrl_in[0] inst_control_tower/mem_ctrl_in[10] inst_control_tower/mem_ctrl_in[11]
+ inst_control_tower/mem_ctrl_in[12] inst_control_tower/mem_ctrl_in[13] inst_control_tower/mem_ctrl_in[14]
+ inst_control_tower/mem_ctrl_in[15] inst_control_tower/mem_ctrl_in[16] inst_control_tower/mem_ctrl_in[17]
+ inst_control_tower/mem_ctrl_in[18] inst_control_tower/mem_ctrl_in[19] inst_control_tower/mem_ctrl_in[1]
+ inst_control_tower/mem_ctrl_in[20] inst_control_tower/mem_ctrl_in[21] inst_control_tower/mem_ctrl_in[22]
+ inst_control_tower/mem_ctrl_in[23] inst_control_tower/mem_ctrl_in[24] inst_control_tower/mem_ctrl_in[25]
+ inst_control_tower/mem_ctrl_in[26] inst_control_tower/mem_ctrl_in[27] inst_control_tower/mem_ctrl_in[28]
+ inst_control_tower/mem_ctrl_in[29] inst_control_tower/mem_ctrl_in[2] inst_control_tower/mem_ctrl_in[30]
+ inst_control_tower/mem_ctrl_in[31] inst_control_tower/mem_ctrl_in[3] inst_control_tower/mem_ctrl_in[4]
+ inst_control_tower/mem_ctrl_in[5] inst_control_tower/mem_ctrl_in[6] inst_control_tower/mem_ctrl_in[7]
+ inst_control_tower/mem_ctrl_in[8] inst_control_tower/mem_ctrl_in[9] inst_control_tower/mem_ctrl_out[0]
+ inst_control_tower/mem_ctrl_out[10] inst_control_tower/mem_ctrl_out[11] inst_control_tower/mem_ctrl_out[12]
+ inst_control_tower/mem_ctrl_out[13] inst_control_tower/mem_ctrl_out[14] inst_control_tower/mem_ctrl_out[15]
+ inst_control_tower/mem_ctrl_out[16] inst_control_tower/mem_ctrl_out[17] inst_control_tower/mem_ctrl_out[18]
+ inst_control_tower/mem_ctrl_out[19] inst_control_tower/mem_ctrl_out[1] inst_control_tower/mem_ctrl_out[20]
+ inst_control_tower/mem_ctrl_out[21] inst_control_tower/mem_ctrl_out[22] inst_control_tower/mem_ctrl_out[23]
+ inst_control_tower/mem_ctrl_out[24] inst_control_tower/mem_ctrl_out[25] inst_control_tower/mem_ctrl_out[26]
+ inst_control_tower/mem_ctrl_out[27] inst_control_tower/mem_ctrl_out[28] inst_control_tower/mem_ctrl_out[29]
+ inst_control_tower/mem_ctrl_out[2] inst_control_tower/mem_ctrl_out[30] inst_control_tower/mem_ctrl_out[31]
+ inst_control_tower/mem_ctrl_out[3] inst_control_tower/mem_ctrl_out[4] inst_control_tower/mem_ctrl_out[5]
+ inst_control_tower/mem_ctrl_out[6] inst_control_tower/mem_ctrl_out[7] inst_control_tower/mem_ctrl_out[8]
+ inst_control_tower/mem_ctrl_out[9] inst_control_tower/mem_ctrl_req inst_control_tower/mem_ctrl_vld
+ inst_control_tower/mem_ctrl_we inst_uart/reset vccd1 vssd1 VerySimpleCPU_core
Xinst_main_memory inst_main_memory/addra[0] inst_main_memory/addra[1] inst_main_memory/addra[2]
+ inst_main_memory/addra[3] inst_main_memory/addra[4] inst_main_memory/addra[5] wb_clk_i
+ inst_main_memory/dina[0] inst_main_memory/dina[10] inst_main_memory/dina[11] inst_main_memory/dina[12]
+ inst_main_memory/dina[13] inst_main_memory/dina[14] inst_main_memory/dina[15] inst_main_memory/dina[16]
+ inst_main_memory/dina[17] inst_main_memory/dina[18] inst_main_memory/dina[19] inst_main_memory/dina[1]
+ inst_main_memory/dina[20] inst_main_memory/dina[21] inst_main_memory/dina[22] inst_main_memory/dina[23]
+ inst_main_memory/dina[24] inst_main_memory/dina[25] inst_main_memory/dina[26] inst_main_memory/dina[27]
+ inst_main_memory/dina[28] inst_main_memory/dina[29] inst_main_memory/dina[2] inst_main_memory/dina[30]
+ inst_main_memory/dina[31] inst_main_memory/dina[3] inst_main_memory/dina[4] inst_main_memory/dina[5]
+ inst_main_memory/dina[6] inst_main_memory/dina[7] inst_main_memory/dina[8] inst_main_memory/dina[9]
+ inst_main_memory/douta[0] inst_main_memory/douta[10] inst_main_memory/douta[11]
+ inst_main_memory/douta[12] inst_main_memory/douta[13] inst_main_memory/douta[14]
+ inst_main_memory/douta[15] inst_main_memory/douta[16] inst_main_memory/douta[17]
+ inst_main_memory/douta[18] inst_main_memory/douta[19] inst_main_memory/douta[1]
+ inst_main_memory/douta[20] inst_main_memory/douta[21] inst_main_memory/douta[22]
+ inst_main_memory/douta[23] inst_main_memory/douta[24] inst_main_memory/douta[25]
+ inst_main_memory/douta[26] inst_main_memory/douta[27] inst_main_memory/douta[28]
+ inst_main_memory/douta[29] inst_main_memory/douta[2] inst_main_memory/douta[30]
+ inst_main_memory/douta[31] inst_main_memory/douta[3] inst_main_memory/douta[4] inst_main_memory/douta[5]
+ inst_main_memory/douta[6] inst_main_memory/douta[7] inst_main_memory/douta[8] inst_main_memory/douta[9]
+ io_in[16] io_in[26] io_in[17] io_in[18] io_in[19] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_out[27] io_out[37] io_out[28] io_out[29] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] vccd1 vssd1 inst_main_memory/wea
+ main_memory
Xinst_uart wb_clk_i inst_uart/r_data[0] inst_uart/r_data[1] inst_uart/r_data[2] inst_uart/r_data[3]
+ inst_uart/r_data[4] inst_uart/r_data[5] inst_uart/r_data[6] inst_uart/r_data[7]
+ inst_uart/rd_uart inst_uart/reset io_in[11] inst_uart/rx_empty inst_uart/rx_fifo_flush_enable
+ io_out[12] inst_uart/tx_full vccd1 vssd1 inst_uart/w_data[0] inst_uart/w_data[1]
+ inst_uart/w_data[2] inst_uart/w_data[3] inst_uart/w_data[4] inst_uart/w_data[5]
+ inst_uart/w_data[6] inst_uart/w_data[7] inst_uart/wr_uart uart
Xinst_main_controller inst_agent_1/mem_ctrl_addr[0] inst_agent_1/mem_ctrl_addr[10]
+ inst_agent_1/mem_ctrl_addr[11] inst_agent_1/mem_ctrl_addr[12] inst_agent_1/mem_ctrl_addr[13]
+ inst_agent_1/mem_ctrl_addr[1] inst_agent_1/mem_ctrl_addr[2] inst_agent_1/mem_ctrl_addr[3]
+ inst_agent_1/mem_ctrl_addr[4] inst_agent_1/mem_ctrl_addr[5] inst_agent_1/mem_ctrl_addr[6]
+ inst_agent_1/mem_ctrl_addr[7] inst_agent_1/mem_ctrl_addr[8] inst_agent_1/mem_ctrl_addr[9]
+ inst_agent_1/mem_ctrl_in[0] inst_agent_1/mem_ctrl_in[10] inst_agent_1/mem_ctrl_in[11]
+ inst_agent_1/mem_ctrl_in[12] inst_agent_1/mem_ctrl_in[13] inst_agent_1/mem_ctrl_in[14]
+ inst_agent_1/mem_ctrl_in[15] inst_agent_1/mem_ctrl_in[16] inst_agent_1/mem_ctrl_in[17]
+ inst_agent_1/mem_ctrl_in[18] inst_agent_1/mem_ctrl_in[19] inst_agent_1/mem_ctrl_in[1]
+ inst_agent_1/mem_ctrl_in[20] inst_agent_1/mem_ctrl_in[21] inst_agent_1/mem_ctrl_in[22]
+ inst_agent_1/mem_ctrl_in[23] inst_agent_1/mem_ctrl_in[24] inst_agent_1/mem_ctrl_in[25]
+ inst_agent_1/mem_ctrl_in[26] inst_agent_1/mem_ctrl_in[27] inst_agent_1/mem_ctrl_in[28]
+ inst_agent_1/mem_ctrl_in[29] inst_agent_1/mem_ctrl_in[2] inst_agent_1/mem_ctrl_in[30]
+ inst_agent_1/mem_ctrl_in[31] inst_agent_1/mem_ctrl_in[3] inst_agent_1/mem_ctrl_in[4]
+ inst_agent_1/mem_ctrl_in[5] inst_agent_1/mem_ctrl_in[6] inst_agent_1/mem_ctrl_in[7]
+ inst_agent_1/mem_ctrl_in[8] inst_agent_1/mem_ctrl_in[9] inst_agent_1/mem_ctrl_out[0]
+ inst_agent_1/mem_ctrl_out[10] inst_agent_1/mem_ctrl_out[11] inst_agent_1/mem_ctrl_out[12]
+ inst_agent_1/mem_ctrl_out[13] inst_agent_1/mem_ctrl_out[14] inst_agent_1/mem_ctrl_out[15]
+ inst_agent_1/mem_ctrl_out[16] inst_agent_1/mem_ctrl_out[17] inst_agent_1/mem_ctrl_out[18]
+ inst_agent_1/mem_ctrl_out[19] inst_agent_1/mem_ctrl_out[1] inst_agent_1/mem_ctrl_out[20]
+ inst_agent_1/mem_ctrl_out[21] inst_agent_1/mem_ctrl_out[22] inst_agent_1/mem_ctrl_out[23]
+ inst_agent_1/mem_ctrl_out[24] inst_agent_1/mem_ctrl_out[25] inst_agent_1/mem_ctrl_out[26]
+ inst_agent_1/mem_ctrl_out[27] inst_agent_1/mem_ctrl_out[28] inst_agent_1/mem_ctrl_out[29]
+ inst_agent_1/mem_ctrl_out[2] inst_agent_1/mem_ctrl_out[30] inst_agent_1/mem_ctrl_out[31]
+ inst_agent_1/mem_ctrl_out[3] inst_agent_1/mem_ctrl_out[4] inst_agent_1/mem_ctrl_out[5]
+ inst_agent_1/mem_ctrl_out[6] inst_agent_1/mem_ctrl_out[7] inst_agent_1/mem_ctrl_out[8]
+ inst_agent_1/mem_ctrl_out[9] inst_agent_1/mem_ctrl_req inst_agent_1/mem_ctrl_vld
+ inst_agent_1/mem_ctrl_we agent_1_sram2k_inst0/csb0 agent_1_sram2k_inst0/dout0[0]
+ agent_1_sram2k_inst0/dout0[10] agent_1_sram2k_inst0/dout0[11] agent_1_sram2k_inst0/dout0[12]
+ agent_1_sram2k_inst0/dout0[13] agent_1_sram2k_inst0/dout0[14] agent_1_sram2k_inst0/dout0[15]
+ agent_1_sram2k_inst0/dout0[16] agent_1_sram2k_inst0/dout0[17] agent_1_sram2k_inst0/dout0[18]
+ agent_1_sram2k_inst0/dout0[19] agent_1_sram2k_inst0/dout0[1] agent_1_sram2k_inst0/dout0[20]
+ agent_1_sram2k_inst0/dout0[21] agent_1_sram2k_inst0/dout0[22] agent_1_sram2k_inst0/dout0[23]
+ agent_1_sram2k_inst0/dout0[24] agent_1_sram2k_inst0/dout0[25] agent_1_sram2k_inst0/dout0[26]
+ agent_1_sram2k_inst0/dout0[27] agent_1_sram2k_inst0/dout0[28] agent_1_sram2k_inst0/dout0[29]
+ agent_1_sram2k_inst0/dout0[2] agent_1_sram2k_inst0/dout0[30] agent_1_sram2k_inst0/dout0[31]
+ agent_1_sram2k_inst0/dout0[3] agent_1_sram2k_inst0/dout0[4] agent_1_sram2k_inst0/dout0[5]
+ agent_1_sram2k_inst0/dout0[6] agent_1_sram2k_inst0/dout0[7] agent_1_sram2k_inst0/dout0[8]
+ agent_1_sram2k_inst0/dout0[9] agent_1_sram2k_inst0/web0 agent_1_sram2k_inst1/csb0
+ agent_1_sram2k_inst1/dout0[0] agent_1_sram2k_inst1/dout0[10] agent_1_sram2k_inst1/dout0[11]
+ agent_1_sram2k_inst1/dout0[12] agent_1_sram2k_inst1/dout0[13] agent_1_sram2k_inst1/dout0[14]
+ agent_1_sram2k_inst1/dout0[15] agent_1_sram2k_inst1/dout0[16] agent_1_sram2k_inst1/dout0[17]
+ agent_1_sram2k_inst1/dout0[18] agent_1_sram2k_inst1/dout0[19] agent_1_sram2k_inst1/dout0[1]
+ agent_1_sram2k_inst1/dout0[20] agent_1_sram2k_inst1/dout0[21] agent_1_sram2k_inst1/dout0[22]
+ agent_1_sram2k_inst1/dout0[23] agent_1_sram2k_inst1/dout0[24] agent_1_sram2k_inst1/dout0[25]
+ agent_1_sram2k_inst1/dout0[26] agent_1_sram2k_inst1/dout0[27] agent_1_sram2k_inst1/dout0[28]
+ agent_1_sram2k_inst1/dout0[29] agent_1_sram2k_inst1/dout0[2] agent_1_sram2k_inst1/dout0[30]
+ agent_1_sram2k_inst1/dout0[31] agent_1_sram2k_inst1/dout0[3] agent_1_sram2k_inst1/dout0[4]
+ agent_1_sram2k_inst1/dout0[5] agent_1_sram2k_inst1/dout0[6] agent_1_sram2k_inst1/dout0[7]
+ agent_1_sram2k_inst1/dout0[8] agent_1_sram2k_inst1/dout0[9] agent_1_sram2k_inst1/web0
+ agent_1_sram2k_inst2/csb0 agent_1_sram2k_inst2/dout0[0] agent_1_sram2k_inst2/dout0[10]
+ agent_1_sram2k_inst2/dout0[11] agent_1_sram2k_inst2/dout0[12] agent_1_sram2k_inst2/dout0[13]
+ agent_1_sram2k_inst2/dout0[14] agent_1_sram2k_inst2/dout0[15] agent_1_sram2k_inst2/dout0[16]
+ agent_1_sram2k_inst2/dout0[17] agent_1_sram2k_inst2/dout0[18] agent_1_sram2k_inst2/dout0[19]
+ agent_1_sram2k_inst2/dout0[1] agent_1_sram2k_inst2/dout0[20] agent_1_sram2k_inst2/dout0[21]
+ agent_1_sram2k_inst2/dout0[22] agent_1_sram2k_inst2/dout0[23] agent_1_sram2k_inst2/dout0[24]
+ agent_1_sram2k_inst2/dout0[25] agent_1_sram2k_inst2/dout0[26] agent_1_sram2k_inst2/dout0[27]
+ agent_1_sram2k_inst2/dout0[28] agent_1_sram2k_inst2/dout0[29] agent_1_sram2k_inst2/dout0[2]
+ agent_1_sram2k_inst2/dout0[30] agent_1_sram2k_inst2/dout0[31] agent_1_sram2k_inst2/dout0[3]
+ agent_1_sram2k_inst2/dout0[4] agent_1_sram2k_inst2/dout0[5] agent_1_sram2k_inst2/dout0[6]
+ agent_1_sram2k_inst2/dout0[7] agent_1_sram2k_inst2/dout0[8] agent_1_sram2k_inst2/dout0[9]
+ agent_1_sram2k_inst2/web0 agent_1_sram2k_inst2/addr0[0] agent_1_sram2k_inst2/addr0[1]
+ agent_1_sram2k_inst2/addr0[2] agent_1_sram2k_inst2/addr0[3] agent_1_sram2k_inst2/addr0[4]
+ agent_1_sram2k_inst2/addr0[5] agent_1_sram2k_inst2/addr0[6] agent_1_sram2k_inst2/addr0[7]
+ agent_1_sram2k_inst2/addr0[8] agent_1_sram2k_inst2/din0[0] agent_1_sram2k_inst2/din0[10]
+ agent_1_sram2k_inst2/din0[11] agent_1_sram2k_inst2/din0[12] agent_1_sram2k_inst2/din0[13]
+ agent_1_sram2k_inst2/din0[14] agent_1_sram2k_inst2/din0[15] agent_1_sram2k_inst2/din0[16]
+ agent_1_sram2k_inst2/din0[17] agent_1_sram2k_inst2/din0[18] agent_1_sram2k_inst2/din0[19]
+ agent_1_sram2k_inst2/din0[1] agent_1_sram2k_inst2/din0[20] agent_1_sram2k_inst2/din0[21]
+ agent_1_sram2k_inst2/din0[22] agent_1_sram2k_inst2/din0[23] agent_1_sram2k_inst2/din0[24]
+ agent_1_sram2k_inst2/din0[25] agent_1_sram2k_inst2/din0[26] agent_1_sram2k_inst2/din0[27]
+ agent_1_sram2k_inst2/din0[28] agent_1_sram2k_inst2/din0[29] agent_1_sram2k_inst2/din0[2]
+ agent_1_sram2k_inst2/din0[30] agent_1_sram2k_inst2/din0[31] agent_1_sram2k_inst2/din0[3]
+ agent_1_sram2k_inst2/din0[4] agent_1_sram2k_inst2/din0[5] agent_1_sram2k_inst2/din0[6]
+ agent_1_sram2k_inst2/din0[7] agent_1_sram2k_inst2/din0[8] agent_1_sram2k_inst2/din0[9]
+ wb_clk_i inst_codemaker/mem_ctrl_addr[0] inst_codemaker/mem_ctrl_addr[10] inst_codemaker/mem_ctrl_addr[11]
+ inst_codemaker/mem_ctrl_addr[12] inst_codemaker/mem_ctrl_addr[13] inst_codemaker/mem_ctrl_addr[1]
+ inst_codemaker/mem_ctrl_addr[2] inst_codemaker/mem_ctrl_addr[3] inst_codemaker/mem_ctrl_addr[4]
+ inst_codemaker/mem_ctrl_addr[5] inst_codemaker/mem_ctrl_addr[6] inst_codemaker/mem_ctrl_addr[7]
+ inst_codemaker/mem_ctrl_addr[8] inst_codemaker/mem_ctrl_addr[9] inst_codemaker/mem_ctrl_in[0]
+ inst_codemaker/mem_ctrl_in[10] inst_codemaker/mem_ctrl_in[11] inst_codemaker/mem_ctrl_in[12]
+ inst_codemaker/mem_ctrl_in[13] inst_codemaker/mem_ctrl_in[14] inst_codemaker/mem_ctrl_in[15]
+ inst_codemaker/mem_ctrl_in[16] inst_codemaker/mem_ctrl_in[17] inst_codemaker/mem_ctrl_in[18]
+ inst_codemaker/mem_ctrl_in[19] inst_codemaker/mem_ctrl_in[1] inst_codemaker/mem_ctrl_in[20]
+ inst_codemaker/mem_ctrl_in[21] inst_codemaker/mem_ctrl_in[22] inst_codemaker/mem_ctrl_in[23]
+ inst_codemaker/mem_ctrl_in[24] inst_codemaker/mem_ctrl_in[25] inst_codemaker/mem_ctrl_in[26]
+ inst_codemaker/mem_ctrl_in[27] inst_codemaker/mem_ctrl_in[28] inst_codemaker/mem_ctrl_in[29]
+ inst_codemaker/mem_ctrl_in[2] inst_codemaker/mem_ctrl_in[30] inst_codemaker/mem_ctrl_in[31]
+ inst_codemaker/mem_ctrl_in[3] inst_codemaker/mem_ctrl_in[4] inst_codemaker/mem_ctrl_in[5]
+ inst_codemaker/mem_ctrl_in[6] inst_codemaker/mem_ctrl_in[7] inst_codemaker/mem_ctrl_in[8]
+ inst_codemaker/mem_ctrl_in[9] inst_codemaker/mem_ctrl_out[0] inst_codemaker/mem_ctrl_out[10]
+ inst_codemaker/mem_ctrl_out[11] inst_codemaker/mem_ctrl_out[12] inst_codemaker/mem_ctrl_out[13]
+ inst_codemaker/mem_ctrl_out[14] inst_codemaker/mem_ctrl_out[15] inst_codemaker/mem_ctrl_out[16]
+ inst_codemaker/mem_ctrl_out[17] inst_codemaker/mem_ctrl_out[18] inst_codemaker/mem_ctrl_out[19]
+ inst_codemaker/mem_ctrl_out[1] inst_codemaker/mem_ctrl_out[20] inst_codemaker/mem_ctrl_out[21]
+ inst_codemaker/mem_ctrl_out[22] inst_codemaker/mem_ctrl_out[23] inst_codemaker/mem_ctrl_out[24]
+ inst_codemaker/mem_ctrl_out[25] inst_codemaker/mem_ctrl_out[26] inst_codemaker/mem_ctrl_out[27]
+ inst_codemaker/mem_ctrl_out[28] inst_codemaker/mem_ctrl_out[29] inst_codemaker/mem_ctrl_out[2]
+ inst_codemaker/mem_ctrl_out[30] inst_codemaker/mem_ctrl_out[31] inst_codemaker/mem_ctrl_out[3]
+ inst_codemaker/mem_ctrl_out[4] inst_codemaker/mem_ctrl_out[5] inst_codemaker/mem_ctrl_out[6]
+ inst_codemaker/mem_ctrl_out[7] inst_codemaker/mem_ctrl_out[8] inst_codemaker/mem_ctrl_out[9]
+ inst_codemaker/mem_ctrl_req inst_codemaker/mem_ctrl_vld inst_codemaker/mem_ctrl_we
+ codemaker_sram2k_inst0/csb0 codemaker_sram2k_inst0/dout0[0] codemaker_sram2k_inst0/dout0[10]
+ codemaker_sram2k_inst0/dout0[11] codemaker_sram2k_inst0/dout0[12] codemaker_sram2k_inst0/dout0[13]
+ codemaker_sram2k_inst0/dout0[14] codemaker_sram2k_inst0/dout0[15] codemaker_sram2k_inst0/dout0[16]
+ codemaker_sram2k_inst0/dout0[17] codemaker_sram2k_inst0/dout0[18] codemaker_sram2k_inst0/dout0[19]
+ codemaker_sram2k_inst0/dout0[1] codemaker_sram2k_inst0/dout0[20] codemaker_sram2k_inst0/dout0[21]
+ codemaker_sram2k_inst0/dout0[22] codemaker_sram2k_inst0/dout0[23] codemaker_sram2k_inst0/dout0[24]
+ codemaker_sram2k_inst0/dout0[25] codemaker_sram2k_inst0/dout0[26] codemaker_sram2k_inst0/dout0[27]
+ codemaker_sram2k_inst0/dout0[28] codemaker_sram2k_inst0/dout0[29] codemaker_sram2k_inst0/dout0[2]
+ codemaker_sram2k_inst0/dout0[30] codemaker_sram2k_inst0/dout0[31] codemaker_sram2k_inst0/dout0[3]
+ codemaker_sram2k_inst0/dout0[4] codemaker_sram2k_inst0/dout0[5] codemaker_sram2k_inst0/dout0[6]
+ codemaker_sram2k_inst0/dout0[7] codemaker_sram2k_inst0/dout0[8] codemaker_sram2k_inst0/dout0[9]
+ codemaker_sram2k_inst0/web0 codemaker_sram2k_inst1/csb0 codemaker_sram2k_inst1/dout0[0]
+ codemaker_sram2k_inst1/dout0[10] codemaker_sram2k_inst1/dout0[11] codemaker_sram2k_inst1/dout0[12]
+ codemaker_sram2k_inst1/dout0[13] codemaker_sram2k_inst1/dout0[14] codemaker_sram2k_inst1/dout0[15]
+ codemaker_sram2k_inst1/dout0[16] codemaker_sram2k_inst1/dout0[17] codemaker_sram2k_inst1/dout0[18]
+ codemaker_sram2k_inst1/dout0[19] codemaker_sram2k_inst1/dout0[1] codemaker_sram2k_inst1/dout0[20]
+ codemaker_sram2k_inst1/dout0[21] codemaker_sram2k_inst1/dout0[22] codemaker_sram2k_inst1/dout0[23]
+ codemaker_sram2k_inst1/dout0[24] codemaker_sram2k_inst1/dout0[25] codemaker_sram2k_inst1/dout0[26]
+ codemaker_sram2k_inst1/dout0[27] codemaker_sram2k_inst1/dout0[28] codemaker_sram2k_inst1/dout0[29]
+ codemaker_sram2k_inst1/dout0[2] codemaker_sram2k_inst1/dout0[30] codemaker_sram2k_inst1/dout0[31]
+ codemaker_sram2k_inst1/dout0[3] codemaker_sram2k_inst1/dout0[4] codemaker_sram2k_inst1/dout0[5]
+ codemaker_sram2k_inst1/dout0[6] codemaker_sram2k_inst1/dout0[7] codemaker_sram2k_inst1/dout0[8]
+ codemaker_sram2k_inst1/dout0[9] codemaker_sram2k_inst1/web0 codemaker_sram2k_inst2/csb0
+ codemaker_sram2k_inst2/dout0[0] codemaker_sram2k_inst2/dout0[10] codemaker_sram2k_inst2/dout0[11]
+ codemaker_sram2k_inst2/dout0[12] codemaker_sram2k_inst2/dout0[13] codemaker_sram2k_inst2/dout0[14]
+ codemaker_sram2k_inst2/dout0[15] codemaker_sram2k_inst2/dout0[16] codemaker_sram2k_inst2/dout0[17]
+ codemaker_sram2k_inst2/dout0[18] codemaker_sram2k_inst2/dout0[19] codemaker_sram2k_inst2/dout0[1]
+ codemaker_sram2k_inst2/dout0[20] codemaker_sram2k_inst2/dout0[21] codemaker_sram2k_inst2/dout0[22]
+ codemaker_sram2k_inst2/dout0[23] codemaker_sram2k_inst2/dout0[24] codemaker_sram2k_inst2/dout0[25]
+ codemaker_sram2k_inst2/dout0[26] codemaker_sram2k_inst2/dout0[27] codemaker_sram2k_inst2/dout0[28]
+ codemaker_sram2k_inst2/dout0[29] codemaker_sram2k_inst2/dout0[2] codemaker_sram2k_inst2/dout0[30]
+ codemaker_sram2k_inst2/dout0[31] codemaker_sram2k_inst2/dout0[3] codemaker_sram2k_inst2/dout0[4]
+ codemaker_sram2k_inst2/dout0[5] codemaker_sram2k_inst2/dout0[6] codemaker_sram2k_inst2/dout0[7]
+ codemaker_sram2k_inst2/dout0[8] codemaker_sram2k_inst2/dout0[9] codemaker_sram2k_inst2/web0
+ codemaker_sram2k_inst3/csb0 codemaker_sram2k_inst3/dout0[0] codemaker_sram2k_inst3/dout0[10]
+ codemaker_sram2k_inst3/dout0[11] codemaker_sram2k_inst3/dout0[12] codemaker_sram2k_inst3/dout0[13]
+ codemaker_sram2k_inst3/dout0[14] codemaker_sram2k_inst3/dout0[15] codemaker_sram2k_inst3/dout0[16]
+ codemaker_sram2k_inst3/dout0[17] codemaker_sram2k_inst3/dout0[18] codemaker_sram2k_inst3/dout0[19]
+ codemaker_sram2k_inst3/dout0[1] codemaker_sram2k_inst3/dout0[20] codemaker_sram2k_inst3/dout0[21]
+ codemaker_sram2k_inst3/dout0[22] codemaker_sram2k_inst3/dout0[23] codemaker_sram2k_inst3/dout0[24]
+ codemaker_sram2k_inst3/dout0[25] codemaker_sram2k_inst3/dout0[26] codemaker_sram2k_inst3/dout0[27]
+ codemaker_sram2k_inst3/dout0[28] codemaker_sram2k_inst3/dout0[29] codemaker_sram2k_inst3/dout0[2]
+ codemaker_sram2k_inst3/dout0[30] codemaker_sram2k_inst3/dout0[31] codemaker_sram2k_inst3/dout0[3]
+ codemaker_sram2k_inst3/dout0[4] codemaker_sram2k_inst3/dout0[5] codemaker_sram2k_inst3/dout0[6]
+ codemaker_sram2k_inst3/dout0[7] codemaker_sram2k_inst3/dout0[8] codemaker_sram2k_inst3/dout0[9]
+ codemaker_sram2k_inst3/web0 codemaker_sram2k_inst3/addr0[0] codemaker_sram2k_inst3/addr0[1]
+ codemaker_sram2k_inst3/addr0[2] codemaker_sram2k_inst3/addr0[3] codemaker_sram2k_inst3/addr0[4]
+ codemaker_sram2k_inst3/addr0[5] codemaker_sram2k_inst3/addr0[6] codemaker_sram2k_inst3/addr0[7]
+ codemaker_sram2k_inst3/addr0[8] codemaker_sram2k_inst3/din0[0] codemaker_sram2k_inst3/din0[10]
+ codemaker_sram2k_inst3/din0[11] codemaker_sram2k_inst3/din0[12] codemaker_sram2k_inst3/din0[13]
+ codemaker_sram2k_inst3/din0[14] codemaker_sram2k_inst3/din0[15] codemaker_sram2k_inst3/din0[16]
+ codemaker_sram2k_inst3/din0[17] codemaker_sram2k_inst3/din0[18] codemaker_sram2k_inst3/din0[19]
+ codemaker_sram2k_inst3/din0[1] codemaker_sram2k_inst3/din0[20] codemaker_sram2k_inst3/din0[21]
+ codemaker_sram2k_inst3/din0[22] codemaker_sram2k_inst3/din0[23] codemaker_sram2k_inst3/din0[24]
+ codemaker_sram2k_inst3/din0[25] codemaker_sram2k_inst3/din0[26] codemaker_sram2k_inst3/din0[27]
+ codemaker_sram2k_inst3/din0[28] codemaker_sram2k_inst3/din0[29] codemaker_sram2k_inst3/din0[2]
+ codemaker_sram2k_inst3/din0[30] codemaker_sram2k_inst3/din0[31] codemaker_sram2k_inst3/din0[3]
+ codemaker_sram2k_inst3/din0[4] codemaker_sram2k_inst3/din0[5] codemaker_sram2k_inst3/din0[6]
+ codemaker_sram2k_inst3/din0[7] codemaker_sram2k_inst3/din0[8] codemaker_sram2k_inst3/din0[9]
+ inst_control_tower/mem_ctrl_addr[0] inst_control_tower/mem_ctrl_addr[10] inst_control_tower/mem_ctrl_addr[11]
+ inst_control_tower/mem_ctrl_addr[12] inst_control_tower/mem_ctrl_addr[13] inst_control_tower/mem_ctrl_addr[1]
+ inst_control_tower/mem_ctrl_addr[2] inst_control_tower/mem_ctrl_addr[3] inst_control_tower/mem_ctrl_addr[4]
+ inst_control_tower/mem_ctrl_addr[5] inst_control_tower/mem_ctrl_addr[6] inst_control_tower/mem_ctrl_addr[7]
+ inst_control_tower/mem_ctrl_addr[8] inst_control_tower/mem_ctrl_addr[9] inst_control_tower/mem_ctrl_in[0]
+ inst_control_tower/mem_ctrl_in[10] inst_control_tower/mem_ctrl_in[11] inst_control_tower/mem_ctrl_in[12]
+ inst_control_tower/mem_ctrl_in[13] inst_control_tower/mem_ctrl_in[14] inst_control_tower/mem_ctrl_in[15]
+ inst_control_tower/mem_ctrl_in[16] inst_control_tower/mem_ctrl_in[17] inst_control_tower/mem_ctrl_in[18]
+ inst_control_tower/mem_ctrl_in[19] inst_control_tower/mem_ctrl_in[1] inst_control_tower/mem_ctrl_in[20]
+ inst_control_tower/mem_ctrl_in[21] inst_control_tower/mem_ctrl_in[22] inst_control_tower/mem_ctrl_in[23]
+ inst_control_tower/mem_ctrl_in[24] inst_control_tower/mem_ctrl_in[25] inst_control_tower/mem_ctrl_in[26]
+ inst_control_tower/mem_ctrl_in[27] inst_control_tower/mem_ctrl_in[28] inst_control_tower/mem_ctrl_in[29]
+ inst_control_tower/mem_ctrl_in[2] inst_control_tower/mem_ctrl_in[30] inst_control_tower/mem_ctrl_in[31]
+ inst_control_tower/mem_ctrl_in[3] inst_control_tower/mem_ctrl_in[4] inst_control_tower/mem_ctrl_in[5]
+ inst_control_tower/mem_ctrl_in[6] inst_control_tower/mem_ctrl_in[7] inst_control_tower/mem_ctrl_in[8]
+ inst_control_tower/mem_ctrl_in[9] inst_control_tower/mem_ctrl_out[0] inst_control_tower/mem_ctrl_out[10]
+ inst_control_tower/mem_ctrl_out[11] inst_control_tower/mem_ctrl_out[12] inst_control_tower/mem_ctrl_out[13]
+ inst_control_tower/mem_ctrl_out[14] inst_control_tower/mem_ctrl_out[15] inst_control_tower/mem_ctrl_out[16]
+ inst_control_tower/mem_ctrl_out[17] inst_control_tower/mem_ctrl_out[18] inst_control_tower/mem_ctrl_out[19]
+ inst_control_tower/mem_ctrl_out[1] inst_control_tower/mem_ctrl_out[20] inst_control_tower/mem_ctrl_out[21]
+ inst_control_tower/mem_ctrl_out[22] inst_control_tower/mem_ctrl_out[23] inst_control_tower/mem_ctrl_out[24]
+ inst_control_tower/mem_ctrl_out[25] inst_control_tower/mem_ctrl_out[26] inst_control_tower/mem_ctrl_out[27]
+ inst_control_tower/mem_ctrl_out[28] inst_control_tower/mem_ctrl_out[29] inst_control_tower/mem_ctrl_out[2]
+ inst_control_tower/mem_ctrl_out[30] inst_control_tower/mem_ctrl_out[31] inst_control_tower/mem_ctrl_out[3]
+ inst_control_tower/mem_ctrl_out[4] inst_control_tower/mem_ctrl_out[5] inst_control_tower/mem_ctrl_out[6]
+ inst_control_tower/mem_ctrl_out[7] inst_control_tower/mem_ctrl_out[8] inst_control_tower/mem_ctrl_out[9]
+ inst_control_tower/mem_ctrl_req inst_control_tower/mem_ctrl_vld inst_control_tower/mem_ctrl_we
+ control_tower_sram2k_inst0/csb0 control_tower_sram2k_inst0/dout0[0] control_tower_sram2k_inst0/dout0[10]
+ control_tower_sram2k_inst0/dout0[11] control_tower_sram2k_inst0/dout0[12] control_tower_sram2k_inst0/dout0[13]
+ control_tower_sram2k_inst0/dout0[14] control_tower_sram2k_inst0/dout0[15] control_tower_sram2k_inst0/dout0[16]
+ control_tower_sram2k_inst0/dout0[17] control_tower_sram2k_inst0/dout0[18] control_tower_sram2k_inst0/dout0[19]
+ control_tower_sram2k_inst0/dout0[1] control_tower_sram2k_inst0/dout0[20] control_tower_sram2k_inst0/dout0[21]
+ control_tower_sram2k_inst0/dout0[22] control_tower_sram2k_inst0/dout0[23] control_tower_sram2k_inst0/dout0[24]
+ control_tower_sram2k_inst0/dout0[25] control_tower_sram2k_inst0/dout0[26] control_tower_sram2k_inst0/dout0[27]
+ control_tower_sram2k_inst0/dout0[28] control_tower_sram2k_inst0/dout0[29] control_tower_sram2k_inst0/dout0[2]
+ control_tower_sram2k_inst0/dout0[30] control_tower_sram2k_inst0/dout0[31] control_tower_sram2k_inst0/dout0[3]
+ control_tower_sram2k_inst0/dout0[4] control_tower_sram2k_inst0/dout0[5] control_tower_sram2k_inst0/dout0[6]
+ control_tower_sram2k_inst0/dout0[7] control_tower_sram2k_inst0/dout0[8] control_tower_sram2k_inst0/dout0[9]
+ control_tower_sram2k_inst0/web0 control_tower_sram2k_inst1/csb0 control_tower_sram2k_inst1/dout0[0]
+ control_tower_sram2k_inst1/dout0[10] control_tower_sram2k_inst1/dout0[11] control_tower_sram2k_inst1/dout0[12]
+ control_tower_sram2k_inst1/dout0[13] control_tower_sram2k_inst1/dout0[14] control_tower_sram2k_inst1/dout0[15]
+ control_tower_sram2k_inst1/dout0[16] control_tower_sram2k_inst1/dout0[17] control_tower_sram2k_inst1/dout0[18]
+ control_tower_sram2k_inst1/dout0[19] control_tower_sram2k_inst1/dout0[1] control_tower_sram2k_inst1/dout0[20]
+ control_tower_sram2k_inst1/dout0[21] control_tower_sram2k_inst1/dout0[22] control_tower_sram2k_inst1/dout0[23]
+ control_tower_sram2k_inst1/dout0[24] control_tower_sram2k_inst1/dout0[25] control_tower_sram2k_inst1/dout0[26]
+ control_tower_sram2k_inst1/dout0[27] control_tower_sram2k_inst1/dout0[28] control_tower_sram2k_inst1/dout0[29]
+ control_tower_sram2k_inst1/dout0[2] control_tower_sram2k_inst1/dout0[30] control_tower_sram2k_inst1/dout0[31]
+ control_tower_sram2k_inst1/dout0[3] control_tower_sram2k_inst1/dout0[4] control_tower_sram2k_inst1/dout0[5]
+ control_tower_sram2k_inst1/dout0[6] control_tower_sram2k_inst1/dout0[7] control_tower_sram2k_inst1/dout0[8]
+ control_tower_sram2k_inst1/dout0[9] control_tower_sram2k_inst1/web0 control_tower_sram2k_inst2/csb0
+ control_tower_sram2k_inst2/dout0[0] control_tower_sram2k_inst2/dout0[10] control_tower_sram2k_inst2/dout0[11]
+ control_tower_sram2k_inst2/dout0[12] control_tower_sram2k_inst2/dout0[13] control_tower_sram2k_inst2/dout0[14]
+ control_tower_sram2k_inst2/dout0[15] control_tower_sram2k_inst2/dout0[16] control_tower_sram2k_inst2/dout0[17]
+ control_tower_sram2k_inst2/dout0[18] control_tower_sram2k_inst2/dout0[19] control_tower_sram2k_inst2/dout0[1]
+ control_tower_sram2k_inst2/dout0[20] control_tower_sram2k_inst2/dout0[21] control_tower_sram2k_inst2/dout0[22]
+ control_tower_sram2k_inst2/dout0[23] control_tower_sram2k_inst2/dout0[24] control_tower_sram2k_inst2/dout0[25]
+ control_tower_sram2k_inst2/dout0[26] control_tower_sram2k_inst2/dout0[27] control_tower_sram2k_inst2/dout0[28]
+ control_tower_sram2k_inst2/dout0[29] control_tower_sram2k_inst2/dout0[2] control_tower_sram2k_inst2/dout0[30]
+ control_tower_sram2k_inst2/dout0[31] control_tower_sram2k_inst2/dout0[3] control_tower_sram2k_inst2/dout0[4]
+ control_tower_sram2k_inst2/dout0[5] control_tower_sram2k_inst2/dout0[6] control_tower_sram2k_inst2/dout0[7]
+ control_tower_sram2k_inst2/dout0[8] control_tower_sram2k_inst2/dout0[9] control_tower_sram2k_inst2/web0
+ control_tower_sram2k_inst3/csb0 control_tower_sram2k_inst3/dout0[0] control_tower_sram2k_inst3/dout0[10]
+ control_tower_sram2k_inst3/dout0[11] control_tower_sram2k_inst3/dout0[12] control_tower_sram2k_inst3/dout0[13]
+ control_tower_sram2k_inst3/dout0[14] control_tower_sram2k_inst3/dout0[15] control_tower_sram2k_inst3/dout0[16]
+ control_tower_sram2k_inst3/dout0[17] control_tower_sram2k_inst3/dout0[18] control_tower_sram2k_inst3/dout0[19]
+ control_tower_sram2k_inst3/dout0[1] control_tower_sram2k_inst3/dout0[20] control_tower_sram2k_inst3/dout0[21]
+ control_tower_sram2k_inst3/dout0[22] control_tower_sram2k_inst3/dout0[23] control_tower_sram2k_inst3/dout0[24]
+ control_tower_sram2k_inst3/dout0[25] control_tower_sram2k_inst3/dout0[26] control_tower_sram2k_inst3/dout0[27]
+ control_tower_sram2k_inst3/dout0[28] control_tower_sram2k_inst3/dout0[29] control_tower_sram2k_inst3/dout0[2]
+ control_tower_sram2k_inst3/dout0[30] control_tower_sram2k_inst3/dout0[31] control_tower_sram2k_inst3/dout0[3]
+ control_tower_sram2k_inst3/dout0[4] control_tower_sram2k_inst3/dout0[5] control_tower_sram2k_inst3/dout0[6]
+ control_tower_sram2k_inst3/dout0[7] control_tower_sram2k_inst3/dout0[8] control_tower_sram2k_inst3/dout0[9]
+ control_tower_sram2k_inst3/web0 control_tower_sram2k_inst4/csb0 control_tower_sram2k_inst4/dout0[0]
+ control_tower_sram2k_inst4/dout0[10] control_tower_sram2k_inst4/dout0[11] control_tower_sram2k_inst4/dout0[12]
+ control_tower_sram2k_inst4/dout0[13] control_tower_sram2k_inst4/dout0[14] control_tower_sram2k_inst4/dout0[15]
+ control_tower_sram2k_inst4/dout0[16] control_tower_sram2k_inst4/dout0[17] control_tower_sram2k_inst4/dout0[18]
+ control_tower_sram2k_inst4/dout0[19] control_tower_sram2k_inst4/dout0[1] control_tower_sram2k_inst4/dout0[20]
+ control_tower_sram2k_inst4/dout0[21] control_tower_sram2k_inst4/dout0[22] control_tower_sram2k_inst4/dout0[23]
+ control_tower_sram2k_inst4/dout0[24] control_tower_sram2k_inst4/dout0[25] control_tower_sram2k_inst4/dout0[26]
+ control_tower_sram2k_inst4/dout0[27] control_tower_sram2k_inst4/dout0[28] control_tower_sram2k_inst4/dout0[29]
+ control_tower_sram2k_inst4/dout0[2] control_tower_sram2k_inst4/dout0[30] control_tower_sram2k_inst4/dout0[31]
+ control_tower_sram2k_inst4/dout0[3] control_tower_sram2k_inst4/dout0[4] control_tower_sram2k_inst4/dout0[5]
+ control_tower_sram2k_inst4/dout0[6] control_tower_sram2k_inst4/dout0[7] control_tower_sram2k_inst4/dout0[8]
+ control_tower_sram2k_inst4/dout0[9] control_tower_sram2k_inst4/web0 control_tower_sram2k_inst4/addr0[0]
+ control_tower_sram2k_inst4/addr0[1] control_tower_sram2k_inst4/addr0[2] control_tower_sram2k_inst4/addr0[3]
+ control_tower_sram2k_inst4/addr0[4] control_tower_sram2k_inst4/addr0[5] control_tower_sram2k_inst4/addr0[6]
+ control_tower_sram2k_inst4/addr0[7] control_tower_sram2k_inst4/addr0[8] control_tower_sram2k_inst4/din0[0]
+ control_tower_sram2k_inst4/din0[10] control_tower_sram2k_inst4/din0[11] control_tower_sram2k_inst4/din0[12]
+ control_tower_sram2k_inst4/din0[13] control_tower_sram2k_inst4/din0[14] control_tower_sram2k_inst4/din0[15]
+ control_tower_sram2k_inst4/din0[16] control_tower_sram2k_inst4/din0[17] control_tower_sram2k_inst4/din0[18]
+ control_tower_sram2k_inst4/din0[19] control_tower_sram2k_inst4/din0[1] control_tower_sram2k_inst4/din0[20]
+ control_tower_sram2k_inst4/din0[21] control_tower_sram2k_inst4/din0[22] control_tower_sram2k_inst4/din0[23]
+ control_tower_sram2k_inst4/din0[24] control_tower_sram2k_inst4/din0[25] control_tower_sram2k_inst4/din0[26]
+ control_tower_sram2k_inst4/din0[27] control_tower_sram2k_inst4/din0[28] control_tower_sram2k_inst4/din0[29]
+ control_tower_sram2k_inst4/din0[2] control_tower_sram2k_inst4/din0[30] control_tower_sram2k_inst4/din0[31]
+ control_tower_sram2k_inst4/din0[3] control_tower_sram2k_inst4/din0[4] control_tower_sram2k_inst4/din0[5]
+ control_tower_sram2k_inst4/din0[6] control_tower_sram2k_inst4/din0[7] control_tower_sram2k_inst4/din0[8]
+ control_tower_sram2k_inst4/din0[9] inst_main_memory/addra[0] inst_main_memory/addra[1]
+ inst_main_memory/addra[2] inst_main_memory/addra[3] inst_main_memory/addra[4] inst_main_memory/addra[5]
+ inst_main_memory/dina[0] inst_main_memory/dina[10] inst_main_memory/dina[11] inst_main_memory/dina[12]
+ inst_main_memory/dina[13] inst_main_memory/dina[14] inst_main_memory/dina[15] inst_main_memory/dina[16]
+ inst_main_memory/dina[17] inst_main_memory/dina[18] inst_main_memory/dina[19] inst_main_memory/dina[1]
+ inst_main_memory/dina[20] inst_main_memory/dina[21] inst_main_memory/dina[22] inst_main_memory/dina[23]
+ inst_main_memory/dina[24] inst_main_memory/dina[25] inst_main_memory/dina[26] inst_main_memory/dina[27]
+ inst_main_memory/dina[28] inst_main_memory/dina[29] inst_main_memory/dina[2] inst_main_memory/dina[30]
+ inst_main_memory/dina[31] inst_main_memory/dina[3] inst_main_memory/dina[4] inst_main_memory/dina[5]
+ inst_main_memory/dina[6] inst_main_memory/dina[7] inst_main_memory/dina[8] inst_main_memory/dina[9]
+ inst_main_memory/douta[0] inst_main_memory/douta[10] inst_main_memory/douta[11]
+ inst_main_memory/douta[12] inst_main_memory/douta[13] inst_main_memory/douta[14]
+ inst_main_memory/douta[15] inst_main_memory/douta[16] inst_main_memory/douta[17]
+ inst_main_memory/douta[18] inst_main_memory/douta[19] inst_main_memory/douta[1]
+ inst_main_memory/douta[20] inst_main_memory/douta[21] inst_main_memory/douta[22]
+ inst_main_memory/douta[23] inst_main_memory/douta[24] inst_main_memory/douta[25]
+ inst_main_memory/douta[26] inst_main_memory/douta[27] inst_main_memory/douta[28]
+ inst_main_memory/douta[29] inst_main_memory/douta[2] inst_main_memory/douta[30]
+ inst_main_memory/douta[31] inst_main_memory/douta[3] inst_main_memory/douta[4] inst_main_memory/douta[5]
+ inst_main_memory/douta[6] inst_main_memory/douta[7] inst_main_memory/douta[8] inst_main_memory/douta[9]
+ inst_main_memory/wea io_in[9] io_in[10] inst_uart/r_data[0] inst_uart/r_data[1]
+ inst_uart/r_data[2] inst_uart/r_data[3] inst_uart/r_data[4] inst_uart/r_data[5]
+ inst_uart/r_data[6] inst_uart/r_data[7] inst_uart/rd_uart io_in[8] inst_uart/reset
+ inst_uart/rx_empty inst_uart/rx_fifo_flush_enable io_oeb[0] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] agent_1_sram2k_inst2/csb1
+ agent_1_sram2k_inst2/wmask0[0] agent_1_sram2k_inst2/wmask0[1] agent_1_sram2k_inst2/wmask0[2]
+ agent_1_sram2k_inst2/wmask0[3] inst_uart/tx_full vccd1 vssd1 inst_uart/w_data[0]
+ inst_uart/w_data[1] inst_uart/w_data[2] inst_uart/w_data[3] inst_uart/w_data[4]
+ inst_uart/w_data[5] inst_uart/w_data[6] inst_uart/w_data[7] inst_uart/wr_uart main_controller
.ends

