magic
tech sky130A
magscale 1 2
timestamp 1655291424
<< obsli1 >>
rect 61104 497159 508852 643817
<< obsm1 >>
rect 566 3408 580506 701004
<< metal2 >>
rect 7626 703520 7738 704960
rect 22990 703520 23102 704960
rect 38354 703520 38466 704960
rect 53718 703520 53830 704960
rect 69082 703520 69194 704960
rect 84446 703520 84558 704960
rect 99810 703520 99922 704960
rect 115174 703520 115286 704960
rect 130538 703520 130650 704960
rect 145902 703520 146014 704960
rect 161266 703520 161378 704960
rect 176630 703520 176742 704960
rect 191994 703520 192106 704960
rect 207358 703520 207470 704960
rect 222722 703520 222834 704960
rect 238086 703520 238198 704960
rect 253450 703520 253562 704960
rect 268814 703520 268926 704960
rect 284178 703520 284290 704960
rect 299634 703520 299746 704960
rect 314998 703520 315110 704960
rect 330362 703520 330474 704960
rect 345726 703520 345838 704960
rect 361090 703520 361202 704960
rect 376454 703520 376566 704960
rect 391818 703520 391930 704960
rect 407182 703520 407294 704960
rect 422546 703520 422658 704960
rect 437910 703520 438022 704960
rect 453274 703520 453386 704960
rect 468638 703520 468750 704960
rect 484002 703520 484114 704960
rect 499366 703520 499478 704960
rect 514730 703520 514842 704960
rect 530094 703520 530206 704960
rect 545458 703520 545570 704960
rect 560822 703520 560934 704960
rect 576186 703520 576298 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6338 -960 6450 480
rect 7534 -960 7646 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12226 -960 12338 480
rect 13422 -960 13534 480
rect 14618 -960 14730 480
rect 15814 -960 15926 480
rect 17010 -960 17122 480
rect 18114 -960 18226 480
rect 19310 -960 19422 480
rect 20506 -960 20618 480
rect 21702 -960 21814 480
rect 22898 -960 23010 480
rect 24002 -960 24114 480
rect 25198 -960 25310 480
rect 26394 -960 26506 480
rect 27590 -960 27702 480
rect 28786 -960 28898 480
rect 29890 -960 30002 480
rect 31086 -960 31198 480
rect 32282 -960 32394 480
rect 33478 -960 33590 480
rect 34674 -960 34786 480
rect 35778 -960 35890 480
rect 36974 -960 37086 480
rect 38170 -960 38282 480
rect 39366 -960 39478 480
rect 40562 -960 40674 480
rect 41666 -960 41778 480
rect 42862 -960 42974 480
rect 44058 -960 44170 480
rect 45254 -960 45366 480
rect 46450 -960 46562 480
rect 47554 -960 47666 480
rect 48750 -960 48862 480
rect 49946 -960 50058 480
rect 51142 -960 51254 480
rect 52338 -960 52450 480
rect 53442 -960 53554 480
rect 54638 -960 54750 480
rect 55834 -960 55946 480
rect 57030 -960 57142 480
rect 58226 -960 58338 480
rect 59330 -960 59442 480
rect 60526 -960 60638 480
rect 61722 -960 61834 480
rect 62918 -960 63030 480
rect 64114 -960 64226 480
rect 65218 -960 65330 480
rect 66414 -960 66526 480
rect 67610 -960 67722 480
rect 68806 -960 68918 480
rect 70002 -960 70114 480
rect 71106 -960 71218 480
rect 72302 -960 72414 480
rect 73498 -960 73610 480
rect 74694 -960 74806 480
rect 75890 -960 76002 480
rect 76994 -960 77106 480
rect 78190 -960 78302 480
rect 79386 -960 79498 480
rect 80582 -960 80694 480
rect 81778 -960 81890 480
rect 82882 -960 82994 480
rect 84078 -960 84190 480
rect 85274 -960 85386 480
rect 86470 -960 86582 480
rect 87666 -960 87778 480
rect 88770 -960 88882 480
rect 89966 -960 90078 480
rect 91162 -960 91274 480
rect 92358 -960 92470 480
rect 93554 -960 93666 480
rect 94658 -960 94770 480
rect 95854 -960 95966 480
rect 97050 -960 97162 480
rect 98246 -960 98358 480
rect 99442 -960 99554 480
rect 100546 -960 100658 480
rect 101742 -960 101854 480
rect 102938 -960 103050 480
rect 104134 -960 104246 480
rect 105330 -960 105442 480
rect 106434 -960 106546 480
rect 107630 -960 107742 480
rect 108826 -960 108938 480
rect 110022 -960 110134 480
rect 111218 -960 111330 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124098 -960 124210 480
rect 125294 -960 125406 480
rect 126490 -960 126602 480
rect 127686 -960 127798 480
rect 128882 -960 128994 480
rect 129986 -960 130098 480
rect 131182 -960 131294 480
rect 132378 -960 132490 480
rect 133574 -960 133686 480
rect 134770 -960 134882 480
rect 135874 -960 135986 480
rect 137070 -960 137182 480
rect 138266 -960 138378 480
rect 139462 -960 139574 480
rect 140658 -960 140770 480
rect 141762 -960 141874 480
rect 142958 -960 143070 480
rect 144154 -960 144266 480
rect 145350 -960 145462 480
rect 146546 -960 146658 480
rect 147650 -960 147762 480
rect 148846 -960 148958 480
rect 150042 -960 150154 480
rect 151238 -960 151350 480
rect 152342 -960 152454 480
rect 153538 -960 153650 480
rect 154734 -960 154846 480
rect 155930 -960 156042 480
rect 157126 -960 157238 480
rect 158230 -960 158342 480
rect 159426 -960 159538 480
rect 160622 -960 160734 480
rect 161818 -960 161930 480
rect 163014 -960 163126 480
rect 164118 -960 164230 480
rect 165314 -960 165426 480
rect 166510 -960 166622 480
rect 167706 -960 167818 480
rect 168902 -960 169014 480
rect 170006 -960 170118 480
rect 171202 -960 171314 480
rect 172398 -960 172510 480
rect 173594 -960 173706 480
rect 174790 -960 174902 480
rect 175894 -960 176006 480
rect 177090 -960 177202 480
rect 178286 -960 178398 480
rect 179482 -960 179594 480
rect 180678 -960 180790 480
rect 181782 -960 181894 480
rect 182978 -960 183090 480
rect 184174 -960 184286 480
rect 185370 -960 185482 480
rect 186566 -960 186678 480
rect 187670 -960 187782 480
rect 188866 -960 188978 480
rect 190062 -960 190174 480
rect 191258 -960 191370 480
rect 192454 -960 192566 480
rect 193558 -960 193670 480
rect 194754 -960 194866 480
rect 195950 -960 196062 480
rect 197146 -960 197258 480
rect 198342 -960 198454 480
rect 199446 -960 199558 480
rect 200642 -960 200754 480
rect 201838 -960 201950 480
rect 203034 -960 203146 480
rect 204230 -960 204342 480
rect 205334 -960 205446 480
rect 206530 -960 206642 480
rect 207726 -960 207838 480
rect 208922 -960 209034 480
rect 210118 -960 210230 480
rect 211222 -960 211334 480
rect 212418 -960 212530 480
rect 213614 -960 213726 480
rect 214810 -960 214922 480
rect 216006 -960 216118 480
rect 217110 -960 217222 480
rect 218306 -960 218418 480
rect 219502 -960 219614 480
rect 220698 -960 220810 480
rect 221894 -960 222006 480
rect 222998 -960 223110 480
rect 224194 -960 224306 480
rect 225390 -960 225502 480
rect 226586 -960 226698 480
rect 227782 -960 227894 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240662 -960 240774 480
rect 241858 -960 241970 480
rect 243054 -960 243166 480
rect 244250 -960 244362 480
rect 245446 -960 245558 480
rect 246550 -960 246662 480
rect 247746 -960 247858 480
rect 248942 -960 249054 480
rect 250138 -960 250250 480
rect 251334 -960 251446 480
rect 252438 -960 252550 480
rect 253634 -960 253746 480
rect 254830 -960 254942 480
rect 256026 -960 256138 480
rect 257222 -960 257334 480
rect 258326 -960 258438 480
rect 259522 -960 259634 480
rect 260718 -960 260830 480
rect 261914 -960 262026 480
rect 263110 -960 263222 480
rect 264214 -960 264326 480
rect 265410 -960 265522 480
rect 266606 -960 266718 480
rect 267802 -960 267914 480
rect 268998 -960 269110 480
rect 270102 -960 270214 480
rect 271298 -960 271410 480
rect 272494 -960 272606 480
rect 273690 -960 273802 480
rect 274886 -960 274998 480
rect 275990 -960 276102 480
rect 277186 -960 277298 480
rect 278382 -960 278494 480
rect 279578 -960 279690 480
rect 280774 -960 280886 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285466 -960 285578 480
rect 286662 -960 286774 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298346 -960 298458 480
rect 299542 -960 299654 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304234 -960 304346 480
rect 305430 -960 305542 480
rect 306626 -960 306738 480
rect 307822 -960 307934 480
rect 309018 -960 309130 480
rect 310122 -960 310234 480
rect 311318 -960 311430 480
rect 312514 -960 312626 480
rect 313710 -960 313822 480
rect 314906 -960 315018 480
rect 316010 -960 316122 480
rect 317206 -960 317318 480
rect 318402 -960 318514 480
rect 319598 -960 319710 480
rect 320794 -960 320906 480
rect 321898 -960 322010 480
rect 323094 -960 323206 480
rect 324290 -960 324402 480
rect 325486 -960 325598 480
rect 326682 -960 326794 480
rect 327786 -960 327898 480
rect 328982 -960 329094 480
rect 330178 -960 330290 480
rect 331374 -960 331486 480
rect 332570 -960 332682 480
rect 333674 -960 333786 480
rect 334870 -960 334982 480
rect 336066 -960 336178 480
rect 337262 -960 337374 480
rect 338458 -960 338570 480
rect 339562 -960 339674 480
rect 340758 -960 340870 480
rect 341954 -960 342066 480
rect 343150 -960 343262 480
rect 344346 -960 344458 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357226 -960 357338 480
rect 358422 -960 358534 480
rect 359618 -960 359730 480
rect 360814 -960 360926 480
rect 362010 -960 362122 480
rect 363114 -960 363226 480
rect 364310 -960 364422 480
rect 365506 -960 365618 480
rect 366702 -960 366814 480
rect 367898 -960 368010 480
rect 369002 -960 369114 480
rect 370198 -960 370310 480
rect 371394 -960 371506 480
rect 372590 -960 372702 480
rect 373786 -960 373898 480
rect 374890 -960 375002 480
rect 376086 -960 376198 480
rect 377282 -960 377394 480
rect 378478 -960 378590 480
rect 379674 -960 379786 480
rect 380778 -960 380890 480
rect 381974 -960 382086 480
rect 383170 -960 383282 480
rect 384366 -960 384478 480
rect 385562 -960 385674 480
rect 386666 -960 386778 480
rect 387862 -960 387974 480
rect 389058 -960 389170 480
rect 390254 -960 390366 480
rect 391450 -960 391562 480
rect 392554 -960 392666 480
rect 393750 -960 393862 480
rect 394946 -960 395058 480
rect 396142 -960 396254 480
rect 397338 -960 397450 480
rect 398442 -960 398554 480
rect 399638 -960 399750 480
rect 400834 -960 400946 480
rect 402030 -960 402142 480
rect 403226 -960 403338 480
rect 404330 -960 404442 480
rect 405526 -960 405638 480
rect 406722 -960 406834 480
rect 407918 -960 408030 480
rect 409114 -960 409226 480
rect 410218 -960 410330 480
rect 411414 -960 411526 480
rect 412610 -960 412722 480
rect 413806 -960 413918 480
rect 415002 -960 415114 480
rect 416106 -960 416218 480
rect 417302 -960 417414 480
rect 418498 -960 418610 480
rect 419694 -960 419806 480
rect 420890 -960 421002 480
rect 421994 -960 422106 480
rect 423190 -960 423302 480
rect 424386 -960 424498 480
rect 425582 -960 425694 480
rect 426778 -960 426890 480
rect 427882 -960 427994 480
rect 429078 -960 429190 480
rect 430274 -960 430386 480
rect 431470 -960 431582 480
rect 432666 -960 432778 480
rect 433770 -960 433882 480
rect 434966 -960 435078 480
rect 436162 -960 436274 480
rect 437358 -960 437470 480
rect 438554 -960 438666 480
rect 439658 -960 439770 480
rect 440854 -960 440966 480
rect 442050 -960 442162 480
rect 443246 -960 443358 480
rect 444350 -960 444462 480
rect 445546 -960 445658 480
rect 446742 -960 446854 480
rect 447938 -960 448050 480
rect 449134 -960 449246 480
rect 450238 -960 450350 480
rect 451434 -960 451546 480
rect 452630 -960 452742 480
rect 453826 -960 453938 480
rect 455022 -960 455134 480
rect 456126 -960 456238 480
rect 457322 -960 457434 480
rect 458518 -960 458630 480
rect 459714 -960 459826 480
rect 460910 -960 461022 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473790 -960 473902 480
rect 474986 -960 475098 480
rect 476182 -960 476294 480
rect 477378 -960 477490 480
rect 478574 -960 478686 480
rect 479678 -960 479790 480
rect 480874 -960 480986 480
rect 482070 -960 482182 480
rect 483266 -960 483378 480
rect 484462 -960 484574 480
rect 485566 -960 485678 480
rect 486762 -960 486874 480
rect 487958 -960 488070 480
rect 489154 -960 489266 480
rect 490350 -960 490462 480
rect 491454 -960 491566 480
rect 492650 -960 492762 480
rect 493846 -960 493958 480
rect 495042 -960 495154 480
rect 496238 -960 496350 480
rect 497342 -960 497454 480
rect 498538 -960 498650 480
rect 499734 -960 499846 480
rect 500930 -960 501042 480
rect 502126 -960 502238 480
rect 503230 -960 503342 480
rect 504426 -960 504538 480
rect 505622 -960 505734 480
rect 506818 -960 506930 480
rect 508014 -960 508126 480
rect 509118 -960 509230 480
rect 510314 -960 510426 480
rect 511510 -960 511622 480
rect 512706 -960 512818 480
rect 513902 -960 514014 480
rect 515006 -960 515118 480
rect 516202 -960 516314 480
rect 517398 -960 517510 480
rect 518594 -960 518706 480
rect 519790 -960 519902 480
rect 520894 -960 521006 480
rect 522090 -960 522202 480
rect 523286 -960 523398 480
rect 524482 -960 524594 480
rect 525678 -960 525790 480
rect 526782 -960 526894 480
rect 527978 -960 528090 480
rect 529174 -960 529286 480
rect 530370 -960 530482 480
rect 531566 -960 531678 480
rect 532670 -960 532782 480
rect 533866 -960 533978 480
rect 535062 -960 535174 480
rect 536258 -960 536370 480
rect 537454 -960 537566 480
rect 538558 -960 538670 480
rect 539754 -960 539866 480
rect 540950 -960 541062 480
rect 542146 -960 542258 480
rect 543342 -960 543454 480
rect 544446 -960 544558 480
rect 545642 -960 545754 480
rect 546838 -960 546950 480
rect 548034 -960 548146 480
rect 549230 -960 549342 480
rect 550334 -960 550446 480
rect 551530 -960 551642 480
rect 552726 -960 552838 480
rect 553922 -960 554034 480
rect 555118 -960 555230 480
rect 556222 -960 556334 480
rect 557418 -960 557530 480
rect 558614 -960 558726 480
rect 559810 -960 559922 480
rect 561006 -960 561118 480
rect 562110 -960 562222 480
rect 563306 -960 563418 480
rect 564502 -960 564614 480
rect 565698 -960 565810 480
rect 566894 -960 567006 480
rect 567998 -960 568110 480
rect 569194 -960 569306 480
rect 570390 -960 570502 480
rect 571586 -960 571698 480
rect 572782 -960 572894 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577474 -960 577586 480
rect 578670 -960 578782 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 7570 703610
rect 7794 703464 22934 703610
rect 23158 703464 38298 703610
rect 38522 703464 53662 703610
rect 53886 703464 69026 703610
rect 69250 703464 84390 703610
rect 84614 703464 99754 703610
rect 99978 703464 115118 703610
rect 115342 703464 130482 703610
rect 130706 703464 145846 703610
rect 146070 703464 161210 703610
rect 161434 703464 176574 703610
rect 176798 703464 191938 703610
rect 192162 703464 207302 703610
rect 207526 703464 222666 703610
rect 222890 703464 238030 703610
rect 238254 703464 253394 703610
rect 253618 703464 268758 703610
rect 268982 703464 284122 703610
rect 284346 703464 299578 703610
rect 299802 703464 314942 703610
rect 315166 703464 330306 703610
rect 330530 703464 345670 703610
rect 345894 703464 361034 703610
rect 361258 703464 376398 703610
rect 376622 703464 391762 703610
rect 391986 703464 407126 703610
rect 407350 703464 422490 703610
rect 422714 703464 437854 703610
rect 438078 703464 453218 703610
rect 453442 703464 468582 703610
rect 468806 703464 483946 703610
rect 484170 703464 499310 703610
rect 499534 703464 514674 703610
rect 514898 703464 530038 703610
rect 530262 703464 545402 703610
rect 545626 703464 560766 703610
rect 560990 703464 576130 703610
rect 576354 703464 580962 703610
rect 572 536 580962 703464
rect 710 480 1590 536
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6282 536
rect 6506 480 7478 536
rect 7702 480 8674 536
rect 8898 480 9870 536
rect 10094 480 11066 536
rect 11290 480 12170 536
rect 12394 480 13366 536
rect 13590 480 14562 536
rect 14786 480 15758 536
rect 15982 480 16954 536
rect 17178 480 18058 536
rect 18282 480 19254 536
rect 19478 480 20450 536
rect 20674 480 21646 536
rect 21870 480 22842 536
rect 23066 480 23946 536
rect 24170 480 25142 536
rect 25366 480 26338 536
rect 26562 480 27534 536
rect 27758 480 28730 536
rect 28954 480 29834 536
rect 30058 480 31030 536
rect 31254 480 32226 536
rect 32450 480 33422 536
rect 33646 480 34618 536
rect 34842 480 35722 536
rect 35946 480 36918 536
rect 37142 480 38114 536
rect 38338 480 39310 536
rect 39534 480 40506 536
rect 40730 480 41610 536
rect 41834 480 42806 536
rect 43030 480 44002 536
rect 44226 480 45198 536
rect 45422 480 46394 536
rect 46618 480 47498 536
rect 47722 480 48694 536
rect 48918 480 49890 536
rect 50114 480 51086 536
rect 51310 480 52282 536
rect 52506 480 53386 536
rect 53610 480 54582 536
rect 54806 480 55778 536
rect 56002 480 56974 536
rect 57198 480 58170 536
rect 58394 480 59274 536
rect 59498 480 60470 536
rect 60694 480 61666 536
rect 61890 480 62862 536
rect 63086 480 64058 536
rect 64282 480 65162 536
rect 65386 480 66358 536
rect 66582 480 67554 536
rect 67778 480 68750 536
rect 68974 480 69946 536
rect 70170 480 71050 536
rect 71274 480 72246 536
rect 72470 480 73442 536
rect 73666 480 74638 536
rect 74862 480 75834 536
rect 76058 480 76938 536
rect 77162 480 78134 536
rect 78358 480 79330 536
rect 79554 480 80526 536
rect 80750 480 81722 536
rect 81946 480 82826 536
rect 83050 480 84022 536
rect 84246 480 85218 536
rect 85442 480 86414 536
rect 86638 480 87610 536
rect 87834 480 88714 536
rect 88938 480 89910 536
rect 90134 480 91106 536
rect 91330 480 92302 536
rect 92526 480 93498 536
rect 93722 480 94602 536
rect 94826 480 95798 536
rect 96022 480 96994 536
rect 97218 480 98190 536
rect 98414 480 99386 536
rect 99610 480 100490 536
rect 100714 480 101686 536
rect 101910 480 102882 536
rect 103106 480 104078 536
rect 104302 480 105274 536
rect 105498 480 106378 536
rect 106602 480 107574 536
rect 107798 480 108770 536
rect 108994 480 109966 536
rect 110190 480 111162 536
rect 111386 480 112266 536
rect 112490 480 113462 536
rect 113686 480 114658 536
rect 114882 480 115854 536
rect 116078 480 117050 536
rect 117274 480 118154 536
rect 118378 480 119350 536
rect 119574 480 120546 536
rect 120770 480 121742 536
rect 121966 480 122938 536
rect 123162 480 124042 536
rect 124266 480 125238 536
rect 125462 480 126434 536
rect 126658 480 127630 536
rect 127854 480 128826 536
rect 129050 480 129930 536
rect 130154 480 131126 536
rect 131350 480 132322 536
rect 132546 480 133518 536
rect 133742 480 134714 536
rect 134938 480 135818 536
rect 136042 480 137014 536
rect 137238 480 138210 536
rect 138434 480 139406 536
rect 139630 480 140602 536
rect 140826 480 141706 536
rect 141930 480 142902 536
rect 143126 480 144098 536
rect 144322 480 145294 536
rect 145518 480 146490 536
rect 146714 480 147594 536
rect 147818 480 148790 536
rect 149014 480 149986 536
rect 150210 480 151182 536
rect 151406 480 152286 536
rect 152510 480 153482 536
rect 153706 480 154678 536
rect 154902 480 155874 536
rect 156098 480 157070 536
rect 157294 480 158174 536
rect 158398 480 159370 536
rect 159594 480 160566 536
rect 160790 480 161762 536
rect 161986 480 162958 536
rect 163182 480 164062 536
rect 164286 480 165258 536
rect 165482 480 166454 536
rect 166678 480 167650 536
rect 167874 480 168846 536
rect 169070 480 169950 536
rect 170174 480 171146 536
rect 171370 480 172342 536
rect 172566 480 173538 536
rect 173762 480 174734 536
rect 174958 480 175838 536
rect 176062 480 177034 536
rect 177258 480 178230 536
rect 178454 480 179426 536
rect 179650 480 180622 536
rect 180846 480 181726 536
rect 181950 480 182922 536
rect 183146 480 184118 536
rect 184342 480 185314 536
rect 185538 480 186510 536
rect 186734 480 187614 536
rect 187838 480 188810 536
rect 189034 480 190006 536
rect 190230 480 191202 536
rect 191426 480 192398 536
rect 192622 480 193502 536
rect 193726 480 194698 536
rect 194922 480 195894 536
rect 196118 480 197090 536
rect 197314 480 198286 536
rect 198510 480 199390 536
rect 199614 480 200586 536
rect 200810 480 201782 536
rect 202006 480 202978 536
rect 203202 480 204174 536
rect 204398 480 205278 536
rect 205502 480 206474 536
rect 206698 480 207670 536
rect 207894 480 208866 536
rect 209090 480 210062 536
rect 210286 480 211166 536
rect 211390 480 212362 536
rect 212586 480 213558 536
rect 213782 480 214754 536
rect 214978 480 215950 536
rect 216174 480 217054 536
rect 217278 480 218250 536
rect 218474 480 219446 536
rect 219670 480 220642 536
rect 220866 480 221838 536
rect 222062 480 222942 536
rect 223166 480 224138 536
rect 224362 480 225334 536
rect 225558 480 226530 536
rect 226754 480 227726 536
rect 227950 480 228830 536
rect 229054 480 230026 536
rect 230250 480 231222 536
rect 231446 480 232418 536
rect 232642 480 233614 536
rect 233838 480 234718 536
rect 234942 480 235914 536
rect 236138 480 237110 536
rect 237334 480 238306 536
rect 238530 480 239502 536
rect 239726 480 240606 536
rect 240830 480 241802 536
rect 242026 480 242998 536
rect 243222 480 244194 536
rect 244418 480 245390 536
rect 245614 480 246494 536
rect 246718 480 247690 536
rect 247914 480 248886 536
rect 249110 480 250082 536
rect 250306 480 251278 536
rect 251502 480 252382 536
rect 252606 480 253578 536
rect 253802 480 254774 536
rect 254998 480 255970 536
rect 256194 480 257166 536
rect 257390 480 258270 536
rect 258494 480 259466 536
rect 259690 480 260662 536
rect 260886 480 261858 536
rect 262082 480 263054 536
rect 263278 480 264158 536
rect 264382 480 265354 536
rect 265578 480 266550 536
rect 266774 480 267746 536
rect 267970 480 268942 536
rect 269166 480 270046 536
rect 270270 480 271242 536
rect 271466 480 272438 536
rect 272662 480 273634 536
rect 273858 480 274830 536
rect 275054 480 275934 536
rect 276158 480 277130 536
rect 277354 480 278326 536
rect 278550 480 279522 536
rect 279746 480 280718 536
rect 280942 480 281822 536
rect 282046 480 283018 536
rect 283242 480 284214 536
rect 284438 480 285410 536
rect 285634 480 286606 536
rect 286830 480 287710 536
rect 287934 480 288906 536
rect 289130 480 290102 536
rect 290326 480 291298 536
rect 291522 480 292494 536
rect 292718 480 293598 536
rect 293822 480 294794 536
rect 295018 480 295990 536
rect 296214 480 297186 536
rect 297410 480 298290 536
rect 298514 480 299486 536
rect 299710 480 300682 536
rect 300906 480 301878 536
rect 302102 480 303074 536
rect 303298 480 304178 536
rect 304402 480 305374 536
rect 305598 480 306570 536
rect 306794 480 307766 536
rect 307990 480 308962 536
rect 309186 480 310066 536
rect 310290 480 311262 536
rect 311486 480 312458 536
rect 312682 480 313654 536
rect 313878 480 314850 536
rect 315074 480 315954 536
rect 316178 480 317150 536
rect 317374 480 318346 536
rect 318570 480 319542 536
rect 319766 480 320738 536
rect 320962 480 321842 536
rect 322066 480 323038 536
rect 323262 480 324234 536
rect 324458 480 325430 536
rect 325654 480 326626 536
rect 326850 480 327730 536
rect 327954 480 328926 536
rect 329150 480 330122 536
rect 330346 480 331318 536
rect 331542 480 332514 536
rect 332738 480 333618 536
rect 333842 480 334814 536
rect 335038 480 336010 536
rect 336234 480 337206 536
rect 337430 480 338402 536
rect 338626 480 339506 536
rect 339730 480 340702 536
rect 340926 480 341898 536
rect 342122 480 343094 536
rect 343318 480 344290 536
rect 344514 480 345394 536
rect 345618 480 346590 536
rect 346814 480 347786 536
rect 348010 480 348982 536
rect 349206 480 350178 536
rect 350402 480 351282 536
rect 351506 480 352478 536
rect 352702 480 353674 536
rect 353898 480 354870 536
rect 355094 480 356066 536
rect 356290 480 357170 536
rect 357394 480 358366 536
rect 358590 480 359562 536
rect 359786 480 360758 536
rect 360982 480 361954 536
rect 362178 480 363058 536
rect 363282 480 364254 536
rect 364478 480 365450 536
rect 365674 480 366646 536
rect 366870 480 367842 536
rect 368066 480 368946 536
rect 369170 480 370142 536
rect 370366 480 371338 536
rect 371562 480 372534 536
rect 372758 480 373730 536
rect 373954 480 374834 536
rect 375058 480 376030 536
rect 376254 480 377226 536
rect 377450 480 378422 536
rect 378646 480 379618 536
rect 379842 480 380722 536
rect 380946 480 381918 536
rect 382142 480 383114 536
rect 383338 480 384310 536
rect 384534 480 385506 536
rect 385730 480 386610 536
rect 386834 480 387806 536
rect 388030 480 389002 536
rect 389226 480 390198 536
rect 390422 480 391394 536
rect 391618 480 392498 536
rect 392722 480 393694 536
rect 393918 480 394890 536
rect 395114 480 396086 536
rect 396310 480 397282 536
rect 397506 480 398386 536
rect 398610 480 399582 536
rect 399806 480 400778 536
rect 401002 480 401974 536
rect 402198 480 403170 536
rect 403394 480 404274 536
rect 404498 480 405470 536
rect 405694 480 406666 536
rect 406890 480 407862 536
rect 408086 480 409058 536
rect 409282 480 410162 536
rect 410386 480 411358 536
rect 411582 480 412554 536
rect 412778 480 413750 536
rect 413974 480 414946 536
rect 415170 480 416050 536
rect 416274 480 417246 536
rect 417470 480 418442 536
rect 418666 480 419638 536
rect 419862 480 420834 536
rect 421058 480 421938 536
rect 422162 480 423134 536
rect 423358 480 424330 536
rect 424554 480 425526 536
rect 425750 480 426722 536
rect 426946 480 427826 536
rect 428050 480 429022 536
rect 429246 480 430218 536
rect 430442 480 431414 536
rect 431638 480 432610 536
rect 432834 480 433714 536
rect 433938 480 434910 536
rect 435134 480 436106 536
rect 436330 480 437302 536
rect 437526 480 438498 536
rect 438722 480 439602 536
rect 439826 480 440798 536
rect 441022 480 441994 536
rect 442218 480 443190 536
rect 443414 480 444294 536
rect 444518 480 445490 536
rect 445714 480 446686 536
rect 446910 480 447882 536
rect 448106 480 449078 536
rect 449302 480 450182 536
rect 450406 480 451378 536
rect 451602 480 452574 536
rect 452798 480 453770 536
rect 453994 480 454966 536
rect 455190 480 456070 536
rect 456294 480 457266 536
rect 457490 480 458462 536
rect 458686 480 459658 536
rect 459882 480 460854 536
rect 461078 480 461958 536
rect 462182 480 463154 536
rect 463378 480 464350 536
rect 464574 480 465546 536
rect 465770 480 466742 536
rect 466966 480 467846 536
rect 468070 480 469042 536
rect 469266 480 470238 536
rect 470462 480 471434 536
rect 471658 480 472630 536
rect 472854 480 473734 536
rect 473958 480 474930 536
rect 475154 480 476126 536
rect 476350 480 477322 536
rect 477546 480 478518 536
rect 478742 480 479622 536
rect 479846 480 480818 536
rect 481042 480 482014 536
rect 482238 480 483210 536
rect 483434 480 484406 536
rect 484630 480 485510 536
rect 485734 480 486706 536
rect 486930 480 487902 536
rect 488126 480 489098 536
rect 489322 480 490294 536
rect 490518 480 491398 536
rect 491622 480 492594 536
rect 492818 480 493790 536
rect 494014 480 494986 536
rect 495210 480 496182 536
rect 496406 480 497286 536
rect 497510 480 498482 536
rect 498706 480 499678 536
rect 499902 480 500874 536
rect 501098 480 502070 536
rect 502294 480 503174 536
rect 503398 480 504370 536
rect 504594 480 505566 536
rect 505790 480 506762 536
rect 506986 480 507958 536
rect 508182 480 509062 536
rect 509286 480 510258 536
rect 510482 480 511454 536
rect 511678 480 512650 536
rect 512874 480 513846 536
rect 514070 480 514950 536
rect 515174 480 516146 536
rect 516370 480 517342 536
rect 517566 480 518538 536
rect 518762 480 519734 536
rect 519958 480 520838 536
rect 521062 480 522034 536
rect 522258 480 523230 536
rect 523454 480 524426 536
rect 524650 480 525622 536
rect 525846 480 526726 536
rect 526950 480 527922 536
rect 528146 480 529118 536
rect 529342 480 530314 536
rect 530538 480 531510 536
rect 531734 480 532614 536
rect 532838 480 533810 536
rect 534034 480 535006 536
rect 535230 480 536202 536
rect 536426 480 537398 536
rect 537622 480 538502 536
rect 538726 480 539698 536
rect 539922 480 540894 536
rect 541118 480 542090 536
rect 542314 480 543286 536
rect 543510 480 544390 536
rect 544614 480 545586 536
rect 545810 480 546782 536
rect 547006 480 547978 536
rect 548202 480 549174 536
rect 549398 480 550278 536
rect 550502 480 551474 536
rect 551698 480 552670 536
rect 552894 480 553866 536
rect 554090 480 555062 536
rect 555286 480 556166 536
rect 556390 480 557362 536
rect 557586 480 558558 536
rect 558782 480 559754 536
rect 559978 480 560950 536
rect 561174 480 562054 536
rect 562278 480 563250 536
rect 563474 480 564446 536
rect 564670 480 565642 536
rect 565866 480 566838 536
rect 567062 480 567942 536
rect 568166 480 569138 536
rect 569362 480 570334 536
rect 570558 480 571530 536
rect 571754 480 572726 536
rect 572950 480 573830 536
rect 574054 480 575026 536
rect 575250 480 576222 536
rect 576446 480 577418 536
rect 577642 480 578614 536
rect 578838 480 579718 536
rect 579942 480 580914 536
<< metal3 >>
rect -960 697492 480 697732
rect 583520 697356 584960 697596
rect -960 684980 480 685220
rect 583520 684572 584960 684812
rect -960 672332 480 672572
rect 583520 671788 584960 672028
rect -960 659820 480 660060
rect 583520 659004 584960 659244
rect -960 647172 480 647412
rect 583520 646220 584960 646460
rect -960 634660 480 634900
rect 583520 633436 584960 633676
rect -960 622148 480 622388
rect 583520 620652 584960 620892
rect -960 609500 480 609740
rect 583520 607868 584960 608108
rect -960 596988 480 597228
rect 583520 595084 584960 595324
rect -960 584340 480 584580
rect 583520 582164 584960 582404
rect -960 571828 480 572068
rect 583520 569380 584960 569620
rect -960 559180 480 559420
rect 583520 556596 584960 556836
rect -960 546668 480 546908
rect 583520 543812 584960 544052
rect -960 534156 480 534396
rect 583520 531028 584960 531268
rect -960 521508 480 521748
rect 583520 518244 584960 518484
rect -960 508996 480 509236
rect 583520 505460 584960 505700
rect -960 496348 480 496588
rect 583520 492676 584960 492916
rect -960 483836 480 484076
rect 583520 479892 584960 480132
rect -960 471188 480 471428
rect 583520 466972 584960 467212
rect -960 458676 480 458916
rect 583520 454188 584960 454428
rect -960 446164 480 446404
rect 583520 441404 584960 441644
rect -960 433516 480 433756
rect 583520 428620 584960 428860
rect -960 421004 480 421244
rect 583520 415836 584960 416076
rect -960 408356 480 408596
rect 583520 403052 584960 403292
rect -960 395844 480 396084
rect 583520 390268 584960 390508
rect -960 383196 480 383436
rect 583520 377484 584960 377724
rect -960 370684 480 370924
rect 583520 364700 584960 364940
rect -960 358172 480 358412
rect 583520 351780 584960 352020
rect -960 345524 480 345764
rect 583520 338996 584960 339236
rect -960 333012 480 333252
rect 583520 326212 584960 326452
rect -960 320364 480 320604
rect 583520 313428 584960 313668
rect -960 307852 480 308092
rect 583520 300644 584960 300884
rect -960 295204 480 295444
rect 583520 287860 584960 288100
rect -960 282692 480 282932
rect 583520 275076 584960 275316
rect -960 270180 480 270420
rect 583520 262292 584960 262532
rect -960 257532 480 257772
rect 583520 249508 584960 249748
rect -960 245020 480 245260
rect 583520 236588 584960 236828
rect -960 232372 480 232612
rect 583520 223804 584960 224044
rect -960 219860 480 220100
rect 583520 211020 584960 211260
rect -960 207212 480 207452
rect 583520 198236 584960 198476
rect -960 194700 480 194940
rect 583520 185452 584960 185692
rect -960 182188 480 182428
rect 583520 172668 584960 172908
rect -960 169540 480 169780
rect 583520 159884 584960 160124
rect -960 157028 480 157268
rect 583520 147100 584960 147340
rect -960 144380 480 144620
rect 583520 134316 584960 134556
rect -960 131868 480 132108
rect 583520 121396 584960 121636
rect -960 119220 480 119460
rect 583520 108612 584960 108852
rect -960 106708 480 106948
rect 583520 95828 584960 96068
rect -960 94196 480 94436
rect 583520 83044 584960 83284
rect -960 81548 480 81788
rect 583520 70260 584960 70500
rect -960 69036 480 69276
rect 583520 57476 584960 57716
rect -960 56388 480 56628
rect 583520 44692 584960 44932
rect -960 43876 480 44116
rect 583520 31908 584960 32148
rect -960 31228 480 31468
rect 583520 19124 584960 19364
rect -960 18716 480 18956
rect -960 6204 480 6444
rect 583520 6340 584960 6580
<< obsm3 >>
rect 560 684900 583520 685133
rect 246 684892 583520 684900
rect 246 684492 583440 684892
rect 246 672652 583520 684492
rect 560 672252 583520 672652
rect 246 672108 583520 672252
rect 246 671708 583440 672108
rect 246 660140 583520 671708
rect 560 659740 583520 660140
rect 246 659324 583520 659740
rect 246 658924 583440 659324
rect 246 647492 583520 658924
rect 560 647092 583520 647492
rect 246 646540 583520 647092
rect 246 646140 583440 646540
rect 246 634980 583520 646140
rect 560 634580 583520 634980
rect 246 633756 583520 634580
rect 246 633356 583440 633756
rect 246 622468 583520 633356
rect 560 622068 583520 622468
rect 246 620972 583520 622068
rect 246 620572 583440 620972
rect 246 609820 583520 620572
rect 560 609420 583520 609820
rect 246 608188 583520 609420
rect 246 607788 583440 608188
rect 246 597308 583520 607788
rect 560 596908 583520 597308
rect 246 595404 583520 596908
rect 246 595004 583440 595404
rect 246 584660 583520 595004
rect 560 584260 583520 584660
rect 246 582484 583520 584260
rect 246 582084 583440 582484
rect 246 572148 583520 582084
rect 560 571748 583520 572148
rect 246 569700 583520 571748
rect 246 569300 583440 569700
rect 246 559500 583520 569300
rect 560 559100 583520 559500
rect 246 556916 583520 559100
rect 246 556516 583440 556916
rect 246 546988 583520 556516
rect 560 546588 583520 546988
rect 246 544132 583520 546588
rect 246 543732 583440 544132
rect 246 534476 583520 543732
rect 560 534076 583520 534476
rect 246 531348 583520 534076
rect 246 530948 583440 531348
rect 246 521828 583520 530948
rect 560 521428 583520 521828
rect 246 518564 583520 521428
rect 246 518164 583440 518564
rect 246 509316 583520 518164
rect 560 508916 583520 509316
rect 246 505780 583520 508916
rect 246 505380 583440 505780
rect 246 496668 583520 505380
rect 560 496268 583520 496668
rect 246 492996 583520 496268
rect 246 492596 583440 492996
rect 246 484156 583520 492596
rect 560 483756 583520 484156
rect 246 480212 583520 483756
rect 246 479812 583440 480212
rect 246 471508 583520 479812
rect 560 471108 583520 471508
rect 246 467292 583520 471108
rect 246 466892 583440 467292
rect 246 458996 583520 466892
rect 560 458596 583520 458996
rect 246 454508 583520 458596
rect 246 454108 583440 454508
rect 246 446484 583520 454108
rect 560 446084 583520 446484
rect 246 441724 583520 446084
rect 246 441324 583440 441724
rect 246 433836 583520 441324
rect 560 433436 583520 433836
rect 246 428940 583520 433436
rect 246 428540 583440 428940
rect 246 421324 583520 428540
rect 560 420924 583520 421324
rect 246 416156 583520 420924
rect 246 415756 583440 416156
rect 246 408676 583520 415756
rect 560 408276 583520 408676
rect 246 403372 583520 408276
rect 246 402972 583440 403372
rect 246 396164 583520 402972
rect 560 395764 583520 396164
rect 246 390588 583520 395764
rect 246 390188 583440 390588
rect 246 383516 583520 390188
rect 560 383116 583520 383516
rect 246 377804 583520 383116
rect 246 377404 583440 377804
rect 246 371004 583520 377404
rect 560 370604 583520 371004
rect 246 365020 583520 370604
rect 246 364620 583440 365020
rect 246 358492 583520 364620
rect 560 358092 583520 358492
rect 246 352100 583520 358092
rect 246 351700 583440 352100
rect 246 345844 583520 351700
rect 560 345444 583520 345844
rect 246 339316 583520 345444
rect 246 338916 583440 339316
rect 246 333332 583520 338916
rect 560 332932 583520 333332
rect 246 326532 583520 332932
rect 246 326132 583440 326532
rect 246 320684 583520 326132
rect 560 320284 583520 320684
rect 246 313748 583520 320284
rect 246 313348 583440 313748
rect 246 308172 583520 313348
rect 560 307772 583520 308172
rect 246 300964 583520 307772
rect 246 300564 583440 300964
rect 246 295524 583520 300564
rect 560 295124 583520 295524
rect 246 288180 583520 295124
rect 246 287780 583440 288180
rect 246 283012 583520 287780
rect 560 282612 583520 283012
rect 246 275396 583520 282612
rect 246 274996 583440 275396
rect 246 270500 583520 274996
rect 560 270100 583520 270500
rect 246 262612 583520 270100
rect 246 262212 583440 262612
rect 246 257852 583520 262212
rect 560 257452 583520 257852
rect 246 249828 583520 257452
rect 246 249428 583440 249828
rect 246 245340 583520 249428
rect 560 244940 583520 245340
rect 246 236908 583520 244940
rect 246 236508 583440 236908
rect 246 232692 583520 236508
rect 560 232292 583520 232692
rect 246 224124 583520 232292
rect 246 223724 583440 224124
rect 246 220180 583520 223724
rect 560 219780 583520 220180
rect 246 211340 583520 219780
rect 246 210940 583440 211340
rect 246 207532 583520 210940
rect 560 207132 583520 207532
rect 246 198556 583520 207132
rect 246 198156 583440 198556
rect 246 195020 583520 198156
rect 560 194620 583520 195020
rect 246 185772 583520 194620
rect 246 185372 583440 185772
rect 246 182508 583520 185372
rect 560 182108 583520 182508
rect 246 172988 583520 182108
rect 246 172588 583440 172988
rect 246 169860 583520 172588
rect 560 169460 583520 169860
rect 246 160204 583520 169460
rect 246 159804 583440 160204
rect 246 157348 583520 159804
rect 560 156948 583520 157348
rect 246 147420 583520 156948
rect 246 147020 583440 147420
rect 246 144700 583520 147020
rect 560 144300 583520 144700
rect 246 134636 583520 144300
rect 246 134236 583440 134636
rect 246 132188 583520 134236
rect 560 131788 583520 132188
rect 246 121716 583520 131788
rect 246 121316 583440 121716
rect 246 119540 583520 121316
rect 560 119140 583520 119540
rect 246 108932 583520 119140
rect 246 108532 583440 108932
rect 246 107028 583520 108532
rect 560 106628 583520 107028
rect 246 96148 583520 106628
rect 246 95748 583440 96148
rect 246 94516 583520 95748
rect 560 94116 583520 94516
rect 246 83364 583520 94116
rect 246 82964 583440 83364
rect 246 81868 583520 82964
rect 560 81468 583520 81868
rect 246 70580 583520 81468
rect 246 70180 583440 70580
rect 246 69356 583520 70180
rect 560 68956 583520 69356
rect 246 57796 583520 68956
rect 246 57396 583440 57796
rect 246 56708 583520 57396
rect 560 56308 583520 56708
rect 246 45012 583520 56308
rect 246 44612 583440 45012
rect 246 44196 583520 44612
rect 560 43796 583520 44196
rect 246 32228 583520 43796
rect 246 31828 583440 32228
rect 246 31548 583520 31828
rect 560 31315 583520 31548
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 -5734 9854 709670
rect 12954 -7654 13574 711590
rect 19794 -1894 20414 705830
rect 23514 -3814 24134 707750
rect 27234 -5734 27854 709670
rect 30954 -7654 31574 711590
rect 37794 -1894 38414 705830
rect 41514 -3814 42134 707750
rect 45234 -5734 45854 709670
rect 48954 -7654 49574 711590
rect 55794 -1894 56414 705830
rect 59514 640099 60134 707750
rect 63234 640099 63854 709670
rect 66954 640099 67574 711590
rect 73794 640099 74414 705830
rect 77514 640099 78134 707750
rect 81234 640099 81854 709670
rect 84954 640099 85574 711590
rect 91794 640099 92414 705830
rect 95514 640099 96134 707750
rect 99234 640099 99854 709670
rect 102954 640099 103574 711590
rect 109794 640099 110414 705830
rect 113514 640099 114134 707750
rect 117234 640099 117854 709670
rect 120954 640099 121574 711590
rect 59514 557000 60134 573000
rect 63234 557000 63854 573000
rect 66954 557000 67574 573000
rect 73794 557000 74414 573000
rect 77514 557000 78134 573000
rect 81234 557000 81854 573000
rect 84954 557000 85574 573000
rect 91794 557000 92414 573000
rect 95514 557000 96134 573000
rect 99234 557000 99854 573000
rect 102954 557000 103574 573000
rect 109794 557000 110414 573000
rect 113514 557000 114134 573000
rect 117234 557000 117854 573000
rect 120954 557000 121574 573000
rect 127794 557000 128414 705830
rect 131514 557000 132134 707750
rect 135234 557000 135854 709670
rect 138954 640099 139574 711590
rect 145794 640099 146414 705830
rect 149514 640099 150134 707750
rect 153234 640099 153854 709670
rect 156954 640099 157574 711590
rect 163794 640099 164414 705830
rect 167514 640099 168134 707750
rect 171234 640099 171854 709670
rect 174954 640099 175574 711590
rect 181794 640099 182414 705830
rect 185514 640099 186134 707750
rect 189234 640099 189854 709670
rect 192954 640099 193574 711590
rect 199794 640099 200414 705830
rect 138954 557000 139574 573000
rect 145794 557000 146414 573000
rect 149514 557000 150134 573000
rect 153234 557000 153854 573000
rect 156954 557000 157574 573000
rect 163794 557000 164414 573000
rect 167514 557000 168134 573000
rect 171234 557000 171854 573000
rect 174954 557000 175574 573000
rect 181794 557000 182414 573000
rect 185514 557000 186134 573000
rect 189234 557000 189854 573000
rect 192954 557000 193574 573000
rect 199794 557000 200414 573000
rect 203514 557000 204134 707750
rect 207234 557000 207854 709670
rect 210954 557000 211574 711590
rect 217794 640099 218414 705830
rect 221514 640099 222134 707750
rect 225234 640099 225854 709670
rect 228954 640099 229574 711590
rect 235794 640099 236414 705830
rect 239514 640099 240134 707750
rect 243234 640099 243854 709670
rect 246954 640099 247574 711590
rect 253794 640099 254414 705830
rect 257514 640099 258134 707750
rect 261234 640099 261854 709670
rect 264954 640099 265574 711590
rect 271794 640099 272414 705830
rect 275514 640099 276134 707750
rect 279234 640099 279854 709670
rect 282954 640099 283574 711590
rect 217794 557000 218414 573000
rect 221514 557000 222134 573000
rect 225234 557000 225854 573000
rect 228954 557000 229574 573000
rect 235794 557000 236414 573000
rect 239514 557000 240134 573000
rect 243234 557000 243854 573000
rect 246954 557000 247574 573000
rect 253794 557000 254414 573000
rect 257514 557000 258134 573000
rect 261234 557000 261854 573000
rect 264954 557000 265574 573000
rect 271794 557000 272414 573000
rect 275514 557000 276134 573000
rect 279234 557000 279854 573000
rect 282954 557000 283574 573000
rect 289794 557000 290414 705830
rect 293514 557000 294134 707750
rect 297234 557000 297854 709670
rect 300954 557000 301574 711590
rect 59514 460308 60134 493000
rect 63234 460308 63854 493000
rect 66954 460308 67574 493000
rect 73794 460308 74414 493000
rect 77514 460308 78134 493000
rect 81234 460308 81854 493000
rect 84954 460308 85574 493000
rect 91794 460308 92414 493000
rect 95514 460308 96134 493000
rect 99234 460308 99854 493000
rect 102954 460308 103574 493000
rect 109794 460308 110414 493000
rect 113514 460308 114134 493000
rect 117234 460308 117854 493000
rect 120954 460308 121574 493000
rect 127794 460308 128414 493000
rect 131514 460308 132134 493000
rect 135234 460308 135854 493000
rect 138954 460308 139574 493000
rect 145794 460308 146414 493000
rect 149514 460308 150134 493000
rect 153234 460308 153854 493000
rect 156954 460308 157574 493000
rect 163794 460308 164414 493000
rect 167514 460308 168134 493000
rect 171234 460308 171854 493000
rect 174954 460308 175574 493000
rect 181794 460308 182414 493000
rect 185514 460308 186134 493000
rect 189234 460308 189854 493000
rect 192954 460308 193574 493000
rect 59514 350308 60134 373000
rect 63234 350308 63854 373000
rect 66954 350308 67574 373000
rect 73794 350308 74414 373000
rect 77514 350308 78134 373000
rect 81234 350308 81854 373000
rect 84954 350308 85574 373000
rect 91794 350308 92414 373000
rect 95514 350308 96134 373000
rect 99234 350308 99854 373000
rect 102954 350308 103574 373000
rect 109794 350308 110414 373000
rect 113514 350308 114134 373000
rect 117234 350308 117854 373000
rect 120954 350308 121574 373000
rect 127794 350308 128414 373000
rect 131514 350308 132134 373000
rect 135234 350308 135854 373000
rect 138954 350308 139574 373000
rect 145794 350308 146414 373000
rect 149514 350308 150134 373000
rect 153234 350308 153854 373000
rect 156954 350308 157574 373000
rect 163794 350308 164414 373000
rect 167514 350308 168134 373000
rect 171234 350308 171854 373000
rect 174954 350308 175574 373000
rect 181794 350308 182414 373000
rect 185514 350308 186134 373000
rect 189234 350308 189854 373000
rect 192954 350308 193574 373000
rect 59514 240308 60134 263000
rect 63234 240308 63854 263000
rect 66954 240308 67574 263000
rect 73794 240308 74414 263000
rect 77514 240308 78134 263000
rect 81234 240308 81854 263000
rect 84954 240308 85574 263000
rect 91794 240308 92414 263000
rect 95514 240308 96134 263000
rect 99234 240308 99854 263000
rect 102954 240308 103574 263000
rect 109794 240308 110414 263000
rect 113514 240308 114134 263000
rect 117234 240308 117854 263000
rect 120954 240308 121574 263000
rect 127794 240308 128414 263000
rect 131514 240308 132134 263000
rect 135234 240308 135854 263000
rect 138954 240308 139574 263000
rect 145794 240308 146414 263000
rect 149514 240308 150134 263000
rect 153234 240308 153854 263000
rect 156954 240308 157574 263000
rect 163794 240308 164414 263000
rect 167514 240308 168134 263000
rect 171234 240308 171854 263000
rect 174954 240308 175574 263000
rect 181794 240308 182414 263000
rect 185514 240308 186134 263000
rect 189234 240308 189854 263000
rect 192954 240308 193574 263000
rect 59514 130308 60134 153000
rect 63234 130308 63854 153000
rect 66954 130308 67574 153000
rect 73794 130308 74414 153000
rect 77514 130308 78134 153000
rect 81234 130308 81854 153000
rect 84954 130308 85574 153000
rect 91794 130308 92414 153000
rect 95514 130308 96134 153000
rect 99234 130308 99854 153000
rect 102954 130308 103574 153000
rect 109794 130308 110414 153000
rect 113514 130308 114134 153000
rect 117234 130308 117854 153000
rect 120954 130308 121574 153000
rect 127794 130308 128414 153000
rect 131514 130308 132134 153000
rect 135234 130308 135854 153000
rect 138954 130308 139574 153000
rect 145794 130308 146414 153000
rect 149514 130308 150134 153000
rect 153234 130308 153854 153000
rect 156954 130308 157574 153000
rect 163794 130308 164414 153000
rect 167514 130308 168134 153000
rect 171234 130308 171854 153000
rect 174954 130308 175574 153000
rect 181794 130308 182414 153000
rect 185514 130308 186134 153000
rect 189234 130308 189854 153000
rect 192954 130308 193574 153000
rect 59514 -3814 60134 43000
rect 63234 -5734 63854 43000
rect 66954 -7654 67574 43000
rect 73794 -1894 74414 43000
rect 77514 -3814 78134 43000
rect 81234 -5734 81854 43000
rect 84954 -7654 85574 43000
rect 91794 -1894 92414 43000
rect 95514 -3814 96134 43000
rect 99234 -5734 99854 43000
rect 102954 -7654 103574 43000
rect 109794 -1894 110414 43000
rect 113514 -3814 114134 43000
rect 117234 -5734 117854 43000
rect 120954 -7654 121574 43000
rect 127794 -1894 128414 43000
rect 131514 -3814 132134 43000
rect 135234 -5734 135854 43000
rect 138954 -7654 139574 43000
rect 145794 -1894 146414 43000
rect 149514 -3814 150134 43000
rect 153234 -5734 153854 43000
rect 156954 -7654 157574 43000
rect 163794 -1894 164414 43000
rect 167514 -3814 168134 43000
rect 171234 -5734 171854 43000
rect 174954 -7654 175574 43000
rect 181794 -1894 182414 43000
rect 185514 -3814 186134 43000
rect 189234 -5734 189854 43000
rect 192954 -7654 193574 43000
rect 199794 -1894 200414 493000
rect 203514 -3814 204134 493000
rect 207234 -5734 207854 493000
rect 210954 -7654 211574 493000
rect 217794 460308 218414 493000
rect 221514 460308 222134 493000
rect 225234 460308 225854 493000
rect 228954 460308 229574 493000
rect 235794 460308 236414 493000
rect 239514 460308 240134 493000
rect 243234 460308 243854 493000
rect 246954 460308 247574 493000
rect 253794 460308 254414 493000
rect 257514 460308 258134 493000
rect 261234 460308 261854 493000
rect 264954 460308 265574 493000
rect 271794 460308 272414 493000
rect 275514 460308 276134 493000
rect 279234 460308 279854 493000
rect 282954 460308 283574 493000
rect 289794 460308 290414 493000
rect 293514 460308 294134 493000
rect 297234 460308 297854 493000
rect 300954 460308 301574 493000
rect 307794 460308 308414 705830
rect 311514 460308 312134 707750
rect 315234 460308 315854 709670
rect 318954 648033 319574 711590
rect 325794 648033 326414 705830
rect 329514 648033 330134 707750
rect 333234 648033 333854 709670
rect 336954 648033 337574 711590
rect 343794 648033 344414 705830
rect 347514 648033 348134 707750
rect 351234 648033 351854 709670
rect 354954 648033 355574 711590
rect 361794 648033 362414 705830
rect 365514 648033 366134 707750
rect 369234 648033 369854 709670
rect 372954 648033 373574 711590
rect 379794 648033 380414 705830
rect 383514 648033 384134 707750
rect 387234 648033 387854 709670
rect 390954 648033 391574 711590
rect 397794 648033 398414 705830
rect 401514 648033 402134 707750
rect 405234 648033 405854 709670
rect 408954 648033 409574 711590
rect 415794 648033 416414 705830
rect 419514 648033 420134 707750
rect 423234 648033 423854 709670
rect 426954 648033 427574 711590
rect 318954 460308 319574 533000
rect 325794 460308 326414 533000
rect 329514 460308 330134 533000
rect 333234 460308 333854 533000
rect 336954 460308 337574 533000
rect 343794 460308 344414 533000
rect 347514 460308 348134 533000
rect 351234 460308 351854 533000
rect 354954 460308 355574 533000
rect 217794 350308 218414 373000
rect 221514 350308 222134 373000
rect 225234 350308 225854 373000
rect 228954 350308 229574 373000
rect 235794 350308 236414 373000
rect 239514 350308 240134 373000
rect 243234 350308 243854 373000
rect 246954 350308 247574 373000
rect 253794 350308 254414 373000
rect 257514 350308 258134 373000
rect 261234 350308 261854 373000
rect 264954 350308 265574 373000
rect 271794 350308 272414 373000
rect 275514 350308 276134 373000
rect 279234 350308 279854 373000
rect 282954 350308 283574 373000
rect 289794 350308 290414 373000
rect 293514 350308 294134 373000
rect 297234 350308 297854 373000
rect 300954 350308 301574 373000
rect 307794 350308 308414 373000
rect 311514 350308 312134 373000
rect 315234 350308 315854 373000
rect 318954 350308 319574 373000
rect 325794 350308 326414 373000
rect 329514 350308 330134 373000
rect 333234 350308 333854 373000
rect 336954 350308 337574 373000
rect 343794 350308 344414 373000
rect 347514 350308 348134 373000
rect 351234 350308 351854 373000
rect 354954 350308 355574 373000
rect 217794 240308 218414 263000
rect 221514 240308 222134 263000
rect 225234 240308 225854 263000
rect 228954 240308 229574 263000
rect 235794 240308 236414 263000
rect 239514 240308 240134 263000
rect 243234 240308 243854 263000
rect 246954 240308 247574 263000
rect 253794 240308 254414 263000
rect 257514 240308 258134 263000
rect 261234 240308 261854 263000
rect 264954 240308 265574 263000
rect 271794 240308 272414 263000
rect 275514 240308 276134 263000
rect 279234 240308 279854 263000
rect 282954 240308 283574 263000
rect 289794 240308 290414 263000
rect 293514 240308 294134 263000
rect 297234 240308 297854 263000
rect 300954 240308 301574 263000
rect 307794 240308 308414 263000
rect 311514 240308 312134 263000
rect 315234 240308 315854 263000
rect 318954 240308 319574 263000
rect 325794 240308 326414 263000
rect 329514 240308 330134 263000
rect 333234 240308 333854 263000
rect 336954 240308 337574 263000
rect 343794 240308 344414 263000
rect 347514 240308 348134 263000
rect 351234 240308 351854 263000
rect 354954 240308 355574 263000
rect 217794 130308 218414 153000
rect 221514 130308 222134 153000
rect 225234 130308 225854 153000
rect 228954 130308 229574 153000
rect 235794 130308 236414 153000
rect 239514 130308 240134 153000
rect 243234 130308 243854 153000
rect 246954 130308 247574 153000
rect 253794 130308 254414 153000
rect 257514 130308 258134 153000
rect 261234 130308 261854 153000
rect 264954 130308 265574 153000
rect 271794 130308 272414 153000
rect 275514 130308 276134 153000
rect 279234 130308 279854 153000
rect 282954 130308 283574 153000
rect 289794 130308 290414 153000
rect 293514 130308 294134 153000
rect 297234 130308 297854 153000
rect 300954 130308 301574 153000
rect 307794 130308 308414 153000
rect 311514 130308 312134 153000
rect 315234 130308 315854 153000
rect 318954 130308 319574 153000
rect 325794 130308 326414 153000
rect 329514 130308 330134 153000
rect 333234 130308 333854 153000
rect 336954 130308 337574 153000
rect 343794 130308 344414 153000
rect 347514 130308 348134 153000
rect 351234 130308 351854 153000
rect 354954 130308 355574 153000
rect 217794 -1894 218414 43000
rect 221514 -3814 222134 43000
rect 225234 -5734 225854 43000
rect 228954 -7654 229574 43000
rect 235794 -1894 236414 43000
rect 239514 -3814 240134 43000
rect 243234 -5734 243854 43000
rect 246954 -7654 247574 43000
rect 253794 -1894 254414 43000
rect 257514 -3814 258134 43000
rect 261234 -5734 261854 43000
rect 264954 -7654 265574 43000
rect 271794 -1894 272414 43000
rect 275514 -3814 276134 43000
rect 279234 -5734 279854 43000
rect 282954 -7654 283574 43000
rect 289794 -1894 290414 43000
rect 293514 -3814 294134 43000
rect 297234 -5734 297854 43000
rect 300954 -7654 301574 43000
rect 307794 -1894 308414 43000
rect 311514 -3814 312134 43000
rect 315234 -5734 315854 43000
rect 318954 -7654 319574 43000
rect 325794 -1894 326414 43000
rect 329514 -3814 330134 43000
rect 333234 -5734 333854 43000
rect 336954 -7654 337574 43000
rect 343794 -1894 344414 43000
rect 347514 -3814 348134 43000
rect 351234 -5734 351854 43000
rect 354954 -7654 355574 43000
rect 361794 -1894 362414 533000
rect 365514 -3814 366134 533000
rect 369234 -5734 369854 533000
rect 372954 -7654 373574 533000
rect 379794 460308 380414 533000
rect 383514 460308 384134 533000
rect 387234 460308 387854 533000
rect 390954 460308 391574 533000
rect 397794 460308 398414 533000
rect 401514 460308 402134 533000
rect 405234 460308 405854 533000
rect 408954 460308 409574 533000
rect 415794 460308 416414 533000
rect 419514 460308 420134 533000
rect 423234 460308 423854 533000
rect 426954 460308 427574 533000
rect 433794 460308 434414 705830
rect 437514 460308 438134 707750
rect 441234 460308 441854 709670
rect 444954 460308 445574 711590
rect 451794 460308 452414 705830
rect 455514 460308 456134 707750
rect 459234 637000 459854 709670
rect 462954 637000 463574 711590
rect 469794 637000 470414 705830
rect 473514 637000 474134 707750
rect 477234 637000 477854 709670
rect 480954 637000 481574 711590
rect 487794 637000 488414 705830
rect 491514 637000 492134 707750
rect 495234 637000 495854 709670
rect 498954 637000 499574 711590
rect 505794 637000 506414 705830
rect 509514 637000 510134 707750
rect 459234 460308 459854 583000
rect 462954 460308 463574 583000
rect 469794 460308 470414 583000
rect 473514 460308 474134 583000
rect 477234 460308 477854 583000
rect 480954 460308 481574 583000
rect 487794 460308 488414 583000
rect 491514 460308 492134 583000
rect 495234 460308 495854 583000
rect 498954 460308 499574 583000
rect 505794 460308 506414 583000
rect 509514 460308 510134 583000
rect 513234 460308 513854 709670
rect 516954 460308 517574 711590
rect 379794 350308 380414 373000
rect 383514 350308 384134 373000
rect 387234 350308 387854 373000
rect 390954 350308 391574 373000
rect 397794 350308 398414 373000
rect 401514 350308 402134 373000
rect 405234 350308 405854 373000
rect 408954 350308 409574 373000
rect 415794 350308 416414 373000
rect 419514 350308 420134 373000
rect 423234 350308 423854 373000
rect 426954 350308 427574 373000
rect 433794 350308 434414 373000
rect 437514 350308 438134 373000
rect 441234 350308 441854 373000
rect 444954 350308 445574 373000
rect 451794 350308 452414 373000
rect 455514 350308 456134 373000
rect 459234 350308 459854 373000
rect 462954 350308 463574 373000
rect 469794 350308 470414 373000
rect 473514 350308 474134 373000
rect 477234 350308 477854 373000
rect 480954 350308 481574 373000
rect 487794 350308 488414 373000
rect 491514 350308 492134 373000
rect 495234 350308 495854 373000
rect 498954 350308 499574 373000
rect 505794 350308 506414 373000
rect 509514 350308 510134 373000
rect 513234 350308 513854 373000
rect 516954 350308 517574 373000
rect 379794 240308 380414 263000
rect 383514 240308 384134 263000
rect 387234 240308 387854 263000
rect 390954 240308 391574 263000
rect 397794 240308 398414 263000
rect 401514 240308 402134 263000
rect 405234 240308 405854 263000
rect 408954 240308 409574 263000
rect 415794 240308 416414 263000
rect 419514 240308 420134 263000
rect 423234 240308 423854 263000
rect 426954 240308 427574 263000
rect 433794 240308 434414 263000
rect 437514 240308 438134 263000
rect 441234 240308 441854 263000
rect 444954 240308 445574 263000
rect 451794 240308 452414 263000
rect 455514 240308 456134 263000
rect 459234 240308 459854 263000
rect 462954 240308 463574 263000
rect 469794 240308 470414 263000
rect 473514 240308 474134 263000
rect 477234 240308 477854 263000
rect 480954 240308 481574 263000
rect 487794 240308 488414 263000
rect 491514 240308 492134 263000
rect 495234 240308 495854 263000
rect 498954 240308 499574 263000
rect 505794 240308 506414 263000
rect 509514 240308 510134 263000
rect 513234 240308 513854 263000
rect 516954 240308 517574 263000
rect 379794 130308 380414 153000
rect 383514 130308 384134 153000
rect 387234 130308 387854 153000
rect 390954 130308 391574 153000
rect 397794 130308 398414 153000
rect 401514 130308 402134 153000
rect 405234 130308 405854 153000
rect 408954 130308 409574 153000
rect 415794 130308 416414 153000
rect 419514 130308 420134 153000
rect 423234 130308 423854 153000
rect 426954 130308 427574 153000
rect 433794 130308 434414 153000
rect 437514 130308 438134 153000
rect 441234 130308 441854 153000
rect 444954 130308 445574 153000
rect 451794 130308 452414 153000
rect 455514 130308 456134 153000
rect 459234 130308 459854 153000
rect 462954 130308 463574 153000
rect 469794 130308 470414 153000
rect 473514 130308 474134 153000
rect 477234 130308 477854 153000
rect 480954 130308 481574 153000
rect 487794 130308 488414 153000
rect 491514 130308 492134 153000
rect 495234 130308 495854 153000
rect 498954 130308 499574 153000
rect 505794 130308 506414 153000
rect 509514 130308 510134 153000
rect 513234 130308 513854 153000
rect 516954 130308 517574 153000
rect 379794 -1894 380414 43000
rect 383514 -3814 384134 43000
rect 387234 -5734 387854 43000
rect 390954 -7654 391574 43000
rect 397794 -1894 398414 43000
rect 401514 -3814 402134 43000
rect 405234 -5734 405854 43000
rect 408954 -7654 409574 43000
rect 415794 -1894 416414 43000
rect 419514 -3814 420134 43000
rect 423234 -5734 423854 43000
rect 426954 -7654 427574 43000
rect 433794 -1894 434414 43000
rect 437514 -3814 438134 43000
rect 441234 -5734 441854 43000
rect 444954 -7654 445574 43000
rect 451794 -1894 452414 43000
rect 455514 -3814 456134 43000
rect 459234 -5734 459854 43000
rect 462954 -7654 463574 43000
rect 469794 -1894 470414 43000
rect 473514 -3814 474134 43000
rect 477234 -5734 477854 43000
rect 480954 -7654 481574 43000
rect 487794 -1894 488414 43000
rect 491514 -3814 492134 43000
rect 495234 -5734 495854 43000
rect 498954 -7654 499574 43000
rect 505794 -1894 506414 43000
rect 509514 -3814 510134 43000
rect 513234 -5734 513854 43000
rect 516954 -7654 517574 43000
rect 523794 -1894 524414 705830
rect 527514 -3814 528134 707750
rect 531234 -5734 531854 709670
rect 534954 -7654 535574 711590
rect 541794 -1894 542414 705830
rect 545514 -3814 546134 707750
rect 549234 -5734 549854 709670
rect 552954 -7654 553574 711590
rect 559794 -1894 560414 705830
rect 563514 -3814 564134 707750
rect 567234 -5734 567854 709670
rect 570954 -7654 571574 711590
rect 577794 -1894 578414 705830
rect 581514 -3814 582134 707750
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 44771 39883 45154 646237
rect 45934 39883 48874 646237
rect 49654 39883 55714 646237
rect 56494 640019 59434 646237
rect 60214 640019 63154 646237
rect 63934 640019 66874 646237
rect 67654 640019 73714 646237
rect 74494 640019 77434 646237
rect 78214 640019 81154 646237
rect 81934 640019 84874 646237
rect 85654 640019 91714 646237
rect 92494 640019 95434 646237
rect 96214 640019 99154 646237
rect 99934 640019 102874 646237
rect 103654 640019 109714 646237
rect 110494 640019 113434 646237
rect 114214 640019 117154 646237
rect 117934 640019 120874 646237
rect 121654 640019 127714 646237
rect 56494 573080 127714 640019
rect 56494 556920 59434 573080
rect 60214 556920 63154 573080
rect 63934 556920 66874 573080
rect 67654 556920 73714 573080
rect 74494 556920 77434 573080
rect 78214 556920 81154 573080
rect 81934 556920 84874 573080
rect 85654 556920 91714 573080
rect 92494 556920 95434 573080
rect 96214 556920 99154 573080
rect 99934 556920 102874 573080
rect 103654 556920 109714 573080
rect 110494 556920 113434 573080
rect 114214 556920 117154 573080
rect 117934 556920 120874 573080
rect 121654 556920 127714 573080
rect 128494 556920 131434 646237
rect 132214 556920 135154 646237
rect 135934 640019 138874 646237
rect 139654 640019 145714 646237
rect 146494 640019 149434 646237
rect 150214 640019 153154 646237
rect 153934 640019 156874 646237
rect 157654 640019 163714 646237
rect 164494 640019 167434 646237
rect 168214 640019 171154 646237
rect 171934 640019 174874 646237
rect 175654 640019 181714 646237
rect 182494 640019 185434 646237
rect 186214 640019 189154 646237
rect 189934 640019 192874 646237
rect 193654 640019 199714 646237
rect 200494 640019 203434 646237
rect 135934 573080 203434 640019
rect 135934 556920 138874 573080
rect 139654 556920 145714 573080
rect 146494 556920 149434 573080
rect 150214 556920 153154 573080
rect 153934 556920 156874 573080
rect 157654 556920 163714 573080
rect 164494 556920 167434 573080
rect 168214 556920 171154 573080
rect 171934 556920 174874 573080
rect 175654 556920 181714 573080
rect 182494 556920 185434 573080
rect 186214 556920 189154 573080
rect 189934 556920 192874 573080
rect 193654 556920 199714 573080
rect 200494 556920 203434 573080
rect 204214 556920 207154 646237
rect 207934 556920 210874 646237
rect 211654 640019 217714 646237
rect 218494 640019 221434 646237
rect 222214 640019 225154 646237
rect 225934 640019 228874 646237
rect 229654 640019 235714 646237
rect 236494 640019 239434 646237
rect 240214 640019 243154 646237
rect 243934 640019 246874 646237
rect 247654 640019 253714 646237
rect 254494 640019 257434 646237
rect 258214 640019 261154 646237
rect 261934 640019 264874 646237
rect 265654 640019 271714 646237
rect 272494 640019 275434 646237
rect 276214 640019 279154 646237
rect 279934 640019 282874 646237
rect 283654 640019 289714 646237
rect 211654 573080 289714 640019
rect 211654 556920 217714 573080
rect 218494 556920 221434 573080
rect 222214 556920 225154 573080
rect 225934 556920 228874 573080
rect 229654 556920 235714 573080
rect 236494 556920 239434 573080
rect 240214 556920 243154 573080
rect 243934 556920 246874 573080
rect 247654 556920 253714 573080
rect 254494 556920 257434 573080
rect 258214 556920 261154 573080
rect 261934 556920 264874 573080
rect 265654 556920 271714 573080
rect 272494 556920 275434 573080
rect 276214 556920 279154 573080
rect 279934 556920 282874 573080
rect 283654 556920 289714 573080
rect 290494 556920 293434 646237
rect 294214 556920 297154 646237
rect 297934 556920 300874 646237
rect 301654 556920 307714 646237
rect 56494 493080 307714 556920
rect 56494 460228 59434 493080
rect 60214 460228 63154 493080
rect 63934 460228 66874 493080
rect 67654 460228 73714 493080
rect 74494 460228 77434 493080
rect 78214 460228 81154 493080
rect 81934 460228 84874 493080
rect 85654 460228 91714 493080
rect 92494 460228 95434 493080
rect 96214 460228 99154 493080
rect 99934 460228 102874 493080
rect 103654 460228 109714 493080
rect 110494 460228 113434 493080
rect 114214 460228 117154 493080
rect 117934 460228 120874 493080
rect 121654 460228 127714 493080
rect 128494 460228 131434 493080
rect 132214 460228 135154 493080
rect 135934 460228 138874 493080
rect 139654 460228 145714 493080
rect 146494 460228 149434 493080
rect 150214 460228 153154 493080
rect 153934 460228 156874 493080
rect 157654 460228 163714 493080
rect 164494 460228 167434 493080
rect 168214 460228 171154 493080
rect 171934 460228 174874 493080
rect 175654 460228 181714 493080
rect 182494 460228 185434 493080
rect 186214 460228 189154 493080
rect 189934 460228 192874 493080
rect 193654 460228 199714 493080
rect 56494 373080 199714 460228
rect 56494 350228 59434 373080
rect 60214 350228 63154 373080
rect 63934 350228 66874 373080
rect 67654 350228 73714 373080
rect 74494 350228 77434 373080
rect 78214 350228 81154 373080
rect 81934 350228 84874 373080
rect 85654 350228 91714 373080
rect 92494 350228 95434 373080
rect 96214 350228 99154 373080
rect 99934 350228 102874 373080
rect 103654 350228 109714 373080
rect 110494 350228 113434 373080
rect 114214 350228 117154 373080
rect 117934 350228 120874 373080
rect 121654 350228 127714 373080
rect 128494 350228 131434 373080
rect 132214 350228 135154 373080
rect 135934 350228 138874 373080
rect 139654 350228 145714 373080
rect 146494 350228 149434 373080
rect 150214 350228 153154 373080
rect 153934 350228 156874 373080
rect 157654 350228 163714 373080
rect 164494 350228 167434 373080
rect 168214 350228 171154 373080
rect 171934 350228 174874 373080
rect 175654 350228 181714 373080
rect 182494 350228 185434 373080
rect 186214 350228 189154 373080
rect 189934 350228 192874 373080
rect 193654 350228 199714 373080
rect 56494 263080 199714 350228
rect 56494 240228 59434 263080
rect 60214 240228 63154 263080
rect 63934 240228 66874 263080
rect 67654 240228 73714 263080
rect 74494 240228 77434 263080
rect 78214 240228 81154 263080
rect 81934 240228 84874 263080
rect 85654 240228 91714 263080
rect 92494 240228 95434 263080
rect 96214 240228 99154 263080
rect 99934 240228 102874 263080
rect 103654 240228 109714 263080
rect 110494 240228 113434 263080
rect 114214 240228 117154 263080
rect 117934 240228 120874 263080
rect 121654 240228 127714 263080
rect 128494 240228 131434 263080
rect 132214 240228 135154 263080
rect 135934 240228 138874 263080
rect 139654 240228 145714 263080
rect 146494 240228 149434 263080
rect 150214 240228 153154 263080
rect 153934 240228 156874 263080
rect 157654 240228 163714 263080
rect 164494 240228 167434 263080
rect 168214 240228 171154 263080
rect 171934 240228 174874 263080
rect 175654 240228 181714 263080
rect 182494 240228 185434 263080
rect 186214 240228 189154 263080
rect 189934 240228 192874 263080
rect 193654 240228 199714 263080
rect 56494 153080 199714 240228
rect 56494 130228 59434 153080
rect 60214 130228 63154 153080
rect 63934 130228 66874 153080
rect 67654 130228 73714 153080
rect 74494 130228 77434 153080
rect 78214 130228 81154 153080
rect 81934 130228 84874 153080
rect 85654 130228 91714 153080
rect 92494 130228 95434 153080
rect 96214 130228 99154 153080
rect 99934 130228 102874 153080
rect 103654 130228 109714 153080
rect 110494 130228 113434 153080
rect 114214 130228 117154 153080
rect 117934 130228 120874 153080
rect 121654 130228 127714 153080
rect 128494 130228 131434 153080
rect 132214 130228 135154 153080
rect 135934 130228 138874 153080
rect 139654 130228 145714 153080
rect 146494 130228 149434 153080
rect 150214 130228 153154 153080
rect 153934 130228 156874 153080
rect 157654 130228 163714 153080
rect 164494 130228 167434 153080
rect 168214 130228 171154 153080
rect 171934 130228 174874 153080
rect 175654 130228 181714 153080
rect 182494 130228 185434 153080
rect 186214 130228 189154 153080
rect 189934 130228 192874 153080
rect 193654 130228 199714 153080
rect 56494 43080 199714 130228
rect 56494 39883 59434 43080
rect 60214 39883 63154 43080
rect 63934 39883 66874 43080
rect 67654 39883 73714 43080
rect 74494 39883 77434 43080
rect 78214 39883 81154 43080
rect 81934 39883 84874 43080
rect 85654 39883 91714 43080
rect 92494 39883 95434 43080
rect 96214 39883 99154 43080
rect 99934 39883 102874 43080
rect 103654 39883 109714 43080
rect 110494 39883 113434 43080
rect 114214 39883 117154 43080
rect 117934 39883 120874 43080
rect 121654 39883 127714 43080
rect 128494 39883 131434 43080
rect 132214 39883 135154 43080
rect 135934 39883 138874 43080
rect 139654 39883 145714 43080
rect 146494 39883 149434 43080
rect 150214 39883 153154 43080
rect 153934 39883 156874 43080
rect 157654 39883 163714 43080
rect 164494 39883 167434 43080
rect 168214 39883 171154 43080
rect 171934 39883 174874 43080
rect 175654 39883 181714 43080
rect 182494 39883 185434 43080
rect 186214 39883 189154 43080
rect 189934 39883 192874 43080
rect 193654 39883 199714 43080
rect 200494 39883 203434 493080
rect 204214 39883 207154 493080
rect 207934 39883 210874 493080
rect 211654 460228 217714 493080
rect 218494 460228 221434 493080
rect 222214 460228 225154 493080
rect 225934 460228 228874 493080
rect 229654 460228 235714 493080
rect 236494 460228 239434 493080
rect 240214 460228 243154 493080
rect 243934 460228 246874 493080
rect 247654 460228 253714 493080
rect 254494 460228 257434 493080
rect 258214 460228 261154 493080
rect 261934 460228 264874 493080
rect 265654 460228 271714 493080
rect 272494 460228 275434 493080
rect 276214 460228 279154 493080
rect 279934 460228 282874 493080
rect 283654 460228 289714 493080
rect 290494 460228 293434 493080
rect 294214 460228 297154 493080
rect 297934 460228 300874 493080
rect 301654 460228 307714 493080
rect 308494 460228 311434 646237
rect 312214 460228 315154 646237
rect 315934 533080 433714 646237
rect 315934 460228 318874 533080
rect 319654 460228 325714 533080
rect 326494 460228 329434 533080
rect 330214 460228 333154 533080
rect 333934 460228 336874 533080
rect 337654 460228 343714 533080
rect 344494 460228 347434 533080
rect 348214 460228 351154 533080
rect 351934 460228 354874 533080
rect 355654 460228 361714 533080
rect 211654 373080 361714 460228
rect 211654 350228 217714 373080
rect 218494 350228 221434 373080
rect 222214 350228 225154 373080
rect 225934 350228 228874 373080
rect 229654 350228 235714 373080
rect 236494 350228 239434 373080
rect 240214 350228 243154 373080
rect 243934 350228 246874 373080
rect 247654 350228 253714 373080
rect 254494 350228 257434 373080
rect 258214 350228 261154 373080
rect 261934 350228 264874 373080
rect 265654 350228 271714 373080
rect 272494 350228 275434 373080
rect 276214 350228 279154 373080
rect 279934 350228 282874 373080
rect 283654 350228 289714 373080
rect 290494 350228 293434 373080
rect 294214 350228 297154 373080
rect 297934 350228 300874 373080
rect 301654 350228 307714 373080
rect 308494 350228 311434 373080
rect 312214 350228 315154 373080
rect 315934 350228 318874 373080
rect 319654 350228 325714 373080
rect 326494 350228 329434 373080
rect 330214 350228 333154 373080
rect 333934 350228 336874 373080
rect 337654 350228 343714 373080
rect 344494 350228 347434 373080
rect 348214 350228 351154 373080
rect 351934 350228 354874 373080
rect 355654 350228 361714 373080
rect 211654 263080 361714 350228
rect 211654 240228 217714 263080
rect 218494 240228 221434 263080
rect 222214 240228 225154 263080
rect 225934 240228 228874 263080
rect 229654 240228 235714 263080
rect 236494 240228 239434 263080
rect 240214 240228 243154 263080
rect 243934 240228 246874 263080
rect 247654 240228 253714 263080
rect 254494 240228 257434 263080
rect 258214 240228 261154 263080
rect 261934 240228 264874 263080
rect 265654 240228 271714 263080
rect 272494 240228 275434 263080
rect 276214 240228 279154 263080
rect 279934 240228 282874 263080
rect 283654 240228 289714 263080
rect 290494 240228 293434 263080
rect 294214 240228 297154 263080
rect 297934 240228 300874 263080
rect 301654 240228 307714 263080
rect 308494 240228 311434 263080
rect 312214 240228 315154 263080
rect 315934 240228 318874 263080
rect 319654 240228 325714 263080
rect 326494 240228 329434 263080
rect 330214 240228 333154 263080
rect 333934 240228 336874 263080
rect 337654 240228 343714 263080
rect 344494 240228 347434 263080
rect 348214 240228 351154 263080
rect 351934 240228 354874 263080
rect 355654 240228 361714 263080
rect 211654 153080 361714 240228
rect 211654 130228 217714 153080
rect 218494 130228 221434 153080
rect 222214 130228 225154 153080
rect 225934 130228 228874 153080
rect 229654 130228 235714 153080
rect 236494 130228 239434 153080
rect 240214 130228 243154 153080
rect 243934 130228 246874 153080
rect 247654 130228 253714 153080
rect 254494 130228 257434 153080
rect 258214 130228 261154 153080
rect 261934 130228 264874 153080
rect 265654 130228 271714 153080
rect 272494 130228 275434 153080
rect 276214 130228 279154 153080
rect 279934 130228 282874 153080
rect 283654 130228 289714 153080
rect 290494 130228 293434 153080
rect 294214 130228 297154 153080
rect 297934 130228 300874 153080
rect 301654 130228 307714 153080
rect 308494 130228 311434 153080
rect 312214 130228 315154 153080
rect 315934 130228 318874 153080
rect 319654 130228 325714 153080
rect 326494 130228 329434 153080
rect 330214 130228 333154 153080
rect 333934 130228 336874 153080
rect 337654 130228 343714 153080
rect 344494 130228 347434 153080
rect 348214 130228 351154 153080
rect 351934 130228 354874 153080
rect 355654 130228 361714 153080
rect 211654 43080 361714 130228
rect 211654 39883 217714 43080
rect 218494 39883 221434 43080
rect 222214 39883 225154 43080
rect 225934 39883 228874 43080
rect 229654 39883 235714 43080
rect 236494 39883 239434 43080
rect 240214 39883 243154 43080
rect 243934 39883 246874 43080
rect 247654 39883 253714 43080
rect 254494 39883 257434 43080
rect 258214 39883 261154 43080
rect 261934 39883 264874 43080
rect 265654 39883 271714 43080
rect 272494 39883 275434 43080
rect 276214 39883 279154 43080
rect 279934 39883 282874 43080
rect 283654 39883 289714 43080
rect 290494 39883 293434 43080
rect 294214 39883 297154 43080
rect 297934 39883 300874 43080
rect 301654 39883 307714 43080
rect 308494 39883 311434 43080
rect 312214 39883 315154 43080
rect 315934 39883 318874 43080
rect 319654 39883 325714 43080
rect 326494 39883 329434 43080
rect 330214 39883 333154 43080
rect 333934 39883 336874 43080
rect 337654 39883 343714 43080
rect 344494 39883 347434 43080
rect 348214 39883 351154 43080
rect 351934 39883 354874 43080
rect 355654 39883 361714 43080
rect 362494 39883 365434 533080
rect 366214 39883 369154 533080
rect 369934 39883 372874 533080
rect 373654 460228 379714 533080
rect 380494 460228 383434 533080
rect 384214 460228 387154 533080
rect 387934 460228 390874 533080
rect 391654 460228 397714 533080
rect 398494 460228 401434 533080
rect 402214 460228 405154 533080
rect 405934 460228 408874 533080
rect 409654 460228 415714 533080
rect 416494 460228 419434 533080
rect 420214 460228 423154 533080
rect 423934 460228 426874 533080
rect 427654 460228 433714 533080
rect 434494 460228 437434 646237
rect 438214 460228 441154 646237
rect 441934 460228 444874 646237
rect 445654 460228 451714 646237
rect 452494 460228 455434 646237
rect 456214 636920 459154 646237
rect 459934 636920 462874 646237
rect 463654 636920 469714 646237
rect 470494 636920 473434 646237
rect 474214 636920 477154 646237
rect 477934 636920 480874 646237
rect 481654 636920 487714 646237
rect 488494 636920 491434 646237
rect 492214 636920 495154 646237
rect 495934 636920 498874 646237
rect 499654 636920 505714 646237
rect 506494 636920 509434 646237
rect 510214 636920 513154 646237
rect 456214 583080 513154 636920
rect 456214 460228 459154 583080
rect 459934 460228 462874 583080
rect 463654 460228 469714 583080
rect 470494 460228 473434 583080
rect 474214 460228 477154 583080
rect 477934 460228 480874 583080
rect 481654 460228 487714 583080
rect 488494 460228 491434 583080
rect 492214 460228 495154 583080
rect 495934 460228 498874 583080
rect 499654 460228 505714 583080
rect 506494 460228 509434 583080
rect 510214 460228 513154 583080
rect 513934 460228 516496 646237
rect 373654 373080 516496 460228
rect 373654 350228 379714 373080
rect 380494 350228 383434 373080
rect 384214 350228 387154 373080
rect 387934 350228 390874 373080
rect 391654 350228 397714 373080
rect 398494 350228 401434 373080
rect 402214 350228 405154 373080
rect 405934 350228 408874 373080
rect 409654 350228 415714 373080
rect 416494 350228 419434 373080
rect 420214 350228 423154 373080
rect 423934 350228 426874 373080
rect 427654 350228 433714 373080
rect 434494 350228 437434 373080
rect 438214 350228 441154 373080
rect 441934 350228 444874 373080
rect 445654 350228 451714 373080
rect 452494 350228 455434 373080
rect 456214 350228 459154 373080
rect 459934 350228 462874 373080
rect 463654 350228 469714 373080
rect 470494 350228 473434 373080
rect 474214 350228 477154 373080
rect 477934 350228 480874 373080
rect 481654 350228 487714 373080
rect 488494 350228 491434 373080
rect 492214 350228 495154 373080
rect 495934 350228 498874 373080
rect 499654 350228 505714 373080
rect 506494 350228 509434 373080
rect 510214 350228 513154 373080
rect 513934 350228 516496 373080
rect 373654 263080 516496 350228
rect 373654 240228 379714 263080
rect 380494 240228 383434 263080
rect 384214 240228 387154 263080
rect 387934 240228 390874 263080
rect 391654 240228 397714 263080
rect 398494 240228 401434 263080
rect 402214 240228 405154 263080
rect 405934 240228 408874 263080
rect 409654 240228 415714 263080
rect 416494 240228 419434 263080
rect 420214 240228 423154 263080
rect 423934 240228 426874 263080
rect 427654 240228 433714 263080
rect 434494 240228 437434 263080
rect 438214 240228 441154 263080
rect 441934 240228 444874 263080
rect 445654 240228 451714 263080
rect 452494 240228 455434 263080
rect 456214 240228 459154 263080
rect 459934 240228 462874 263080
rect 463654 240228 469714 263080
rect 470494 240228 473434 263080
rect 474214 240228 477154 263080
rect 477934 240228 480874 263080
rect 481654 240228 487714 263080
rect 488494 240228 491434 263080
rect 492214 240228 495154 263080
rect 495934 240228 498874 263080
rect 499654 240228 505714 263080
rect 506494 240228 509434 263080
rect 510214 240228 513154 263080
rect 513934 240228 516496 263080
rect 373654 153080 516496 240228
rect 373654 130228 379714 153080
rect 380494 130228 383434 153080
rect 384214 130228 387154 153080
rect 387934 130228 390874 153080
rect 391654 130228 397714 153080
rect 398494 130228 401434 153080
rect 402214 130228 405154 153080
rect 405934 130228 408874 153080
rect 409654 130228 415714 153080
rect 416494 130228 419434 153080
rect 420214 130228 423154 153080
rect 423934 130228 426874 153080
rect 427654 130228 433714 153080
rect 434494 130228 437434 153080
rect 438214 130228 441154 153080
rect 441934 130228 444874 153080
rect 445654 130228 451714 153080
rect 452494 130228 455434 153080
rect 456214 130228 459154 153080
rect 459934 130228 462874 153080
rect 463654 130228 469714 153080
rect 470494 130228 473434 153080
rect 474214 130228 477154 153080
rect 477934 130228 480874 153080
rect 481654 130228 487714 153080
rect 488494 130228 491434 153080
rect 492214 130228 495154 153080
rect 495934 130228 498874 153080
rect 499654 130228 505714 153080
rect 506494 130228 509434 153080
rect 510214 130228 513154 153080
rect 513934 130228 516496 153080
rect 373654 43080 516496 130228
rect 373654 39883 379714 43080
rect 380494 39883 383434 43080
rect 384214 39883 387154 43080
rect 387934 39883 390874 43080
rect 391654 39883 397714 43080
rect 398494 39883 401434 43080
rect 402214 39883 405154 43080
rect 405934 39883 408874 43080
rect 409654 39883 415714 43080
rect 416494 39883 419434 43080
rect 420214 39883 423154 43080
rect 423934 39883 426874 43080
rect 427654 39883 433714 43080
rect 434494 39883 437434 43080
rect 438214 39883 441154 43080
rect 441934 39883 444874 43080
rect 445654 39883 451714 43080
rect 452494 39883 455434 43080
rect 456214 39883 459154 43080
rect 459934 39883 462874 43080
rect 463654 39883 469714 43080
rect 470494 39883 473434 43080
rect 474214 39883 477154 43080
rect 477934 39883 480874 43080
rect 481654 39883 487714 43080
rect 488494 39883 491434 43080
rect 492214 39883 495154 43080
rect 495934 39883 498874 43080
rect 499654 39883 505714 43080
rect 506494 39883 509434 43080
rect 510214 39883 513154 43080
rect 513934 39883 516496 43080
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -6806 694306 590730 694926
rect -4886 690586 588810 691206
rect -2966 686866 586890 687486
rect -8726 680026 592650 680646
rect -6806 676306 590730 676926
rect -4886 672586 588810 673206
rect -2966 668866 586890 669486
rect -8726 662026 592650 662646
rect -6806 658306 590730 658926
rect -4886 654586 588810 655206
rect -2966 650866 586890 651486
rect -8726 644026 592650 644646
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -2966 632866 586890 633486
rect -8726 626026 592650 626646
rect -6806 622306 590730 622926
rect -4886 618586 588810 619206
rect -2966 614866 586890 615486
rect -8726 608026 592650 608646
rect -6806 604306 590730 604926
rect -4886 600586 588810 601206
rect -2966 596866 586890 597486
rect -8726 590026 592650 590646
rect -6806 586306 590730 586926
rect -4886 582586 588810 583206
rect -2966 578866 586890 579486
rect -8726 572026 592650 572646
rect 84954 571086 265574 571706
rect -6806 568306 590730 568926
rect 81234 567366 261854 567986
rect 77514 565526 258134 566146
rect -4886 564586 588810 565206
rect 73794 561806 254414 562426
rect -2966 560866 586890 561486
rect -8726 554026 592650 554646
rect -6806 550306 590730 550926
rect -4886 546586 588810 547206
rect -2966 542866 586890 543486
rect -8726 536026 592650 536646
rect -6806 532306 590730 532926
rect -4886 528586 588810 529206
rect -2966 524866 586890 525486
rect -8726 518026 592650 518646
rect -6806 514306 590730 514926
rect -4886 510586 588810 511206
rect -2966 506866 586890 507486
rect -8726 500026 592650 500646
rect -6806 496306 590730 496926
rect -4886 492586 588810 493206
rect -2966 488866 586890 489486
rect -8726 482026 592650 482646
rect -6806 478306 590730 478926
rect 63234 477366 279854 477986
rect 59514 475526 276134 476146
rect -4886 474586 588810 475206
rect -2966 470866 586890 471486
rect -8726 464026 592650 464646
rect -6806 460306 590730 460926
rect -4886 456586 588810 457206
rect -2966 452866 586890 453486
rect -8726 446026 592650 446646
rect -6806 442306 590730 442926
rect -4886 438586 588810 439206
rect -2966 434866 586890 435486
rect -8726 428026 592650 428646
rect -6806 424306 590730 424926
rect -4886 420586 588810 421206
rect -2966 416866 586890 417486
rect -8726 410026 592650 410646
rect -6806 406306 590730 406926
rect -4886 402586 588810 403206
rect -2966 398866 586890 399486
rect -8726 392026 592650 392646
rect -6806 388306 590730 388926
rect -4886 384586 588810 385206
rect -2966 380866 586890 381486
rect -8726 374026 592650 374646
rect -6806 370306 590730 370926
rect -4886 366586 588810 367206
rect 59514 365646 492134 366266
rect -2966 362866 586890 363486
rect 91794 361926 488414 362546
rect 84954 356966 517574 357586
rect -8726 356026 592650 356646
rect -6806 352306 590730 352926
rect -4886 348586 588810 349206
rect -2966 344866 586890 345486
rect -8726 338026 592650 338646
rect -6806 334306 590730 334926
rect -4886 330586 588810 331206
rect -2966 326866 586890 327486
rect -8726 320026 592650 320646
rect -6806 316306 590730 316926
rect -4886 312586 588810 313206
rect -2966 308866 586890 309486
rect -8726 302026 592650 302646
rect -6806 298306 590730 298926
rect -4886 294586 588810 295206
rect -2966 290866 586890 291486
rect -8726 284026 592650 284646
rect -6806 280306 590730 280926
rect -4886 276586 588810 277206
rect -2966 272866 586890 273486
rect -8726 266026 592650 266646
rect -6806 262306 590730 262926
rect -4886 258586 588810 259206
rect -2966 254866 586890 255486
rect 91794 253926 488414 254546
rect 84954 248966 517574 249586
rect -8726 248026 592650 248646
rect -6806 244306 590730 244926
rect -4886 240586 588810 241206
rect -2966 236866 586890 237486
rect -8726 230026 592650 230646
rect -6806 226306 590730 226926
rect -4886 222586 588810 223206
rect -2966 218866 586890 219486
rect -8726 212026 592650 212646
rect -6806 208306 590730 208926
rect -4886 204586 588810 205206
rect -2966 200866 586890 201486
rect -8726 194026 592650 194646
rect -6806 190306 590730 190926
rect -4886 186586 588810 187206
rect -2966 182866 586890 183486
rect -8726 176026 592650 176646
rect -6806 172306 590730 172926
rect -4886 168586 588810 169206
rect -2966 164866 586890 165486
rect -8726 158026 592650 158646
rect -6806 154306 590730 154926
rect -4886 150586 588810 151206
rect -2966 146866 586890 147486
rect 91794 145926 488414 146546
rect 84954 140966 517574 141586
rect -8726 140026 592650 140646
rect 81234 137246 513854 137866
rect -6806 136306 590730 136926
rect -4886 132586 588810 133206
rect -2966 128866 586890 129486
rect -8726 122026 592650 122646
rect -6806 118306 590730 118926
rect -4886 114586 588810 115206
rect -2966 110866 586890 111486
rect -8726 104026 592650 104646
rect -6806 100306 590730 100926
rect -4886 96586 588810 97206
rect -2966 92866 586890 93486
rect -8726 86026 592650 86646
rect -6806 82306 590730 82926
rect -4886 78586 588810 79206
rect -2966 74866 586890 75486
rect -8726 68026 592650 68646
rect -6806 64306 590730 64926
rect -4886 60586 588810 61206
rect -2966 56866 586890 57486
rect -8726 50026 592650 50646
rect -6806 46306 590730 46926
rect -4886 42586 588810 43206
rect -2966 38866 586890 39486
rect -8726 32026 592650 32646
rect -6806 28306 590730 28926
rect -4886 24586 588810 25206
rect -2966 20866 586890 21486
rect -8726 14026 592650 14646
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 275076 584960 275316 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 453274 703520 453386 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 391818 703520 391930 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 330362 703520 330474 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 268814 703520 268926 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 207358 703520 207470 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 145902 703520 146014 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 84446 703520 84558 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697492 480 697732 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 647172 480 647412 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 596988 480 597228 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 326212 584960 326452 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 546668 480 546908 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 496348 480 496588 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 446164 480 446404 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 395844 480 396084 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 345524 480 345764 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 295204 480 295444 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 245020 480 245260 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 194700 480 194940 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 144380 480 144620 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 377484 584960 377724 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 428620 584960 428860 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 479892 584960 480132 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 531028 584960 531268 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 582164 584960 582404 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 633436 584960 633676 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 576186 703520 576298 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 514730 703520 514842 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6340 584960 6580 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 441404 584960 441644 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 492676 584960 492916 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 543812 584960 544052 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 595084 584960 595324 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 646220 584960 646460 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 560822 703520 560934 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 499366 703520 499478 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 437910 703520 438022 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 376454 703520 376566 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 314998 703520 315110 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 44692 584960 44932 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 253450 703520 253562 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 191994 703520 192106 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 130538 703520 130650 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 69082 703520 69194 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684980 480 685220 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 634660 480 634900 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 584340 480 584580 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 534156 480 534396 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 483836 480 484076 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 433516 480 433756 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 83044 584960 83284 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 383196 480 383436 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 333012 480 333252 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 282692 480 282932 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 232372 480 232612 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 182188 480 182428 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 131868 480 132108 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 94196 480 94436 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 56388 480 56628 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 121396 584960 121636 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 159884 584960 160124 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 198236 584960 198476 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 236588 584960 236828 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 287860 584960 288100 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 338996 584960 339236 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 390268 584960 390508 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 31908 584960 32148 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 466972 584960 467212 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 518244 584960 518484 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 569380 584960 569620 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 620652 584960 620892 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 671788 584960 672028 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 530094 703520 530206 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 468638 703520 468750 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 407182 703520 407294 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 345726 703520 345838 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 284178 703520 284290 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 70260 584960 70500 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 222722 703520 222834 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 161266 703520 161378 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 99810 703520 99922 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 38354 703520 38466 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 659820 480 660060 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 609500 480 609740 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 559180 480 559420 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 508996 480 509236 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 458676 480 458916 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 408356 480 408596 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 108612 584960 108852 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 358172 480 358412 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 307852 480 308092 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 257532 480 257772 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 207212 480 207452 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 157028 480 157268 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 106708 480 106948 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 69036 480 69276 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 31228 480 31468 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 147100 584960 147340 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 185452 584960 185692 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 223804 584960 224044 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 262292 584960 262532 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 313428 584960 313668 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 364700 584960 364940 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 415836 584960 416076 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19124 584960 19364 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 454188 584960 454428 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 505460 584960 505700 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 556596 584960 556836 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 607868 584960 608108 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 659004 584960 659244 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 545458 703520 545570 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 484002 703520 484114 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 422546 703520 422658 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 361090 703520 361202 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 299634 703520 299746 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 57476 584960 57716 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 238086 703520 238198 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 176630 703520 176742 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 115174 703520 115286 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 53718 703520 53830 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 672332 480 672572 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 622148 480 622388 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 571828 480 572068 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 521508 480 521748 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 471188 480 471428 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 421004 480 421244 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 95828 584960 96068 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 370684 480 370924 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 320364 480 320604 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 270180 480 270420 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 219860 480 220100 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 169540 480 169780 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 119220 480 119460 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 81548 480 81788 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 43876 480 44116 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 134316 584960 134556 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 172668 584960 172908 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 211020 584960 211260 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 249508 584960 249748 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 300644 584960 300884 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 351780 584960 352020 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 403052 584960 403292 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125294 -960 125406 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 478574 -960 478686 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 482070 -960 482182 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 485566 -960 485678 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 489154 -960 489266 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 492650 -960 492762 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 496238 -960 496350 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 499734 -960 499846 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 503230 -960 503342 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 506818 -960 506930 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 510314 -960 510426 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 160622 -960 160734 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 513902 -960 514014 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 517398 -960 517510 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 520894 -960 521006 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 524482 -960 524594 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 527978 -960 528090 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 531566 -960 531678 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 535062 -960 535174 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 538558 -960 538670 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 542146 -960 542258 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 545642 -960 545754 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164118 -960 164230 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 549230 -960 549342 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 552726 -960 552838 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 556222 -960 556334 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 559810 -960 559922 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 563306 -960 563418 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 566894 -960 567006 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 570390 -960 570502 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 573886 -960 573998 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 167706 -960 167818 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171202 -960 171314 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 174790 -960 174902 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 178286 -960 178398 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 181782 -960 181894 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 185370 -960 185482 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 188866 -960 188978 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 192454 -960 192566 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 128882 -960 128994 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 195950 -960 196062 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 199446 -960 199558 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203034 -960 203146 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 206530 -960 206642 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210118 -960 210230 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 213614 -960 213726 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 217110 -960 217222 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 220698 -960 220810 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 224194 -960 224306 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 227782 -960 227894 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132378 -960 132490 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 231278 -960 231390 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 234774 -960 234886 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 238362 -960 238474 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 241858 -960 241970 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 245446 -960 245558 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 248942 -960 249054 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 252438 -960 252550 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 256026 -960 256138 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 259522 -960 259634 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 263110 -960 263222 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 135874 -960 135986 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 266606 -960 266718 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 270102 -960 270214 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 273690 -960 273802 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 277186 -960 277298 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 280774 -960 280886 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 298346 -960 298458 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 139462 -960 139574 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 305430 -960 305542 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 312514 -960 312626 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 316010 -960 316122 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 319598 -960 319710 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 323094 -960 323206 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 326682 -960 326794 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 330178 -960 330290 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 333674 -960 333786 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 142958 -960 143070 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 337262 -960 337374 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 340758 -960 340870 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 344346 -960 344458 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 358422 -960 358534 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 362010 -960 362122 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 365506 -960 365618 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 369002 -960 369114 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 146546 -960 146658 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 372590 -960 372702 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 376086 -960 376198 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 379674 -960 379786 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 383170 -960 383282 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 386666 -960 386778 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 390254 -960 390366 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 393750 -960 393862 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 397338 -960 397450 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 400834 -960 400946 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 404330 -960 404442 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150042 -960 150154 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 407918 -960 408030 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 411414 -960 411526 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 415002 -960 415114 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 418498 -960 418610 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 421994 -960 422106 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 425582 -960 425694 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 429078 -960 429190 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 432666 -960 432778 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 436162 -960 436274 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 439658 -960 439770 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 153538 -960 153650 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 443246 -960 443358 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 446742 -960 446854 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 450238 -960 450350 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 453826 -960 453938 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 457322 -960 457434 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 460910 -960 461022 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 474986 -960 475098 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157126 -960 157238 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126490 -960 126602 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 479678 -960 479790 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 483266 -960 483378 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 486762 -960 486874 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 490350 -960 490462 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 493846 -960 493958 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 497342 -960 497454 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 500930 -960 501042 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 504426 -960 504538 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 508014 -960 508126 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 511510 -960 511622 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 161818 -960 161930 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 515006 -960 515118 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 518594 -960 518706 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 522090 -960 522202 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 525678 -960 525790 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 529174 -960 529286 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 532670 -960 532782 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 536258 -960 536370 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 539754 -960 539866 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 543342 -960 543454 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 546838 -960 546950 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 165314 -960 165426 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 550334 -960 550446 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 553922 -960 554034 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 557418 -960 557530 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 561006 -960 561118 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 564502 -960 564614 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 567998 -960 568110 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 571586 -960 571698 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 575082 -960 575194 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 168902 -960 169014 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 172398 -960 172510 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 175894 -960 176006 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 179482 -960 179594 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 182978 -960 183090 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 186566 -960 186678 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190062 -960 190174 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 193558 -960 193670 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 129986 -960 130098 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197146 -960 197258 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 200642 -960 200754 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 204230 -960 204342 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 207726 -960 207838 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 211222 -960 211334 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 214810 -960 214922 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 218306 -960 218418 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 221894 -960 222006 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 225390 -960 225502 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 228886 -960 228998 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 133574 -960 133686 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 232474 -960 232586 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 235970 -960 236082 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 239558 -960 239670 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 243054 -960 243166 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 246550 -960 246662 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 250138 -960 250250 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 253634 -960 253746 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 257222 -960 257334 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 260718 -960 260830 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 264214 -960 264326 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137070 -960 137182 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 267802 -960 267914 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 271298 -960 271410 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 274886 -960 274998 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 278382 -960 278494 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 281878 -960 281990 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 285466 -960 285578 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 288962 -960 289074 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 292550 -960 292662 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 296046 -960 296158 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 299542 -960 299654 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 140658 -960 140770 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 303130 -960 303242 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 306626 -960 306738 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 310122 -960 310234 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 313710 -960 313822 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 317206 -960 317318 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 320794 -960 320906 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 324290 -960 324402 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 327786 -960 327898 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 331374 -960 331486 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 334870 -960 334982 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144154 -960 144266 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 338458 -960 338570 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 341954 -960 342066 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 359618 -960 359730 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 363114 -960 363226 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 366702 -960 366814 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 370198 -960 370310 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 147650 -960 147762 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 373786 -960 373898 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 377282 -960 377394 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 380778 -960 380890 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 384366 -960 384478 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 387862 -960 387974 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 391450 -960 391562 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 394946 -960 395058 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 398442 -960 398554 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 402030 -960 402142 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 405526 -960 405638 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151238 -960 151350 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 409114 -960 409226 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 412610 -960 412722 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 416106 -960 416218 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 419694 -960 419806 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 423190 -960 423302 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 426778 -960 426890 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 430274 -960 430386 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 433770 -960 433882 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 437358 -960 437470 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 440854 -960 440966 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 154734 -960 154846 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 444350 -960 444462 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 447938 -960 448050 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 451434 -960 451546 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 455022 -960 455134 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 458518 -960 458630 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 462014 -960 462126 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 465602 -960 465714 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 469098 -960 469210 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 472686 -960 472798 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 476182 -960 476294 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158230 -960 158342 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 127686 -960 127798 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 480874 -960 480986 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 484462 -960 484574 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 487958 -960 488070 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 491454 -960 491566 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 495042 -960 495154 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 498538 -960 498650 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 502126 -960 502238 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 505622 -960 505734 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 509118 -960 509230 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 512706 -960 512818 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163014 -960 163126 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 516202 -960 516314 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 519790 -960 519902 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 523286 -960 523398 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 526782 -960 526894 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 530370 -960 530482 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 533866 -960 533978 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 537454 -960 537566 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 540950 -960 541062 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 544446 -960 544558 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 548034 -960 548146 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 166510 -960 166622 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 551530 -960 551642 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 555118 -960 555230 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 558614 -960 558726 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 562110 -960 562222 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 565698 -960 565810 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 569194 -960 569306 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 572782 -960 572894 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170006 -960 170118 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 173594 -960 173706 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177090 -960 177202 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 180678 -960 180790 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184174 -960 184286 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 187670 -960 187782 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191258 -960 191370 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 194754 -960 194866 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131182 -960 131294 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 198342 -960 198454 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 201838 -960 201950 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 205334 -960 205446 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 208922 -960 209034 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 212418 -960 212530 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216006 -960 216118 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 219502 -960 219614 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 222998 -960 223110 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 226586 -960 226698 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 134770 -960 134882 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 240662 -960 240774 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 244250 -960 244362 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 247746 -960 247858 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 251334 -960 251446 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 254830 -960 254942 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 258326 -960 258438 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 261914 -960 262026 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 265410 -960 265522 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138266 -960 138378 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 268998 -960 269110 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 272494 -960 272606 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 275990 -960 276102 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 279578 -960 279690 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 283074 -960 283186 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 286662 -960 286774 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 290158 -960 290270 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 293654 -960 293766 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 297242 -960 297354 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 300738 -960 300850 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 141762 -960 141874 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 304234 -960 304346 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 307822 -960 307934 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 311318 -960 311430 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 314906 -960 315018 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 318402 -960 318514 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 321898 -960 322010 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 325486 -960 325598 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 328982 -960 329094 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 332570 -960 332682 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 336066 -960 336178 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145350 -960 145462 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 339562 -960 339674 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 343150 -960 343262 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 357226 -960 357338 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 360814 -960 360926 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 364310 -960 364422 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 367898 -960 368010 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 371394 -960 371506 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 148846 -960 148958 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 374890 -960 375002 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 378478 -960 378590 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 381974 -960 382086 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 385562 -960 385674 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 389058 -960 389170 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 392554 -960 392666 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 396142 -960 396254 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 399638 -960 399750 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 403226 -960 403338 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 406722 -960 406834 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152342 -960 152454 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 410218 -960 410330 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 413806 -960 413918 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 417302 -960 417414 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 420890 -960 421002 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 424386 -960 424498 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 427882 -960 427994 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 431470 -960 431582 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 434966 -960 435078 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 438554 -960 438666 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 442050 -960 442162 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 155930 -960 156042 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 445546 -960 445658 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 449134 -960 449246 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 452630 -960 452742 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 456126 -960 456238 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 459714 -960 459826 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 463210 -960 463322 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 466798 -960 466910 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 470294 -960 470406 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 473790 -960 473902 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 477378 -960 477490 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 159426 -960 159538 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 577474 -960 577586 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 578670 -960 578782 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 579774 -960 579886 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 580970 -960 581082 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 73794 561806 254414 562426 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 -1894 74414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 -1894 110414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 -1894 146414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 -1894 182414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 -1894 218414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 -1894 254414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 -1894 290414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 -1894 326414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 -1894 398414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 -1894 434414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 -1894 470414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 -1894 506414 43000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 130308 74414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 130308 110414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 130308 146414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 130308 182414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 130308 218414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 130308 254414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 130308 290414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 130308 326414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 130308 398414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 130308 434414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 130308 470414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 130308 506414 153000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 240308 74414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 240308 110414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 240308 146414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 240308 182414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 240308 218414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 240308 254414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 240308 290414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 240308 326414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 240308 398414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 240308 434414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 240308 470414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 240308 506414 263000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 350308 74414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 350308 110414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 350308 146414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 350308 182414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 350308 218414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 350308 254414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 350308 290414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 350308 326414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 350308 398414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 350308 434414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 350308 470414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 350308 506414 373000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 460308 74414 493000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 460308 110414 493000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 460308 146414 493000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 460308 182414 493000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 460308 218414 493000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 460308 254414 493000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 460308 290414 493000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 460308 326414 533000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 -1894 362414 533000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 460308 398414 533000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 557000 74414 573000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 557000 110414 573000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 557000 146414 573000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 557000 182414 573000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 557000 218414 573000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 557000 254414 573000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 460308 470414 583000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 460308 506414 583000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 640099 74414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 640099 110414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 640099 146414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 640099 182414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 640099 218414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 640099 254414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 557000 290414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 648033 326414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 648033 362414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 648033 398414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 460308 434414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 637000 470414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 637000 506414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 532 nsew power bidirectional
rlabel metal2 s 22990 703520 23102 704960 6 vccd1
port 533 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s 77514 565526 258134 566146 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 77514 -3814 78134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 113514 -3814 114134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 149514 -3814 150134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 185514 -3814 186134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 221514 -3814 222134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 257514 -3814 258134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 293514 -3814 294134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 329514 -3814 330134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 401514 -3814 402134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 437514 -3814 438134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 473514 -3814 474134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 509514 -3814 510134 43000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 77514 130308 78134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 113514 130308 114134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 149514 130308 150134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 185514 130308 186134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 221514 130308 222134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 257514 130308 258134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 293514 130308 294134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 329514 130308 330134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 401514 130308 402134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 437514 130308 438134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 473514 130308 474134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 509514 130308 510134 153000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 77514 240308 78134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 113514 240308 114134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 149514 240308 150134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 185514 240308 186134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 221514 240308 222134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 257514 240308 258134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 293514 240308 294134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 329514 240308 330134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 401514 240308 402134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 437514 240308 438134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 473514 240308 474134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 509514 240308 510134 263000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 77514 350308 78134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 113514 350308 114134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 149514 350308 150134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 185514 350308 186134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 221514 350308 222134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 257514 350308 258134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 293514 350308 294134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 329514 350308 330134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 401514 350308 402134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 437514 350308 438134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 473514 350308 474134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 509514 350308 510134 373000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 77514 460308 78134 493000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 113514 460308 114134 493000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 149514 460308 150134 493000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 185514 460308 186134 493000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 221514 460308 222134 493000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 257514 460308 258134 493000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 293514 460308 294134 493000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 329514 460308 330134 533000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 365514 -3814 366134 533000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 401514 460308 402134 533000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 77514 557000 78134 573000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 113514 557000 114134 573000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 149514 557000 150134 573000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 185514 557000 186134 573000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 221514 557000 222134 573000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 257514 557000 258134 573000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 473514 460308 474134 583000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 509514 460308 510134 583000 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 77514 640099 78134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 113514 640099 114134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 149514 640099 150134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 185514 640099 186134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 221514 640099 222134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 257514 640099 258134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 293514 557000 294134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 329514 648033 330134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 365514 648033 366134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 401514 648033 402134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 437514 460308 438134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 473514 637000 474134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 509514 637000 510134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 534 nsew power bidirectional
rlabel metal2 s 582166 -960 582278 480 8 vccd2
port 535 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s 81234 137246 513854 137866 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s 81234 567366 261854 567986 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 81234 -5734 81854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 117234 -5734 117854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 153234 -5734 153854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 189234 -5734 189854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 225234 -5734 225854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 261234 -5734 261854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 297234 -5734 297854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 333234 -5734 333854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 405234 -5734 405854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 441234 -5734 441854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 477234 -5734 477854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 513234 -5734 513854 43000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 81234 130308 81854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 117234 130308 117854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 153234 130308 153854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 189234 130308 189854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 225234 130308 225854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 261234 130308 261854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 297234 130308 297854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 333234 130308 333854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 405234 130308 405854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 441234 130308 441854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 477234 130308 477854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 513234 130308 513854 153000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 81234 240308 81854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 117234 240308 117854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 153234 240308 153854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 189234 240308 189854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 225234 240308 225854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 261234 240308 261854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 297234 240308 297854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 333234 240308 333854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 405234 240308 405854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 441234 240308 441854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 477234 240308 477854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 513234 240308 513854 263000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 81234 350308 81854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 117234 350308 117854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 153234 350308 153854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 189234 350308 189854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 225234 350308 225854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 261234 350308 261854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 297234 350308 297854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 333234 350308 333854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 405234 350308 405854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 441234 350308 441854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 477234 350308 477854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 513234 350308 513854 373000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 81234 460308 81854 493000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 117234 460308 117854 493000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 153234 460308 153854 493000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 189234 460308 189854 493000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 225234 460308 225854 493000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 261234 460308 261854 493000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 297234 460308 297854 493000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 333234 460308 333854 533000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 369234 -5734 369854 533000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 405234 460308 405854 533000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 81234 557000 81854 573000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 117234 557000 117854 573000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 153234 557000 153854 573000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 189234 557000 189854 573000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 225234 557000 225854 573000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 261234 557000 261854 573000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 477234 460308 477854 583000 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 81234 640099 81854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 117234 640099 117854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 153234 640099 153854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 189234 640099 189854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 225234 640099 225854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 261234 640099 261854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 297234 557000 297854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 333234 648033 333854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 369234 648033 369854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 405234 648033 405854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 441234 460308 441854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 477234 637000 477854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 513234 460308 513854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 536 nsew power bidirectional
rlabel metal3 s 583520 684572 584960 684812 6 vdda1
port 537 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s 84954 140966 517574 141586 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s 84954 248966 517574 249586 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s 84954 356966 517574 357586 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s 84954 571086 265574 571706 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 84954 -7654 85574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 120954 -7654 121574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 156954 -7654 157574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 192954 -7654 193574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 228954 -7654 229574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 264954 -7654 265574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 300954 -7654 301574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 336954 -7654 337574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 408954 -7654 409574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 444954 -7654 445574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 480954 -7654 481574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 516954 -7654 517574 43000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 84954 130308 85574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 120954 130308 121574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 156954 130308 157574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 192954 130308 193574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 228954 130308 229574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 264954 130308 265574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 300954 130308 301574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 336954 130308 337574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 408954 130308 409574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 444954 130308 445574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 480954 130308 481574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 516954 130308 517574 153000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 84954 240308 85574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 120954 240308 121574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 156954 240308 157574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 192954 240308 193574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 228954 240308 229574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 264954 240308 265574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 300954 240308 301574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 336954 240308 337574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 408954 240308 409574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 444954 240308 445574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 480954 240308 481574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 516954 240308 517574 263000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 84954 350308 85574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 120954 350308 121574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 156954 350308 157574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 192954 350308 193574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 228954 350308 229574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 264954 350308 265574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 300954 350308 301574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 336954 350308 337574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 408954 350308 409574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 444954 350308 445574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 480954 350308 481574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 516954 350308 517574 373000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 84954 460308 85574 493000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 120954 460308 121574 493000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 156954 460308 157574 493000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 192954 460308 193574 493000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 228954 460308 229574 493000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 264954 460308 265574 493000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 300954 460308 301574 493000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 336954 460308 337574 533000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 372954 -7654 373574 533000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 408954 460308 409574 533000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 84954 557000 85574 573000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 120954 557000 121574 573000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 156954 557000 157574 573000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 192954 557000 193574 573000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 228954 557000 229574 573000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 264954 557000 265574 573000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 480954 460308 481574 583000 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 84954 640099 85574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 120954 640099 121574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 156954 640099 157574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 192954 640099 193574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 228954 640099 229574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 264954 640099 265574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 300954 557000 301574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 336954 648033 337574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 372954 648033 373574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 408954 648033 409574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 444954 460308 445574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 480954 637000 481574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 516954 460308 517574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 538 nsew power bidirectional
rlabel metal2 s 7626 703520 7738 704960 6 vdda2
port 539 nsew power bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s 63234 477366 279854 477986 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 63234 -5734 63854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 99234 -5734 99854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 135234 -5734 135854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 171234 -5734 171854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 243234 -5734 243854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 279234 -5734 279854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 315234 -5734 315854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 351234 -5734 351854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 387234 -5734 387854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 423234 -5734 423854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 459234 -5734 459854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 495234 -5734 495854 43000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 63234 130308 63854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 99234 130308 99854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 135234 130308 135854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 171234 130308 171854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 243234 130308 243854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 279234 130308 279854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 315234 130308 315854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 351234 130308 351854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 387234 130308 387854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 423234 130308 423854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 459234 130308 459854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 495234 130308 495854 153000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 63234 240308 63854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 99234 240308 99854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 135234 240308 135854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 171234 240308 171854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 243234 240308 243854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 279234 240308 279854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 315234 240308 315854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 351234 240308 351854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 387234 240308 387854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 423234 240308 423854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 459234 240308 459854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 495234 240308 495854 263000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 63234 350308 63854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 99234 350308 99854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 135234 350308 135854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 171234 350308 171854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 243234 350308 243854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 279234 350308 279854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 315234 350308 315854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 351234 350308 351854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 387234 350308 387854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 423234 350308 423854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 459234 350308 459854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 495234 350308 495854 373000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 63234 460308 63854 493000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 99234 460308 99854 493000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 135234 460308 135854 493000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 171234 460308 171854 493000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 207234 -5734 207854 493000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 243234 460308 243854 493000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 279234 460308 279854 493000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 351234 460308 351854 533000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 387234 460308 387854 533000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 423234 460308 423854 533000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 63234 557000 63854 573000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 99234 557000 99854 573000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 171234 557000 171854 573000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 243234 557000 243854 573000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 279234 557000 279854 573000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 459234 460308 459854 583000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 495234 460308 495854 583000 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 63234 640099 63854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 99234 640099 99854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 135234 557000 135854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 171234 640099 171854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 207234 557000 207854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 243234 640099 243854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 279234 640099 279854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 315234 460308 315854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 351234 648033 351854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 387234 648033 387854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 423234 648033 423854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 459234 637000 459854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 495234 637000 495854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 540 nsew ground bidirectional
rlabel metal2 s 583362 -960 583474 480 8 vssa1
port 541 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 66954 -7654 67574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 102954 -7654 103574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 138954 -7654 139574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 174954 -7654 175574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 246954 -7654 247574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 282954 -7654 283574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 318954 -7654 319574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 354954 -7654 355574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 390954 -7654 391574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 426954 -7654 427574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 462954 -7654 463574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 498954 -7654 499574 43000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 66954 130308 67574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 102954 130308 103574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 138954 130308 139574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 174954 130308 175574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 246954 130308 247574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 282954 130308 283574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 318954 130308 319574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 354954 130308 355574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 390954 130308 391574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 426954 130308 427574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 462954 130308 463574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 498954 130308 499574 153000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 66954 240308 67574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 102954 240308 103574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 138954 240308 139574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 174954 240308 175574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 246954 240308 247574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 282954 240308 283574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 318954 240308 319574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 354954 240308 355574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 390954 240308 391574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 426954 240308 427574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 462954 240308 463574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 498954 240308 499574 263000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 66954 350308 67574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 102954 350308 103574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 138954 350308 139574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 174954 350308 175574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 246954 350308 247574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 282954 350308 283574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 318954 350308 319574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 354954 350308 355574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 390954 350308 391574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 426954 350308 427574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 462954 350308 463574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 498954 350308 499574 373000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 66954 460308 67574 493000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 102954 460308 103574 493000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 138954 460308 139574 493000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 174954 460308 175574 493000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 210954 -7654 211574 493000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 246954 460308 247574 493000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 282954 460308 283574 493000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 318954 460308 319574 533000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 354954 460308 355574 533000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 390954 460308 391574 533000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 426954 460308 427574 533000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 66954 557000 67574 573000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 102954 557000 103574 573000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 138954 557000 139574 573000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 174954 557000 175574 573000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 246954 557000 247574 573000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 282954 557000 283574 573000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 462954 460308 463574 583000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 498954 460308 499574 583000 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 66954 640099 67574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 102954 640099 103574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 138954 640099 139574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 174954 640099 175574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 210954 557000 211574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 246954 640099 247574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 282954 640099 283574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 318954 648033 319574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 354954 648033 355574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 390954 648033 391574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 426954 648033 427574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 462954 637000 463574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 498954 637000 499574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 542 nsew ground bidirectional
rlabel metal3 s 583520 697356 584960 697596 6 vssa2
port 543 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s 91794 145926 488414 146546 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s 91794 253926 488414 254546 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s 91794 361926 488414 362546 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 91794 -1894 92414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 127794 -1894 128414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 163794 -1894 164414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 235794 -1894 236414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 271794 -1894 272414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 307794 -1894 308414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 343794 -1894 344414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 379794 -1894 380414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 415794 -1894 416414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 451794 -1894 452414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 487794 -1894 488414 43000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 91794 130308 92414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 127794 130308 128414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 163794 130308 164414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 235794 130308 236414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 271794 130308 272414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 307794 130308 308414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 343794 130308 344414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 379794 130308 380414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 415794 130308 416414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 451794 130308 452414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 487794 130308 488414 153000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 91794 240308 92414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 127794 240308 128414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 163794 240308 164414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 235794 240308 236414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 271794 240308 272414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 307794 240308 308414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 343794 240308 344414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 379794 240308 380414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 415794 240308 416414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 451794 240308 452414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 487794 240308 488414 263000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 91794 350308 92414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 127794 350308 128414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 163794 350308 164414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 235794 350308 236414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 271794 350308 272414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 307794 350308 308414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 343794 350308 344414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 379794 350308 380414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 415794 350308 416414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 451794 350308 452414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 487794 350308 488414 373000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 91794 460308 92414 493000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 127794 460308 128414 493000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 163794 460308 164414 493000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 199794 -1894 200414 493000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 235794 460308 236414 493000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 271794 460308 272414 493000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 343794 460308 344414 533000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 379794 460308 380414 533000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 415794 460308 416414 533000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 91794 557000 92414 573000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 163794 557000 164414 573000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 199794 557000 200414 573000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 235794 557000 236414 573000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 271794 557000 272414 573000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 487794 460308 488414 583000 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 91794 640099 92414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 127794 557000 128414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 163794 640099 164414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 199794 640099 200414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 235794 640099 236414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 271794 640099 272414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 307794 460308 308414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 343794 648033 344414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 379794 648033 380414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 415794 648033 416414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 451794 460308 452414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 487794 637000 488414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 544 nsew ground bidirectional
rlabel metal3 s -960 18716 480 18956 4 vssd1
port 545 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s 59514 365646 492134 366266 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s 59514 475526 276134 476146 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 546 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 59514 -3814 60134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 95514 -3814 96134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 131514 -3814 132134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 167514 -3814 168134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 239514 -3814 240134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 275514 -3814 276134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 311514 -3814 312134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 347514 -3814 348134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 383514 -3814 384134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 419514 -3814 420134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 455514 -3814 456134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 491514 -3814 492134 43000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 59514 130308 60134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 95514 130308 96134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 131514 130308 132134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 167514 130308 168134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 239514 130308 240134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 275514 130308 276134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 311514 130308 312134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 347514 130308 348134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 383514 130308 384134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 419514 130308 420134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 455514 130308 456134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 491514 130308 492134 153000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 59514 240308 60134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 95514 240308 96134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 131514 240308 132134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 167514 240308 168134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 239514 240308 240134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 275514 240308 276134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 311514 240308 312134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 347514 240308 348134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 383514 240308 384134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 419514 240308 420134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 455514 240308 456134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 491514 240308 492134 263000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 59514 350308 60134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 95514 350308 96134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 131514 350308 132134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 167514 350308 168134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 239514 350308 240134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 275514 350308 276134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 311514 350308 312134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 347514 350308 348134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 383514 350308 384134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 419514 350308 420134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 455514 350308 456134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 491514 350308 492134 373000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 59514 460308 60134 493000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 95514 460308 96134 493000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 131514 460308 132134 493000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 167514 460308 168134 493000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 203514 -3814 204134 493000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 239514 460308 240134 493000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 275514 460308 276134 493000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 347514 460308 348134 533000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 383514 460308 384134 533000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 419514 460308 420134 533000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 59514 557000 60134 573000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 95514 557000 96134 573000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 167514 557000 168134 573000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 239514 557000 240134 573000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 275514 557000 276134 573000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 491514 460308 492134 583000 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 59514 640099 60134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 95514 640099 96134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 131514 557000 132134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 167514 640099 168134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 203514 557000 204134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 239514 640099 240134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 275514 640099 276134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 311514 460308 312134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 347514 648033 348134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 383514 648033 384134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 419514 648033 420134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 455514 460308 456134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 491514 637000 492134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 546 nsew ground bidirectional
rlabel metal3 s -960 6204 480 6444 4 vssd2
port 547 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 548 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 549 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 550 nsew signal output
rlabel metal2 s 7534 -960 7646 480 8 wbs_adr_i[0]
port 551 nsew signal input
rlabel metal2 s 47554 -960 47666 480 8 wbs_adr_i[10]
port 552 nsew signal input
rlabel metal2 s 51142 -960 51254 480 8 wbs_adr_i[11]
port 553 nsew signal input
rlabel metal2 s 54638 -960 54750 480 8 wbs_adr_i[12]
port 554 nsew signal input
rlabel metal2 s 58226 -960 58338 480 8 wbs_adr_i[13]
port 555 nsew signal input
rlabel metal2 s 61722 -960 61834 480 8 wbs_adr_i[14]
port 556 nsew signal input
rlabel metal2 s 65218 -960 65330 480 8 wbs_adr_i[15]
port 557 nsew signal input
rlabel metal2 s 68806 -960 68918 480 8 wbs_adr_i[16]
port 558 nsew signal input
rlabel metal2 s 72302 -960 72414 480 8 wbs_adr_i[17]
port 559 nsew signal input
rlabel metal2 s 75890 -960 76002 480 8 wbs_adr_i[18]
port 560 nsew signal input
rlabel metal2 s 79386 -960 79498 480 8 wbs_adr_i[19]
port 561 nsew signal input
rlabel metal2 s 12226 -960 12338 480 8 wbs_adr_i[1]
port 562 nsew signal input
rlabel metal2 s 82882 -960 82994 480 8 wbs_adr_i[20]
port 563 nsew signal input
rlabel metal2 s 86470 -960 86582 480 8 wbs_adr_i[21]
port 564 nsew signal input
rlabel metal2 s 89966 -960 90078 480 8 wbs_adr_i[22]
port 565 nsew signal input
rlabel metal2 s 93554 -960 93666 480 8 wbs_adr_i[23]
port 566 nsew signal input
rlabel metal2 s 97050 -960 97162 480 8 wbs_adr_i[24]
port 567 nsew signal input
rlabel metal2 s 100546 -960 100658 480 8 wbs_adr_i[25]
port 568 nsew signal input
rlabel metal2 s 104134 -960 104246 480 8 wbs_adr_i[26]
port 569 nsew signal input
rlabel metal2 s 107630 -960 107742 480 8 wbs_adr_i[27]
port 570 nsew signal input
rlabel metal2 s 111218 -960 111330 480 8 wbs_adr_i[28]
port 571 nsew signal input
rlabel metal2 s 114714 -960 114826 480 8 wbs_adr_i[29]
port 572 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 573 nsew signal input
rlabel metal2 s 118210 -960 118322 480 8 wbs_adr_i[30]
port 574 nsew signal input
rlabel metal2 s 121798 -960 121910 480 8 wbs_adr_i[31]
port 575 nsew signal input
rlabel metal2 s 21702 -960 21814 480 8 wbs_adr_i[3]
port 576 nsew signal input
rlabel metal2 s 26394 -960 26506 480 8 wbs_adr_i[4]
port 577 nsew signal input
rlabel metal2 s 29890 -960 30002 480 8 wbs_adr_i[5]
port 578 nsew signal input
rlabel metal2 s 33478 -960 33590 480 8 wbs_adr_i[6]
port 579 nsew signal input
rlabel metal2 s 36974 -960 37086 480 8 wbs_adr_i[7]
port 580 nsew signal input
rlabel metal2 s 40562 -960 40674 480 8 wbs_adr_i[8]
port 581 nsew signal input
rlabel metal2 s 44058 -960 44170 480 8 wbs_adr_i[9]
port 582 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 583 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 584 nsew signal input
rlabel metal2 s 48750 -960 48862 480 8 wbs_dat_i[10]
port 585 nsew signal input
rlabel metal2 s 52338 -960 52450 480 8 wbs_dat_i[11]
port 586 nsew signal input
rlabel metal2 s 55834 -960 55946 480 8 wbs_dat_i[12]
port 587 nsew signal input
rlabel metal2 s 59330 -960 59442 480 8 wbs_dat_i[13]
port 588 nsew signal input
rlabel metal2 s 62918 -960 63030 480 8 wbs_dat_i[14]
port 589 nsew signal input
rlabel metal2 s 66414 -960 66526 480 8 wbs_dat_i[15]
port 590 nsew signal input
rlabel metal2 s 70002 -960 70114 480 8 wbs_dat_i[16]
port 591 nsew signal input
rlabel metal2 s 73498 -960 73610 480 8 wbs_dat_i[17]
port 592 nsew signal input
rlabel metal2 s 76994 -960 77106 480 8 wbs_dat_i[18]
port 593 nsew signal input
rlabel metal2 s 80582 -960 80694 480 8 wbs_dat_i[19]
port 594 nsew signal input
rlabel metal2 s 13422 -960 13534 480 8 wbs_dat_i[1]
port 595 nsew signal input
rlabel metal2 s 84078 -960 84190 480 8 wbs_dat_i[20]
port 596 nsew signal input
rlabel metal2 s 87666 -960 87778 480 8 wbs_dat_i[21]
port 597 nsew signal input
rlabel metal2 s 91162 -960 91274 480 8 wbs_dat_i[22]
port 598 nsew signal input
rlabel metal2 s 94658 -960 94770 480 8 wbs_dat_i[23]
port 599 nsew signal input
rlabel metal2 s 98246 -960 98358 480 8 wbs_dat_i[24]
port 600 nsew signal input
rlabel metal2 s 101742 -960 101854 480 8 wbs_dat_i[25]
port 601 nsew signal input
rlabel metal2 s 105330 -960 105442 480 8 wbs_dat_i[26]
port 602 nsew signal input
rlabel metal2 s 108826 -960 108938 480 8 wbs_dat_i[27]
port 603 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_dat_i[28]
port 604 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_dat_i[29]
port 605 nsew signal input
rlabel metal2 s 18114 -960 18226 480 8 wbs_dat_i[2]
port 606 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_dat_i[30]
port 607 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_dat_i[31]
port 608 nsew signal input
rlabel metal2 s 22898 -960 23010 480 8 wbs_dat_i[3]
port 609 nsew signal input
rlabel metal2 s 27590 -960 27702 480 8 wbs_dat_i[4]
port 610 nsew signal input
rlabel metal2 s 31086 -960 31198 480 8 wbs_dat_i[5]
port 611 nsew signal input
rlabel metal2 s 34674 -960 34786 480 8 wbs_dat_i[6]
port 612 nsew signal input
rlabel metal2 s 38170 -960 38282 480 8 wbs_dat_i[7]
port 613 nsew signal input
rlabel metal2 s 41666 -960 41778 480 8 wbs_dat_i[8]
port 614 nsew signal input
rlabel metal2 s 45254 -960 45366 480 8 wbs_dat_i[9]
port 615 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 616 nsew signal output
rlabel metal2 s 49946 -960 50058 480 8 wbs_dat_o[10]
port 617 nsew signal output
rlabel metal2 s 53442 -960 53554 480 8 wbs_dat_o[11]
port 618 nsew signal output
rlabel metal2 s 57030 -960 57142 480 8 wbs_dat_o[12]
port 619 nsew signal output
rlabel metal2 s 60526 -960 60638 480 8 wbs_dat_o[13]
port 620 nsew signal output
rlabel metal2 s 64114 -960 64226 480 8 wbs_dat_o[14]
port 621 nsew signal output
rlabel metal2 s 67610 -960 67722 480 8 wbs_dat_o[15]
port 622 nsew signal output
rlabel metal2 s 71106 -960 71218 480 8 wbs_dat_o[16]
port 623 nsew signal output
rlabel metal2 s 74694 -960 74806 480 8 wbs_dat_o[17]
port 624 nsew signal output
rlabel metal2 s 78190 -960 78302 480 8 wbs_dat_o[18]
port 625 nsew signal output
rlabel metal2 s 81778 -960 81890 480 8 wbs_dat_o[19]
port 626 nsew signal output
rlabel metal2 s 14618 -960 14730 480 8 wbs_dat_o[1]
port 627 nsew signal output
rlabel metal2 s 85274 -960 85386 480 8 wbs_dat_o[20]
port 628 nsew signal output
rlabel metal2 s 88770 -960 88882 480 8 wbs_dat_o[21]
port 629 nsew signal output
rlabel metal2 s 92358 -960 92470 480 8 wbs_dat_o[22]
port 630 nsew signal output
rlabel metal2 s 95854 -960 95966 480 8 wbs_dat_o[23]
port 631 nsew signal output
rlabel metal2 s 99442 -960 99554 480 8 wbs_dat_o[24]
port 632 nsew signal output
rlabel metal2 s 102938 -960 103050 480 8 wbs_dat_o[25]
port 633 nsew signal output
rlabel metal2 s 106434 -960 106546 480 8 wbs_dat_o[26]
port 634 nsew signal output
rlabel metal2 s 110022 -960 110134 480 8 wbs_dat_o[27]
port 635 nsew signal output
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_o[28]
port 636 nsew signal output
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_o[29]
port 637 nsew signal output
rlabel metal2 s 19310 -960 19422 480 8 wbs_dat_o[2]
port 638 nsew signal output
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_o[30]
port 639 nsew signal output
rlabel metal2 s 124098 -960 124210 480 8 wbs_dat_o[31]
port 640 nsew signal output
rlabel metal2 s 24002 -960 24114 480 8 wbs_dat_o[3]
port 641 nsew signal output
rlabel metal2 s 28786 -960 28898 480 8 wbs_dat_o[4]
port 642 nsew signal output
rlabel metal2 s 32282 -960 32394 480 8 wbs_dat_o[5]
port 643 nsew signal output
rlabel metal2 s 35778 -960 35890 480 8 wbs_dat_o[6]
port 644 nsew signal output
rlabel metal2 s 39366 -960 39478 480 8 wbs_dat_o[7]
port 645 nsew signal output
rlabel metal2 s 42862 -960 42974 480 8 wbs_dat_o[8]
port 646 nsew signal output
rlabel metal2 s 46450 -960 46562 480 8 wbs_dat_o[9]
port 647 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 648 nsew signal input
rlabel metal2 s 15814 -960 15926 480 8 wbs_sel_i[1]
port 649 nsew signal input
rlabel metal2 s 20506 -960 20618 480 8 wbs_sel_i[2]
port 650 nsew signal input
rlabel metal2 s 25198 -960 25310 480 8 wbs_sel_i[3]
port 651 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 652 nsew signal input
rlabel metal2 s 6338 -960 6450 480 8 wbs_we_i
port 653 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 97600142
string GDS_FILE /home/burak/asic_tools/caravel_vscpu3x/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 94134178
<< end >>

