magic
tech sky130A
magscale 1 2
timestamp 1655395605
<< metal1 >>
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 305638 700380 305644 700392
rect 235224 700352 305644 700380
rect 235224 700340 235230 700352
rect 305638 700340 305644 700352
rect 305696 700340 305702 700392
rect 57882 700272 57888 700324
rect 57940 700312 57946 700324
rect 543458 700312 543464 700324
rect 57940 700284 543464 700312
rect 57940 700272 57946 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 137922 683136 137928 683188
rect 137980 683176 137986 683188
rect 580166 683176 580172 683188
rect 137980 683148 580172 683176
rect 137980 683136 137986 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 169754 640976 169760 641028
rect 169812 641016 169818 641028
rect 430942 641016 430948 641028
rect 169812 640988 430948 641016
rect 169812 640976 169818 640988
rect 430942 640976 430948 640988
rect 431000 640976 431006 641028
rect 3418 639548 3424 639600
rect 3476 639588 3482 639600
rect 317046 639588 317052 639600
rect 3476 639560 317052 639588
rect 3476 639548 3482 639560
rect 317046 639548 317052 639560
rect 317104 639548 317110 639600
rect 104894 638188 104900 638240
rect 104952 638228 104958 638240
rect 429286 638228 429292 638240
rect 104952 638200 429292 638228
rect 104952 638188 104958 638200
rect 429286 638188 429292 638200
rect 429344 638188 429350 638240
rect 299474 636828 299480 636880
rect 299532 636868 299538 636880
rect 401134 636868 401140 636880
rect 299532 636840 401140 636868
rect 299532 636828 299538 636840
rect 401134 636828 401140 636840
rect 401192 636828 401198 636880
rect 364334 635468 364340 635520
rect 364392 635508 364398 635520
rect 423674 635508 423680 635520
rect 364392 635480 423680 635508
rect 364392 635468 364398 635480
rect 423674 635468 423680 635480
rect 423732 635468 423738 635520
rect 316954 634924 316960 634976
rect 317012 634964 317018 634976
rect 430574 634964 430580 634976
rect 317012 634936 430580 634964
rect 317012 634924 317018 634936
rect 430574 634924 430580 634936
rect 430632 634924 430638 634976
rect 316862 634856 316868 634908
rect 316920 634896 316926 634908
rect 430850 634896 430856 634908
rect 316920 634868 430856 634896
rect 316920 634856 316926 634868
rect 430850 634856 430856 634868
rect 430908 634856 430914 634908
rect 291194 634788 291200 634840
rect 291252 634828 291258 634840
rect 457438 634828 457444 634840
rect 291252 634800 457444 634828
rect 291252 634788 291258 634800
rect 457438 634788 457444 634800
rect 457496 634788 457502 634840
rect 318794 634040 318800 634092
rect 318852 634080 318858 634092
rect 494054 634080 494060 634092
rect 318852 634052 494060 634080
rect 318852 634040 318858 634052
rect 494054 634040 494060 634052
rect 494112 634040 494118 634092
rect 280982 633632 280988 633684
rect 281040 633672 281046 633684
rect 383102 633672 383108 633684
rect 281040 633644 383108 633672
rect 281040 633632 281046 633644
rect 383102 633632 383108 633644
rect 383160 633632 383166 633684
rect 281074 633564 281080 633616
rect 281132 633604 281138 633616
rect 430758 633604 430764 633616
rect 281132 633576 430764 633604
rect 281132 633564 281138 633576
rect 430758 633564 430764 633576
rect 430816 633564 430822 633616
rect 289814 633496 289820 633548
rect 289872 633536 289878 633548
rect 489914 633536 489920 633548
rect 289872 633508 489920 633536
rect 289872 633496 289878 633508
rect 489914 633496 489920 633508
rect 489972 633496 489978 633548
rect 288434 633428 288440 633480
rect 288492 633468 288498 633480
rect 511994 633468 512000 633480
rect 288492 633440 512000 633468
rect 288492 633428 288498 633440
rect 511994 633428 512000 633440
rect 512052 633428 512058 633480
rect 313918 632952 313924 633004
rect 313976 632992 313982 633004
rect 337378 632992 337384 633004
rect 313976 632964 337384 632992
rect 313976 632952 313982 632964
rect 337378 632952 337384 632964
rect 337436 632952 337442 633004
rect 309778 632884 309784 632936
rect 309836 632924 309842 632936
rect 332870 632924 332876 632936
rect 309836 632896 332876 632924
rect 309836 632884 309842 632896
rect 332870 632884 332876 632896
rect 332928 632884 332934 632936
rect 295978 632816 295984 632868
rect 296036 632856 296042 632868
rect 378594 632856 378600 632868
rect 296036 632828 378600 632856
rect 296036 632816 296042 632828
rect 378594 632816 378600 632828
rect 378652 632816 378658 632868
rect 291286 632748 291292 632800
rect 291344 632788 291350 632800
rect 432598 632788 432604 632800
rect 291344 632760 432604 632788
rect 291344 632748 291350 632760
rect 432598 632748 432604 632760
rect 432656 632748 432662 632800
rect 319530 632680 319536 632732
rect 319588 632720 319594 632732
rect 355410 632720 355416 632732
rect 319588 632692 355416 632720
rect 319588 632680 319594 632692
rect 355410 632680 355416 632692
rect 355468 632680 355474 632732
rect 311158 632612 311164 632664
rect 311216 632652 311222 632664
rect 350902 632652 350908 632664
rect 311216 632624 350908 632652
rect 311216 632612 311222 632624
rect 350902 632612 350908 632624
rect 350960 632612 350966 632664
rect 319714 632544 319720 632596
rect 319772 632584 319778 632596
rect 364426 632584 364432 632596
rect 319772 632556 364432 632584
rect 319772 632544 319778 632556
rect 364426 632544 364432 632556
rect 364484 632544 364490 632596
rect 312538 632476 312544 632528
rect 312596 632516 312602 632528
rect 359918 632516 359924 632528
rect 312596 632488 359924 632516
rect 312596 632476 312602 632488
rect 359918 632476 359924 632488
rect 359976 632476 359982 632528
rect 319806 632408 319812 632460
rect 319864 632448 319870 632460
rect 373442 632448 373448 632460
rect 319864 632420 373448 632448
rect 319864 632408 319870 632420
rect 373442 632408 373448 632420
rect 373500 632408 373506 632460
rect 316770 632340 316776 632392
rect 316828 632380 316834 632392
rect 387610 632380 387616 632392
rect 316828 632352 387616 632380
rect 316828 632340 316834 632352
rect 387610 632340 387616 632352
rect 387668 632340 387674 632392
rect 316678 632272 316684 632324
rect 316736 632312 316742 632324
rect 396626 632312 396632 632324
rect 316736 632284 396632 632312
rect 316736 632272 316742 632284
rect 396626 632272 396632 632284
rect 396684 632272 396690 632324
rect 320818 632204 320824 632256
rect 320876 632244 320882 632256
rect 341886 632244 341892 632256
rect 320876 632216 341892 632244
rect 320876 632204 320882 632216
rect 341886 632204 341892 632216
rect 341944 632204 341950 632256
rect 318242 632136 318248 632188
rect 318300 632176 318306 632188
rect 428182 632176 428188 632188
rect 318300 632148 428188 632176
rect 318300 632136 318306 632148
rect 428182 632136 428188 632148
rect 428240 632136 428246 632188
rect 319898 632068 319904 632120
rect 319956 632108 319962 632120
rect 323854 632108 323860 632120
rect 319956 632080 323860 632108
rect 319956 632068 319962 632080
rect 323854 632068 323860 632080
rect 323912 632068 323918 632120
rect 284938 631320 284944 631372
rect 284996 631360 285002 631372
rect 368934 631360 368940 631372
rect 284996 631332 368940 631360
rect 284996 631320 285002 631332
rect 368934 631320 368940 631332
rect 368992 631320 368998 631372
rect 318058 631252 318064 631304
rect 318116 631292 318122 631304
rect 430666 631292 430672 631304
rect 318116 631264 430672 631292
rect 318116 631252 318122 631264
rect 430666 631252 430672 631264
rect 430724 631252 430730 631304
rect 298094 631184 298100 631236
rect 298152 631224 298158 631236
rect 429838 631224 429844 631236
rect 298152 631196 429844 631224
rect 298152 631184 298158 631196
rect 429838 631184 429844 631196
rect 429896 631184 429902 631236
rect 296806 631116 296812 631168
rect 296864 631156 296870 631168
rect 435358 631156 435364 631168
rect 296864 631128 435364 631156
rect 296864 631116 296870 631128
rect 435358 631116 435364 631128
rect 435416 631116 435422 631168
rect 293954 631048 293960 631100
rect 294012 631088 294018 631100
rect 432690 631088 432696 631100
rect 294012 631060 432696 631088
rect 294012 631048 294018 631060
rect 432690 631048 432696 631060
rect 432748 631048 432754 631100
rect 288526 630980 288532 631032
rect 288584 631020 288590 631032
rect 428458 631020 428464 631032
rect 288584 630992 428464 631020
rect 288584 630980 288590 630992
rect 428458 630980 428464 630992
rect 428516 630980 428522 631032
rect 319438 630912 319444 630964
rect 319496 630952 319502 630964
rect 466730 630952 466736 630964
rect 319496 630924 466736 630952
rect 319496 630912 319502 630924
rect 466730 630912 466736 630924
rect 466788 630912 466794 630964
rect 296714 630844 296720 630896
rect 296772 630884 296778 630896
rect 510614 630884 510620 630896
rect 296772 630856 510620 630884
rect 296772 630844 296778 630856
rect 510614 630844 510620 630856
rect 510672 630844 510678 630896
rect 319070 630776 319076 630828
rect 319128 630816 319134 630828
rect 580166 630816 580172 630828
rect 319128 630788 580172 630816
rect 319128 630776 319134 630788
rect 580166 630776 580172 630788
rect 580224 630776 580230 630828
rect 18598 630708 18604 630760
rect 18656 630748 18662 630760
rect 409874 630748 409880 630760
rect 18656 630720 409880 630748
rect 18656 630708 18662 630720
rect 409874 630708 409880 630720
rect 409932 630708 409938 630760
rect 218698 630640 218704 630692
rect 218756 630680 218762 630692
rect 414382 630680 414388 630692
rect 218756 630652 414388 630680
rect 218756 630640 218762 630652
rect 414382 630640 414388 630652
rect 414440 630640 414446 630692
rect 320818 630476 320824 630488
rect 316006 630448 320824 630476
rect 280706 629960 280712 630012
rect 280764 630000 280770 630012
rect 316006 630000 316034 630448
rect 320818 630436 320824 630448
rect 320876 630436 320882 630488
rect 280764 629972 316034 630000
rect 280764 629960 280770 629972
rect 217778 629892 217784 629944
rect 217836 629932 217842 629944
rect 319070 629932 319076 629944
rect 217836 629904 319076 629932
rect 217836 629892 217842 629904
rect 319070 629892 319076 629904
rect 319128 629892 319134 629944
rect 314010 629280 314016 629332
rect 314068 629320 314074 629332
rect 317782 629320 317788 629332
rect 314068 629292 317788 629320
rect 314068 629280 314074 629292
rect 317782 629280 317788 629292
rect 317840 629280 317846 629332
rect 214006 625744 214012 625796
rect 214064 625784 214070 625796
rect 225414 625784 225420 625796
rect 214064 625756 225420 625784
rect 214064 625744 214070 625756
rect 225414 625744 225420 625756
rect 225472 625744 225478 625796
rect 100570 625676 100576 625728
rect 100628 625716 100634 625728
rect 124306 625716 124312 625728
rect 100628 625688 124312 625716
rect 100628 625676 100634 625688
rect 124306 625676 124312 625688
rect 124364 625676 124370 625728
rect 137830 625676 137836 625728
rect 137888 625716 137894 625728
rect 186498 625716 186504 625728
rect 137888 625688 186504 625716
rect 137888 625676 137894 625688
rect 186498 625676 186504 625688
rect 186556 625676 186562 625728
rect 206462 625676 206468 625728
rect 206520 625716 206526 625728
rect 231302 625716 231308 625728
rect 206520 625688 231308 625716
rect 206520 625676 206526 625688
rect 231302 625676 231308 625688
rect 231360 625676 231366 625728
rect 112162 625608 112168 625660
rect 112220 625648 112226 625660
rect 122834 625648 122840 625660
rect 112220 625620 122840 625648
rect 112220 625608 112226 625620
rect 122834 625608 122840 625620
rect 122892 625608 122898 625660
rect 135162 625608 135168 625660
rect 135220 625648 135226 625660
rect 160278 625648 160284 625660
rect 135220 625620 160284 625648
rect 135220 625608 135226 625620
rect 160278 625608 160284 625620
rect 160336 625608 160342 625660
rect 212534 625608 212540 625660
rect 212592 625648 212598 625660
rect 271874 625648 271880 625660
rect 212592 625620 271880 625648
rect 212592 625608 212598 625620
rect 271874 625608 271880 625620
rect 271932 625608 271938 625660
rect 94774 625540 94780 625592
rect 94832 625580 94838 625592
rect 122282 625580 122288 625592
rect 94832 625552 122288 625580
rect 94832 625540 94838 625552
rect 122282 625540 122288 625552
rect 122340 625540 122346 625592
rect 136450 625540 136456 625592
rect 136508 625580 136514 625592
rect 162854 625580 162860 625592
rect 136508 625552 162860 625580
rect 136508 625540 136514 625552
rect 162854 625540 162860 625552
rect 162912 625540 162918 625592
rect 217870 625540 217876 625592
rect 217928 625580 217934 625592
rect 242894 625580 242900 625592
rect 217928 625552 242900 625580
rect 217928 625540 217934 625552
rect 242894 625540 242900 625552
rect 242952 625540 242958 625592
rect 83182 625472 83188 625524
rect 83240 625512 83246 625524
rect 124398 625512 124404 625524
rect 83240 625484 124404 625512
rect 83240 625472 83246 625484
rect 124398 625472 124404 625484
rect 124456 625472 124462 625524
rect 139210 625472 139216 625524
rect 139268 625512 139274 625524
rect 166166 625512 166172 625524
rect 139268 625484 166172 625512
rect 139268 625472 139274 625484
rect 166166 625472 166172 625484
rect 166224 625472 166230 625524
rect 218882 625472 218888 625524
rect 218940 625512 218946 625524
rect 251910 625512 251916 625524
rect 218940 625484 251916 625512
rect 218940 625472 218946 625484
rect 251910 625472 251916 625484
rect 251968 625472 251974 625524
rect 109586 625404 109592 625456
rect 109644 625444 109650 625456
rect 120902 625444 120908 625456
rect 109644 625416 120908 625444
rect 109644 625404 109650 625416
rect 120902 625404 120908 625416
rect 120960 625404 120966 625456
rect 139118 625404 139124 625456
rect 139176 625444 139182 625456
rect 174446 625444 174452 625456
rect 139176 625416 174452 625444
rect 139176 625404 139182 625416
rect 174446 625404 174452 625416
rect 174504 625404 174510 625456
rect 218790 625404 218796 625456
rect 218848 625444 218854 625456
rect 263594 625444 263600 625456
rect 218848 625416 263600 625444
rect 218848 625404 218854 625416
rect 263594 625404 263600 625416
rect 263652 625404 263658 625456
rect 103790 625336 103796 625388
rect 103848 625376 103854 625388
rect 121638 625376 121644 625388
rect 103848 625348 121644 625376
rect 103848 625336 103854 625348
rect 121638 625336 121644 625348
rect 121696 625336 121702 625388
rect 137738 625336 137744 625388
rect 137796 625376 137802 625388
rect 180334 625376 180340 625388
rect 137796 625348 180340 625376
rect 137796 625336 137802 625348
rect 180334 625336 180340 625348
rect 180392 625336 180398 625388
rect 189994 625336 190000 625388
rect 190052 625376 190058 625388
rect 204530 625376 204536 625388
rect 190052 625348 204536 625376
rect 190052 625336 190058 625348
rect 204530 625336 204536 625348
rect 204588 625336 204594 625388
rect 209774 625336 209780 625388
rect 209832 625376 209838 625388
rect 260190 625376 260196 625388
rect 209832 625348 260196 625376
rect 209832 625336 209838 625348
rect 260190 625336 260196 625348
rect 260248 625336 260254 625388
rect 54846 625268 54852 625320
rect 54904 625308 54910 625320
rect 88978 625308 88984 625320
rect 54904 625280 88984 625308
rect 54904 625268 54910 625280
rect 88978 625268 88984 625280
rect 89036 625268 89042 625320
rect 124214 625268 124220 625320
rect 124272 625308 124278 625320
rect 171870 625308 171876 625320
rect 124272 625280 171876 625308
rect 124272 625268 124278 625280
rect 171870 625268 171876 625280
rect 171928 625268 171934 625320
rect 213914 625268 213920 625320
rect 213972 625308 213978 625320
rect 269206 625308 269212 625320
rect 213972 625280 269212 625308
rect 213972 625268 213978 625280
rect 269206 625268 269212 625280
rect 269264 625268 269270 625320
rect 55122 625200 55128 625252
rect 55180 625240 55186 625252
rect 92198 625240 92204 625252
rect 55180 625212 92204 625240
rect 55180 625200 55186 625212
rect 92198 625200 92204 625212
rect 92256 625200 92262 625252
rect 115382 625200 115388 625252
rect 115440 625240 115446 625252
rect 124674 625240 124680 625252
rect 115440 625212 124680 625240
rect 115440 625200 115446 625212
rect 124674 625200 124680 625212
rect 124732 625200 124738 625252
rect 135254 625200 135260 625252
rect 135312 625240 135318 625252
rect 183646 625240 183652 625252
rect 135312 625212 183652 625240
rect 135312 625200 135318 625212
rect 183646 625200 183652 625212
rect 183704 625200 183710 625252
rect 192570 625200 192576 625252
rect 192628 625240 192634 625252
rect 204438 625240 204444 625252
rect 192628 625212 204444 625240
rect 192628 625200 192634 625212
rect 204438 625200 204444 625212
rect 204496 625200 204502 625252
rect 219342 625200 219348 625252
rect 219400 625240 219406 625252
rect 275094 625240 275100 625252
rect 219400 625212 275100 625240
rect 219400 625200 219406 625212
rect 275094 625200 275100 625212
rect 275152 625200 275158 625252
rect 56502 625132 56508 625184
rect 56560 625172 56566 625184
rect 77386 625172 77392 625184
rect 56560 625144 77392 625172
rect 56560 625132 56566 625144
rect 77386 625132 77392 625144
rect 77444 625132 77450 625184
rect 133874 625132 133880 625184
rect 133932 625172 133938 625184
rect 133932 625144 139808 625172
rect 133932 625132 133938 625144
rect 139780 625104 139808 625144
rect 139854 625132 139860 625184
rect 139912 625172 139918 625184
rect 157518 625172 157524 625184
rect 139912 625144 157524 625172
rect 139912 625132 139918 625144
rect 157518 625132 157524 625144
rect 157576 625132 157582 625184
rect 195698 625132 195704 625184
rect 195756 625172 195762 625184
rect 201678 625172 201684 625184
rect 195756 625144 201684 625172
rect 195756 625132 195762 625144
rect 201678 625132 201684 625144
rect 201736 625132 201742 625184
rect 140130 625104 140136 625116
rect 139780 625076 140136 625104
rect 140130 625064 140136 625076
rect 140188 625064 140194 625116
rect 215294 624044 215300 624096
rect 215352 624084 215358 624096
rect 234614 624084 234620 624096
rect 215352 624056 234620 624084
rect 215352 624044 215358 624056
rect 234614 624044 234620 624056
rect 234672 624044 234678 624096
rect 219618 623976 219624 624028
rect 219676 624016 219682 624028
rect 246022 624016 246028 624028
rect 219676 623988 246028 624016
rect 219676 623976 219682 623988
rect 246022 623976 246028 623988
rect 246080 623976 246086 624028
rect 59354 623908 59360 623960
rect 59412 623948 59418 623960
rect 97994 623948 98000 623960
rect 59412 623920 98000 623948
rect 59412 623908 59418 623920
rect 97994 623908 98000 623920
rect 98052 623908 98058 623960
rect 210418 623908 210424 623960
rect 210476 623948 210482 623960
rect 237558 623948 237564 623960
rect 210476 623920 237564 623948
rect 210476 623908 210482 623920
rect 237558 623908 237564 623920
rect 237616 623908 237622 623960
rect 57790 623840 57796 623892
rect 57848 623880 57854 623892
rect 80606 623880 80612 623892
rect 57848 623852 80612 623880
rect 57848 623840 57854 623852
rect 80606 623840 80612 623852
rect 80664 623840 80670 623892
rect 86402 623840 86408 623892
rect 86460 623880 86466 623892
rect 124582 623880 124588 623892
rect 86460 623852 124588 623880
rect 86460 623840 86466 623852
rect 124582 623840 124588 623852
rect 124640 623840 124646 623892
rect 133138 623840 133144 623892
rect 133196 623880 133202 623892
rect 151262 623880 151268 623892
rect 133196 623852 151268 623880
rect 133196 623840 133202 623852
rect 151262 623840 151268 623852
rect 151320 623840 151326 623892
rect 206278 623840 206284 623892
rect 206336 623880 206342 623892
rect 254486 623880 254492 623892
rect 206336 623852 254492 623880
rect 206336 623840 206342 623852
rect 254486 623840 254492 623852
rect 254544 623840 254550 623892
rect 69014 623772 69020 623824
rect 69072 623812 69078 623824
rect 124490 623812 124496 623824
rect 69072 623784 124496 623812
rect 69072 623772 69078 623784
rect 124490 623772 124496 623784
rect 124548 623772 124554 623824
rect 136634 623772 136640 623824
rect 136692 623812 136698 623824
rect 168742 623812 168748 623824
rect 136692 623784 168748 623812
rect 136692 623772 136698 623784
rect 168742 623772 168748 623784
rect 168800 623772 168806 623824
rect 204254 623772 204260 623824
rect 204312 623812 204318 623824
rect 277670 623812 277676 623824
rect 204312 623784 277676 623812
rect 204312 623772 204318 623784
rect 277670 623772 277676 623784
rect 277728 623772 277734 623824
rect 217962 622820 217968 622872
rect 218020 622860 218026 622872
rect 228726 622860 228732 622872
rect 218020 622832 228732 622860
rect 218020 622820 218026 622832
rect 228726 622820 228732 622832
rect 228784 622820 228790 622872
rect 126238 622752 126244 622804
rect 126296 622792 126302 622804
rect 177850 622792 177856 622804
rect 126296 622764 177856 622792
rect 126296 622752 126302 622764
rect 177850 622752 177856 622764
rect 177908 622752 177914 622804
rect 214558 622752 214564 622804
rect 214616 622792 214622 622804
rect 257614 622792 257620 622804
rect 214616 622764 257620 622792
rect 214616 622752 214622 622764
rect 257614 622752 257620 622764
rect 257672 622752 257678 622804
rect 136358 622684 136364 622736
rect 136416 622724 136422 622736
rect 145558 622724 145564 622736
rect 136416 622696 145564 622724
rect 136416 622684 136422 622696
rect 145558 622684 145564 622696
rect 145616 622684 145622 622736
rect 204346 622684 204352 622736
rect 204404 622724 204410 622736
rect 222838 622724 222844 622736
rect 204404 622696 222844 622724
rect 204404 622684 204410 622696
rect 222838 622684 222844 622696
rect 222896 622684 222902 622736
rect 56318 622616 56324 622668
rect 56376 622656 56382 622668
rect 74626 622656 74632 622668
rect 56376 622628 74632 622656
rect 56376 622616 56382 622628
rect 74626 622616 74632 622628
rect 74684 622616 74690 622668
rect 135070 622616 135076 622668
rect 135128 622656 135134 622668
rect 149146 622656 149152 622668
rect 135128 622628 149152 622656
rect 135128 622616 135134 622628
rect 149146 622616 149152 622628
rect 149204 622616 149210 622668
rect 208394 622616 208400 622668
rect 208452 622656 208458 622668
rect 240318 622656 240324 622668
rect 208452 622628 240324 622656
rect 208452 622616 208458 622628
rect 240318 622616 240324 622628
rect 240376 622616 240382 622668
rect 54938 622548 54944 622600
rect 54996 622588 55002 622600
rect 65518 622588 65524 622600
rect 54996 622560 65524 622588
rect 54996 622548 55002 622560
rect 65518 622548 65524 622560
rect 65576 622548 65582 622600
rect 134886 622548 134892 622600
rect 134944 622588 134950 622600
rect 154574 622588 154580 622600
rect 134944 622560 154580 622588
rect 134944 622548 134950 622560
rect 154574 622548 154580 622560
rect 154632 622548 154638 622600
rect 206370 622548 206376 622600
rect 206428 622588 206434 622600
rect 248690 622588 248696 622600
rect 206428 622560 248696 622588
rect 206428 622548 206434 622560
rect 248690 622548 248696 622560
rect 248748 622548 248754 622600
rect 56410 622480 56416 622532
rect 56468 622520 56474 622532
rect 71222 622520 71228 622532
rect 56468 622492 71228 622520
rect 56468 622480 56474 622492
rect 71222 622480 71228 622492
rect 71280 622480 71286 622532
rect 134978 622480 134984 622532
rect 135036 622520 135042 622532
rect 142982 622520 142988 622532
rect 135036 622492 142988 622520
rect 135036 622480 135042 622492
rect 142982 622480 142988 622492
rect 143040 622480 143046 622532
rect 211798 622480 211804 622532
rect 211856 622520 211862 622532
rect 266262 622520 266268 622532
rect 211856 622492 266268 622520
rect 211856 622480 211862 622492
rect 266262 622480 266268 622492
rect 266320 622480 266326 622532
rect 280706 622480 280712 622532
rect 280764 622480 280770 622532
rect 55030 622412 55036 622464
rect 55088 622452 55094 622464
rect 62942 622452 62948 622464
rect 55088 622424 62948 622452
rect 55088 622412 55094 622424
rect 62942 622412 62948 622424
rect 63000 622412 63006 622464
rect 136542 622412 136548 622464
rect 136600 622452 136606 622464
rect 218698 622452 218704 622464
rect 136600 622424 218704 622452
rect 136600 622412 136606 622424
rect 218698 622412 218704 622424
rect 218756 622412 218762 622464
rect 118234 622344 118240 622396
rect 118292 622384 118298 622396
rect 121546 622384 121552 622396
rect 118292 622356 121552 622384
rect 118292 622344 118298 622356
rect 121546 622344 121552 622356
rect 121604 622344 121610 622396
rect 198274 622344 198280 622396
rect 198332 622384 198338 622396
rect 201494 622384 201500 622396
rect 198332 622356 201500 622384
rect 198332 622344 198338 622356
rect 201494 622344 201500 622356
rect 201552 622344 201558 622396
rect 217318 622344 217324 622396
rect 217376 622384 217382 622396
rect 219710 622384 219716 622396
rect 217376 622356 219716 622384
rect 217376 622344 217382 622356
rect 219710 622344 219716 622356
rect 219768 622344 219774 622396
rect 280724 622328 280752 622480
rect 280706 622276 280712 622328
rect 280764 622276 280770 622328
rect 435358 621800 435364 621852
rect 435416 621840 435422 621852
rect 474826 621840 474832 621852
rect 435416 621812 474832 621840
rect 435416 621800 435422 621812
rect 474826 621800 474832 621812
rect 474884 621800 474890 621852
rect 432690 621732 432696 621784
rect 432748 621772 432754 621784
rect 498010 621772 498016 621784
rect 432748 621744 498016 621772
rect 432748 621732 432754 621744
rect 498010 621732 498016 621744
rect 498068 621732 498074 621784
rect 429838 621664 429844 621716
rect 429896 621704 429902 621716
rect 505738 621704 505744 621716
rect 429896 621676 505744 621704
rect 429896 621664 429902 621676
rect 505738 621664 505744 621676
rect 505796 621664 505802 621716
rect 482554 620984 482560 621036
rect 482612 621024 482618 621036
rect 509878 621024 509884 621036
rect 482612 620996 509884 621024
rect 482612 620984 482618 620996
rect 509878 620984 509884 620996
rect 509936 620984 509942 621036
rect 213178 619624 213184 619676
rect 213236 619664 213242 619676
rect 216674 619664 216680 619676
rect 213236 619636 216680 619664
rect 213236 619624 213242 619636
rect 216674 619624 216680 619636
rect 216732 619624 216738 619676
rect 302878 619624 302884 619676
rect 302936 619664 302942 619676
rect 317966 619664 317972 619676
rect 302936 619636 317972 619664
rect 302936 619624 302942 619636
rect 317966 619624 317972 619636
rect 318024 619624 318030 619676
rect 432598 619556 432604 619608
rect 432656 619596 432662 619608
rect 456794 619596 456800 619608
rect 432656 619568 456800 619596
rect 432656 619556 432662 619568
rect 456794 619556 456800 619568
rect 456852 619556 456858 619608
rect 208486 616836 208492 616888
rect 208544 616876 208550 616888
rect 216674 616876 216680 616888
rect 208544 616848 216680 616876
rect 208544 616836 208550 616848
rect 216674 616836 216680 616848
rect 216732 616836 216738 616888
rect 286318 615476 286324 615528
rect 286376 615516 286382 615528
rect 317966 615516 317972 615528
rect 286376 615488 317972 615516
rect 286376 615476 286382 615488
rect 317966 615476 317972 615488
rect 318024 615476 318030 615528
rect 428458 611260 428464 611312
rect 428516 611300 428522 611312
rect 456794 611300 456800 611312
rect 428516 611272 456800 611300
rect 428516 611260 428522 611272
rect 456794 611260 456800 611272
rect 456852 611260 456858 611312
rect 307018 609968 307024 610020
rect 307076 610008 307082 610020
rect 317874 610008 317880 610020
rect 307076 609980 317880 610008
rect 307076 609968 307082 609980
rect 317874 609968 317880 609980
rect 317932 609968 317938 610020
rect 132494 607180 132500 607232
rect 132552 607220 132558 607232
rect 136726 607220 136732 607232
rect 132552 607192 136732 607220
rect 132552 607180 132558 607192
rect 136726 607180 136732 607192
rect 136784 607180 136790 607232
rect 204898 607180 204904 607232
rect 204956 607220 204962 607232
rect 216674 607220 216680 607232
rect 204956 607192 216680 607220
rect 204956 607180 204962 607192
rect 216674 607180 216680 607192
rect 216732 607180 216738 607232
rect 304258 605820 304264 605872
rect 304316 605860 304322 605872
rect 317966 605860 317972 605872
rect 304316 605832 317972 605860
rect 304316 605820 304322 605832
rect 317966 605820 317972 605832
rect 318024 605820 318030 605872
rect 289078 600312 289084 600364
rect 289136 600352 289142 600364
rect 317598 600352 317604 600364
rect 289136 600324 317604 600352
rect 289136 600312 289142 600324
rect 317598 600312 317604 600324
rect 317656 600312 317662 600364
rect 286410 596164 286416 596216
rect 286468 596204 286474 596216
rect 317598 596204 317604 596216
rect 286468 596176 317604 596204
rect 286468 596164 286474 596176
rect 317598 596164 317604 596176
rect 317656 596164 317662 596216
rect 134518 594804 134524 594856
rect 134576 594844 134582 594856
rect 136542 594844 136548 594856
rect 134576 594816 136548 594844
rect 134576 594804 134582 594816
rect 136542 594804 136548 594816
rect 136600 594804 136606 594856
rect 207014 593376 207020 593428
rect 207072 593416 207078 593428
rect 216674 593416 216680 593428
rect 207072 593388 216680 593416
rect 207072 593376 207078 593388
rect 216674 593376 216680 593388
rect 216732 593376 216738 593428
rect 210510 589364 210516 589416
rect 210568 589404 210574 589416
rect 216674 589404 216680 589416
rect 210568 589376 216680 589404
rect 210568 589364 210574 589376
rect 216674 589364 216680 589376
rect 216732 589364 216738 589416
rect 124122 589296 124128 589348
rect 124180 589336 124186 589348
rect 131758 589336 131764 589348
rect 124180 589308 131764 589336
rect 124180 589296 124186 589308
rect 131758 589296 131764 589308
rect 131816 589296 131822 589348
rect 134610 589296 134616 589348
rect 134668 589336 134674 589348
rect 136910 589336 136916 589348
rect 134668 589308 136916 589336
rect 134668 589296 134674 589308
rect 136910 589296 136916 589308
rect 136968 589296 136974 589348
rect 204162 589296 204168 589348
rect 204220 589336 204226 589348
rect 216766 589336 216772 589348
rect 204220 589308 216772 589336
rect 204220 589296 204226 589308
rect 216766 589296 216772 589308
rect 216824 589296 216830 589348
rect 283558 589296 283564 589348
rect 283616 589336 283622 589348
rect 302234 589336 302240 589348
rect 283616 589308 302240 589336
rect 283616 589296 283622 589308
rect 302234 589296 302240 589308
rect 302292 589296 302298 589348
rect 211154 586848 211160 586900
rect 211212 586888 211218 586900
rect 216674 586888 216680 586900
rect 211212 586860 216680 586888
rect 211212 586848 211218 586860
rect 216674 586848 216680 586860
rect 216732 586848 216738 586900
rect 300118 586508 300124 586560
rect 300176 586548 300182 586560
rect 317414 586548 317420 586560
rect 300176 586520 317420 586548
rect 300176 586508 300182 586520
rect 317414 586508 317420 586520
rect 317472 586508 317478 586560
rect 57514 583720 57520 583772
rect 57572 583760 57578 583772
rect 58618 583760 58624 583772
rect 57572 583732 58624 583760
rect 57572 583720 57578 583732
rect 58618 583720 58624 583732
rect 58676 583720 58682 583772
rect 291838 582360 291844 582412
rect 291896 582400 291902 582412
rect 317966 582400 317972 582412
rect 291896 582372 317972 582400
rect 291896 582360 291902 582372
rect 317966 582360 317972 582372
rect 318024 582360 318030 582412
rect 217686 581680 217692 581732
rect 217744 581720 217750 581732
rect 218698 581720 218704 581732
rect 217744 581692 218704 581720
rect 217744 581680 217750 581692
rect 218698 581680 218704 581692
rect 218756 581680 218762 581732
rect 509878 578144 509884 578196
rect 509936 578184 509942 578196
rect 580166 578184 580172 578196
rect 509936 578156 580172 578184
rect 509936 578144 509942 578156
rect 580166 578144 580172 578156
rect 580224 578144 580230 578196
rect 125594 576852 125600 576904
rect 125652 576892 125658 576904
rect 136726 576892 136732 576904
rect 125652 576864 136732 576892
rect 125652 576852 125658 576864
rect 136726 576852 136732 576864
rect 136784 576852 136790 576904
rect 287698 576852 287704 576904
rect 287756 576892 287762 576904
rect 317874 576892 317880 576904
rect 287756 576864 317880 576892
rect 287756 576852 287762 576864
rect 317874 576852 317880 576864
rect 317932 576852 317938 576904
rect 206554 574064 206560 574116
rect 206612 574104 206618 574116
rect 216674 574104 216680 574116
rect 206612 574076 216680 574104
rect 206612 574064 206618 574076
rect 216674 574064 216680 574076
rect 216732 574064 216738 574116
rect 57330 572296 57336 572348
rect 57388 572336 57394 572348
rect 58710 572336 58716 572348
rect 57388 572308 58716 572336
rect 57388 572296 57394 572308
rect 58710 572296 58716 572308
rect 58768 572296 58774 572348
rect 210602 571344 210608 571396
rect 210660 571384 210666 571396
rect 216674 571384 216680 571396
rect 210660 571356 216680 571384
rect 210660 571344 210666 571356
rect 216674 571344 216680 571356
rect 216732 571344 216738 571396
rect 286502 571344 286508 571396
rect 286560 571384 286566 571396
rect 317966 571384 317972 571396
rect 286560 571356 317972 571384
rect 286560 571344 286566 571356
rect 317966 571344 317972 571356
rect 318024 571344 318030 571396
rect 209038 562300 209044 562352
rect 209096 562340 209102 562352
rect 217410 562340 217416 562352
rect 209096 562312 217416 562340
rect 209096 562300 209102 562312
rect 217410 562300 217416 562312
rect 217468 562300 217474 562352
rect 319346 562300 319352 562352
rect 319404 562340 319410 562352
rect 319806 562340 319812 562352
rect 319404 562312 319812 562340
rect 319404 562300 319410 562312
rect 319806 562300 319812 562312
rect 319864 562300 319870 562352
rect 281534 562232 281540 562284
rect 281592 562272 281598 562284
rect 282086 562272 282092 562284
rect 281592 562244 282092 562272
rect 281592 562232 281598 562244
rect 282086 562232 282092 562244
rect 282144 562232 282150 562284
rect 57882 561144 57888 561196
rect 57940 561184 57946 561196
rect 134518 561184 134524 561196
rect 57940 561156 134524 561184
rect 57940 561144 57946 561156
rect 134518 561144 134524 561156
rect 134576 561144 134582 561196
rect 3418 561076 3424 561128
rect 3476 561116 3482 561128
rect 291838 561116 291844 561128
rect 3476 561088 291844 561116
rect 3476 561076 3482 561088
rect 291838 561076 291844 561088
rect 291896 561076 291902 561128
rect 217686 560260 217692 560312
rect 217744 560300 217750 560312
rect 220170 560300 220176 560312
rect 217744 560272 220176 560300
rect 217744 560260 217750 560272
rect 220170 560260 220176 560272
rect 220228 560260 220234 560312
rect 57146 560192 57152 560244
rect 57204 560232 57210 560244
rect 62114 560232 62120 560244
rect 57204 560204 62120 560232
rect 57204 560192 57210 560204
rect 62114 560192 62120 560204
rect 62172 560192 62178 560244
rect 131758 560192 131764 560244
rect 131816 560232 131822 560244
rect 216766 560232 216772 560244
rect 131816 560204 216772 560232
rect 131816 560192 131822 560204
rect 216766 560192 216772 560204
rect 216824 560232 216830 560244
rect 302234 560232 302240 560244
rect 216824 560204 302240 560232
rect 216824 560192 216830 560204
rect 302234 560192 302240 560204
rect 302292 560192 302298 560244
rect 137646 560124 137652 560176
rect 137704 560164 137710 560176
rect 140774 560164 140780 560176
rect 137704 560136 140780 560164
rect 137704 560124 137710 560136
rect 140774 560124 140780 560136
rect 140832 560124 140838 560176
rect 106274 560056 106280 560108
rect 106332 560096 106338 560108
rect 124674 560096 124680 560108
rect 106332 560068 124680 560096
rect 106332 560056 106338 560068
rect 124674 560056 124680 560068
rect 124732 560056 124738 560108
rect 98086 559988 98092 560040
rect 98144 560028 98150 560040
rect 120902 560028 120908 560040
rect 98144 560000 120908 560028
rect 98144 559988 98150 560000
rect 120902 559988 120908 560000
rect 120960 559988 120966 560040
rect 182358 559988 182364 560040
rect 182416 560028 182422 560040
rect 218882 560028 218888 560040
rect 182416 560000 218888 560028
rect 182416 559988 182422 560000
rect 218882 559988 218888 560000
rect 218940 559988 218946 560040
rect 255958 559988 255964 560040
rect 256016 560028 256022 560040
rect 282914 560028 282920 560040
rect 256016 560000 282920 560028
rect 256016 559988 256022 560000
rect 282914 559988 282920 560000
rect 282972 559988 282978 560040
rect 96798 559920 96804 559972
rect 96856 559960 96862 559972
rect 122834 559960 122840 559972
rect 96856 559932 122840 559960
rect 96856 559920 96862 559932
rect 122834 559920 122840 559932
rect 122892 559920 122898 559972
rect 164326 559920 164332 559972
rect 164384 559960 164390 559972
rect 201678 559960 201684 559972
rect 164384 559932 201684 559960
rect 164384 559920 164390 559932
rect 201678 559920 201684 559932
rect 201736 559920 201742 559972
rect 273254 559920 273260 559972
rect 273312 559960 273318 559972
rect 318242 559960 318248 559972
rect 273312 559932 318248 559960
rect 273312 559920 273318 559932
rect 318242 559920 318248 559932
rect 318300 559920 318306 559972
rect 57054 559852 57060 559904
rect 57112 559892 57118 559904
rect 67726 559892 67732 559904
rect 57112 559864 67732 559892
rect 57112 559852 57118 559864
rect 67726 559852 67732 559864
rect 67784 559852 67790 559904
rect 93854 559852 93860 559904
rect 93912 559892 93918 559904
rect 124306 559892 124312 559904
rect 93912 559864 124312 559892
rect 93912 559852 93918 559864
rect 124306 559852 124312 559864
rect 124364 559852 124370 559904
rect 157978 559852 157984 559904
rect 158036 559892 158042 559904
rect 203242 559892 203248 559904
rect 158036 559864 203248 559892
rect 158036 559852 158042 559864
rect 203242 559852 203248 559864
rect 203300 559852 203306 559904
rect 260834 559852 260840 559904
rect 260892 559892 260898 559904
rect 316862 559892 316868 559904
rect 260892 559864 316868 559892
rect 260892 559852 260898 559864
rect 316862 559852 316868 559864
rect 316920 559852 316926 559904
rect 59078 559784 59084 559836
rect 59136 559824 59142 559836
rect 82906 559824 82912 559836
rect 59136 559796 82912 559824
rect 59136 559784 59142 559796
rect 82906 559784 82912 559796
rect 82964 559784 82970 559836
rect 87046 559784 87052 559836
rect 87104 559824 87110 559836
rect 121546 559824 121552 559836
rect 87104 559796 121552 559824
rect 87104 559784 87110 559796
rect 121546 559784 121552 559796
rect 121604 559784 121610 559836
rect 139026 559784 139032 559836
rect 139084 559824 139090 559836
rect 150618 559824 150624 559836
rect 139084 559796 150624 559824
rect 139084 559784 139090 559796
rect 150618 559784 150624 559796
rect 150676 559784 150682 559836
rect 156138 559784 156144 559836
rect 156196 559824 156202 559836
rect 204530 559824 204536 559836
rect 156196 559796 204536 559824
rect 156196 559784 156202 559796
rect 204530 559784 204536 559796
rect 204588 559784 204594 559836
rect 258074 559784 258080 559836
rect 258132 559824 258138 559836
rect 316954 559824 316960 559836
rect 258132 559796 316960 559824
rect 258132 559784 258138 559796
rect 316954 559784 316960 559796
rect 317012 559784 317018 559836
rect 54846 559716 54852 559768
rect 54904 559756 54910 559768
rect 78674 559756 78680 559768
rect 54904 559728 78680 559756
rect 54904 559716 54910 559728
rect 78674 559716 78680 559728
rect 78732 559716 78738 559768
rect 85574 559716 85580 559768
rect 85632 559756 85638 559768
rect 121730 559756 121736 559768
rect 85632 559728 121736 559756
rect 85632 559716 85638 559728
rect 121730 559716 121736 559728
rect 121788 559716 121794 559768
rect 139302 559716 139308 559768
rect 139360 559756 139366 559768
rect 160094 559756 160100 559768
rect 139360 559728 160100 559756
rect 139360 559716 139366 559728
rect 160094 559716 160100 559728
rect 160152 559716 160158 559768
rect 182266 559716 182272 559768
rect 182324 559756 182330 559768
rect 281534 559756 281540 559768
rect 182324 559728 281540 559756
rect 182324 559716 182330 559728
rect 281534 559716 281540 559728
rect 281592 559716 281598 559768
rect 67634 559648 67640 559700
rect 67692 559688 67698 559700
rect 121822 559688 121828 559700
rect 67692 559660 121828 559688
rect 67692 559648 67698 559660
rect 121822 559648 121828 559660
rect 121880 559648 121886 559700
rect 137738 559648 137744 559700
rect 137796 559688 137802 559700
rect 151814 559688 151820 559700
rect 137796 559660 151820 559688
rect 137796 559648 137802 559660
rect 151814 559648 151820 559660
rect 151872 559648 151878 559700
rect 154574 559648 154580 559700
rect 154632 559688 154638 559700
rect 204438 559688 204444 559700
rect 154632 559660 204444 559688
rect 154632 559648 154638 559660
rect 204438 559648 204444 559660
rect 204496 559648 204502 559700
rect 216122 559648 216128 559700
rect 216180 559688 216186 559700
rect 283006 559688 283012 559700
rect 216180 559660 283012 559688
rect 216180 559648 216186 559660
rect 283006 559648 283012 559660
rect 283064 559648 283070 559700
rect 302234 559648 302240 559700
rect 302292 559688 302298 559700
rect 302970 559688 302976 559700
rect 302292 559660 302976 559688
rect 302292 559648 302298 559660
rect 302970 559648 302976 559660
rect 303028 559648 303034 559700
rect 63494 559580 63500 559632
rect 63552 559620 63558 559632
rect 123018 559620 123024 559632
rect 63552 559592 123024 559620
rect 63552 559580 63558 559592
rect 123018 559580 123024 559592
rect 123076 559580 123082 559632
rect 139210 559580 139216 559632
rect 139268 559620 139274 559632
rect 161658 559620 161664 559632
rect 139268 559592 161664 559620
rect 139268 559580 139274 559592
rect 161658 559580 161664 559592
rect 161716 559580 161722 559632
rect 179690 559580 179696 559632
rect 179748 559620 179754 559632
rect 282086 559620 282092 559632
rect 179748 559592 282092 559620
rect 179748 559580 179754 559592
rect 282086 559580 282092 559592
rect 282144 559580 282150 559632
rect 3418 559512 3424 559564
rect 3476 559552 3482 559564
rect 286318 559552 286324 559564
rect 3476 559524 286324 559552
rect 3476 559512 3482 559524
rect 286318 559512 286324 559524
rect 286376 559512 286382 559564
rect 217870 559308 217876 559360
rect 217928 559348 217934 559360
rect 222194 559348 222200 559360
rect 217928 559320 222200 559348
rect 217928 559308 217934 559320
rect 222194 559308 222200 559320
rect 222252 559308 222258 559360
rect 139118 559036 139124 559088
rect 139176 559076 139182 559088
rect 142154 559076 142160 559088
rect 139176 559048 142160 559076
rect 139176 559036 139182 559048
rect 142154 559036 142160 559048
rect 142212 559036 142218 559088
rect 219342 559036 219348 559088
rect 219400 559076 219406 559088
rect 223574 559076 223580 559088
rect 219400 559048 223580 559076
rect 219400 559036 219406 559048
rect 223574 559036 223580 559048
rect 223632 559036 223638 559088
rect 57422 558832 57428 558884
rect 57480 558872 57486 558884
rect 60734 558872 60740 558884
rect 57480 558844 60740 558872
rect 57480 558832 57486 558844
rect 60734 558832 60740 558844
rect 60792 558832 60798 558884
rect 100754 558764 100760 558816
rect 100812 558804 100818 558816
rect 102870 558804 102876 558816
rect 100812 558776 102876 558804
rect 100812 558764 100818 558776
rect 102870 558764 102876 558776
rect 102928 558764 102934 558816
rect 116578 558764 116584 558816
rect 116636 558804 116642 558816
rect 120166 558804 120172 558816
rect 116636 558776 120172 558804
rect 116636 558764 116642 558776
rect 120166 558764 120172 558776
rect 120224 558764 120230 558816
rect 161566 558764 161572 558816
rect 161624 558804 161630 558816
rect 168466 558804 168472 558816
rect 161624 558776 168472 558804
rect 161624 558764 161630 558776
rect 168466 558764 168472 558776
rect 168524 558764 168530 558816
rect 173894 558764 173900 558816
rect 173952 558804 173958 558816
rect 179598 558804 179604 558816
rect 173952 558776 179604 558804
rect 173952 558764 173958 558776
rect 179598 558764 179604 558776
rect 179656 558764 179662 558816
rect 225138 558764 225144 558816
rect 225196 558804 225202 558816
rect 227990 558804 227996 558816
rect 225196 558776 227996 558804
rect 225196 558764 225202 558776
rect 227990 558764 227996 558776
rect 228048 558764 228054 558816
rect 260098 558764 260104 558816
rect 260156 558804 260162 558816
rect 262766 558804 262772 558816
rect 260156 558776 262772 558804
rect 260156 558764 260162 558776
rect 262766 558764 262772 558776
rect 262824 558764 262830 558816
rect 278038 558764 278044 558816
rect 278096 558804 278102 558816
rect 280246 558804 280252 558816
rect 278096 558776 280252 558804
rect 278096 558764 278102 558776
rect 280246 558764 280252 558776
rect 280304 558764 280310 558816
rect 60274 558696 60280 558748
rect 60332 558736 60338 558748
rect 62758 558736 62764 558748
rect 60332 558708 62764 558736
rect 60332 558696 60338 558708
rect 62758 558696 62764 558708
rect 62816 558696 62822 558748
rect 119338 558696 119344 558748
rect 119396 558736 119402 558748
rect 120718 558736 120724 558748
rect 119396 558708 120724 558736
rect 119396 558696 119402 558708
rect 120718 558696 120724 558708
rect 120776 558696 120782 558748
rect 147674 558628 147680 558680
rect 147732 558668 147738 558680
rect 162302 558668 162308 558680
rect 147732 558640 162308 558668
rect 147732 558628 147738 558640
rect 162302 558628 162308 558640
rect 162360 558628 162366 558680
rect 151354 558560 151360 558612
rect 151412 558600 151418 558612
rect 164878 558600 164884 558612
rect 151412 558572 164884 558600
rect 151412 558560 151418 558572
rect 164878 558560 164884 558572
rect 164936 558560 164942 558612
rect 231946 558560 231952 558612
rect 232004 558600 232010 558612
rect 259638 558600 259644 558612
rect 232004 558572 259644 558600
rect 232004 558560 232010 558572
rect 259638 558560 259644 558572
rect 259696 558560 259702 558612
rect 142890 558492 142896 558544
rect 142948 558532 142954 558544
rect 160738 558532 160744 558544
rect 142948 558504 160744 558532
rect 142948 558492 142954 558504
rect 160738 558492 160744 558504
rect 160796 558492 160802 558544
rect 199378 558492 199384 558544
rect 199436 558532 199442 558544
rect 202966 558532 202972 558544
rect 199436 558504 202972 558532
rect 199436 558492 199442 558504
rect 202966 558492 202972 558504
rect 203024 558492 203030 558544
rect 222286 558492 222292 558544
rect 222344 558532 222350 558544
rect 253934 558532 253940 558544
rect 222344 558504 253940 558532
rect 222344 558492 222350 558504
rect 253934 558492 253940 558504
rect 253992 558492 253998 558544
rect 68738 558424 68744 558476
rect 68796 558464 68802 558476
rect 71038 558464 71044 558476
rect 68796 558436 71044 558464
rect 68796 558424 68802 558436
rect 71038 558424 71044 558436
rect 71096 558424 71102 558476
rect 82722 558424 82728 558476
rect 82780 558464 82786 558476
rect 88978 558464 88984 558476
rect 82780 558436 88984 558464
rect 82780 558424 82786 558436
rect 88978 558424 88984 558436
rect 89036 558424 89042 558476
rect 140314 558424 140320 558476
rect 140372 558464 140378 558476
rect 159358 558464 159364 558476
rect 140372 558436 159364 558464
rect 140372 558424 140378 558436
rect 159358 558424 159364 558436
rect 159416 558424 159422 558476
rect 188338 558424 188344 558476
rect 188396 558464 188402 558476
rect 200206 558464 200212 558476
rect 188396 558436 200212 558464
rect 188396 558424 188402 558436
rect 200206 558424 200212 558436
rect 200264 558424 200270 558476
rect 212626 558424 212632 558476
rect 212684 558464 212690 558476
rect 251174 558464 251180 558476
rect 212684 558436 251180 558464
rect 212684 558424 212690 558436
rect 251174 558424 251180 558436
rect 251232 558424 251238 558476
rect 77018 558356 77024 558408
rect 77076 558396 77082 558408
rect 85666 558396 85672 558408
rect 77076 558368 85672 558396
rect 77076 558356 77082 558368
rect 85666 558356 85672 558368
rect 85724 558356 85730 558408
rect 94498 558356 94504 558408
rect 94556 558396 94562 558408
rect 104158 558396 104164 558408
rect 94556 558368 104164 558396
rect 94556 558356 94562 558368
rect 104158 558356 104164 558368
rect 104216 558356 104222 558408
rect 111886 558356 111892 558408
rect 111944 558396 111950 558408
rect 123110 558396 123116 558408
rect 111944 558368 123116 558396
rect 111944 558356 111950 558368
rect 123110 558356 123116 558368
rect 123168 558356 123174 558408
rect 129734 558356 129740 558408
rect 129792 558396 129798 558408
rect 153838 558396 153844 558408
rect 129792 558368 153844 558396
rect 129792 558356 129798 558368
rect 153838 558356 153844 558368
rect 153896 558356 153902 558408
rect 154666 558356 154672 558408
rect 154724 558396 154730 558408
rect 171318 558396 171324 558408
rect 154724 558368 171324 558396
rect 154724 558356 154730 558368
rect 171318 558356 171324 558368
rect 171376 558356 171382 558408
rect 187878 558356 187884 558408
rect 187936 558396 187942 558408
rect 233878 558396 233884 558408
rect 187936 558368 233884 558396
rect 187936 558356 187942 558368
rect 233878 558356 233884 558368
rect 233936 558356 233942 558408
rect 62850 558288 62856 558340
rect 62908 558328 62914 558340
rect 80698 558328 80704 558340
rect 62908 558300 80704 558328
rect 62908 558288 62914 558300
rect 80698 558288 80704 558300
rect 80756 558288 80762 558340
rect 86034 558288 86040 558340
rect 86092 558328 86098 558340
rect 108298 558328 108304 558340
rect 86092 558300 108304 558328
rect 86092 558288 86098 558300
rect 108298 558288 108304 558300
rect 108356 558288 108362 558340
rect 112438 558288 112444 558340
rect 112496 558328 112502 558340
rect 117406 558328 117412 558340
rect 112496 558300 117412 558328
rect 112496 558288 112502 558300
rect 117406 558288 117412 558300
rect 117464 558288 117470 558340
rect 118694 558288 118700 558340
rect 118752 558328 118758 558340
rect 144914 558328 144920 558340
rect 118752 558300 144920 558328
rect 118752 558288 118758 558300
rect 144914 558288 144920 558300
rect 144972 558288 144978 558340
rect 158714 558288 158720 558340
rect 158772 558328 158778 558340
rect 182910 558328 182916 558340
rect 158772 558300 182916 558328
rect 158772 558288 158778 558300
rect 182910 558288 182916 558300
rect 182968 558288 182974 558340
rect 190454 558288 190460 558340
rect 190512 558328 190518 558340
rect 257062 558328 257068 558340
rect 190512 558300 257068 558328
rect 190512 558288 190518 558300
rect 257062 558288 257068 558300
rect 257120 558288 257126 558340
rect 269114 558288 269120 558340
rect 269172 558328 269178 558340
rect 287698 558328 287704 558340
rect 269172 558300 287704 558328
rect 269172 558288 269178 558300
rect 287698 558288 287704 558300
rect 287756 558288 287762 558340
rect 71314 558220 71320 558272
rect 71372 558260 71378 558272
rect 93946 558260 93952 558272
rect 71372 558232 93952 558260
rect 71372 558220 71378 558232
rect 93946 558220 93952 558232
rect 94004 558220 94010 558272
rect 100202 558220 100208 558272
rect 100260 558260 100266 558272
rect 115198 558260 115204 558272
rect 100260 558232 115204 558260
rect 100260 558220 100266 558232
rect 115198 558220 115204 558232
rect 115256 558220 115262 558272
rect 133966 558220 133972 558272
rect 134024 558260 134030 558272
rect 197446 558260 197452 558272
rect 134024 558232 197452 558260
rect 134024 558220 134030 558232
rect 197446 558220 197452 558232
rect 197504 558220 197510 558272
rect 199470 558220 199476 558272
rect 199528 558260 199534 558272
rect 203150 558260 203156 558272
rect 199528 558232 203156 558260
rect 199528 558220 199534 558232
rect 203150 558220 203156 558232
rect 203208 558220 203214 558272
rect 227714 558220 227720 558272
rect 227772 558260 227778 558272
rect 245654 558260 245660 558272
rect 227772 558232 245660 558260
rect 227772 558220 227778 558232
rect 245654 558220 245660 558232
rect 245712 558220 245718 558272
rect 249794 558220 249800 558272
rect 249852 558260 249858 558272
rect 319806 558260 319812 558272
rect 249852 558232 319812 558260
rect 249852 558220 249858 558232
rect 319806 558220 319812 558232
rect 319864 558220 319870 558272
rect 58894 558152 58900 558204
rect 58952 558192 58958 558204
rect 74534 558192 74540 558204
rect 58952 558164 74540 558192
rect 58952 558152 58958 558164
rect 74534 558152 74540 558164
rect 74592 558152 74598 558204
rect 79870 558152 79876 558204
rect 79928 558192 79934 558204
rect 114554 558192 114560 558204
rect 79928 558164 114560 558192
rect 79928 558152 79934 558164
rect 114554 558152 114560 558164
rect 114612 558152 114618 558204
rect 132586 558152 132592 558204
rect 132644 558192 132650 558204
rect 177022 558192 177028 558204
rect 132644 558164 177028 558192
rect 132644 558152 132650 558164
rect 177022 558152 177028 558164
rect 177080 558152 177086 558204
rect 177298 558152 177304 558204
rect 177356 558192 177362 558204
rect 188614 558192 188620 558204
rect 177356 558164 188620 558192
rect 177356 558152 177362 558164
rect 188614 558152 188620 558164
rect 188672 558152 188678 558204
rect 191834 558152 191840 558204
rect 191892 558192 191898 558204
rect 276934 558192 276940 558204
rect 191892 558164 276940 558192
rect 191892 558152 191898 558164
rect 276934 558152 276940 558164
rect 276992 558152 276998 558204
rect 71774 557880 71780 557932
rect 71832 557920 71838 557932
rect 73798 557920 73804 557932
rect 71832 557892 73804 557920
rect 71832 557880 71838 557892
rect 73798 557880 73804 557892
rect 73856 557880 73862 557932
rect 184198 557880 184204 557932
rect 184256 557920 184262 557932
rect 185486 557920 185492 557932
rect 184256 557892 185492 557920
rect 184256 557880 184262 557892
rect 185486 557880 185492 557892
rect 185544 557880 185550 557932
rect 264238 557880 264244 557932
rect 264296 557920 264302 557932
rect 265342 557920 265348 557932
rect 264296 557892 265348 557920
rect 264296 557880 264302 557892
rect 265342 557880 265348 557892
rect 265400 557880 265406 557932
rect 262858 557608 262864 557660
rect 262916 557648 262922 557660
rect 268654 557648 268660 557660
rect 262916 557620 268660 557648
rect 262916 557608 262922 557620
rect 268654 557608 268660 557620
rect 268712 557608 268718 557660
rect 64138 557540 64144 557592
rect 64196 557580 64202 557592
rect 65058 557580 65064 557592
rect 64196 557552 65064 557580
rect 64196 557540 64202 557552
rect 65058 557540 65064 557552
rect 65116 557540 65122 557592
rect 222930 557540 222936 557592
rect 222988 557580 222994 557592
rect 224402 557580 224408 557592
rect 222988 557552 224408 557580
rect 222988 557540 222994 557552
rect 224402 557540 224408 557552
rect 224460 557540 224466 557592
rect 267734 557540 267740 557592
rect 267792 557580 267798 557592
rect 317414 557580 317420 557592
rect 267792 557552 317420 557580
rect 267792 557540 267798 557552
rect 317414 557540 317420 557552
rect 317472 557540 317478 557592
rect 219250 557472 219256 557524
rect 219308 557512 219314 557524
rect 223666 557512 223672 557524
rect 219308 557484 223672 557512
rect 219308 557472 219314 557484
rect 223666 557472 223672 557484
rect 223724 557472 223730 557524
rect 178034 557064 178040 557116
rect 178092 557104 178098 557116
rect 206554 557104 206560 557116
rect 178092 557076 206560 557104
rect 178092 557064 178098 557076
rect 206554 557064 206560 557076
rect 206612 557064 206618 557116
rect 57330 556996 57336 557048
rect 57388 557036 57394 557048
rect 81710 557036 81716 557048
rect 57388 557008 81716 557036
rect 57388 556996 57394 557008
rect 81710 556996 81716 557008
rect 81768 556996 81774 557048
rect 122834 556996 122840 557048
rect 122892 557036 122898 557048
rect 202230 557036 202236 557048
rect 122892 557008 202236 557036
rect 122892 556996 122898 557008
rect 202230 556996 202236 557008
rect 202288 556996 202294 557048
rect 78858 556928 78864 556980
rect 78916 556968 78922 556980
rect 121454 556968 121460 556980
rect 78916 556940 121460 556968
rect 78916 556928 78922 556940
rect 121454 556928 121460 556940
rect 121512 556928 121518 556980
rect 137462 556928 137468 556980
rect 137520 556968 137526 556980
rect 149054 556968 149060 556980
rect 137520 556940 149060 556968
rect 137520 556928 137526 556940
rect 149054 556928 149060 556940
rect 149112 556928 149118 556980
rect 194594 556928 194600 556980
rect 194652 556968 194658 556980
rect 283558 556968 283564 556980
rect 194652 556940 283564 556968
rect 194652 556928 194658 556940
rect 283558 556928 283564 556940
rect 283616 556928 283622 556980
rect 63770 556860 63776 556912
rect 63828 556900 63834 556912
rect 122926 556900 122932 556912
rect 63828 556872 122932 556900
rect 63828 556860 63834 556872
rect 122926 556860 122932 556872
rect 122984 556860 122990 556912
rect 138474 556860 138480 556912
rect 138532 556900 138538 556912
rect 159082 556900 159088 556912
rect 138532 556872 159088 556900
rect 138532 556860 138538 556872
rect 159082 556860 159088 556872
rect 159140 556860 159146 556912
rect 159818 556860 159824 556912
rect 159876 556900 159882 556912
rect 173434 556900 173440 556912
rect 159876 556872 173440 556900
rect 159876 556860 159882 556872
rect 173434 556860 173440 556872
rect 173492 556860 173498 556912
rect 179506 556860 179512 556912
rect 179564 556900 179570 556912
rect 281626 556900 281632 556912
rect 179564 556872 281632 556900
rect 179564 556860 179570 556872
rect 281626 556860 281632 556872
rect 281684 556860 281690 556912
rect 4798 556792 4804 556844
rect 4856 556832 4862 556844
rect 318334 556832 318340 556844
rect 4856 556804 318340 556832
rect 4856 556792 4862 556804
rect 318334 556792 318340 556804
rect 318392 556792 318398 556844
rect 193214 555704 193220 555756
rect 193272 555744 193278 555756
rect 218790 555744 218796 555756
rect 193272 555716 218796 555744
rect 193272 555704 193278 555716
rect 218790 555704 218796 555716
rect 218848 555704 218854 555756
rect 143534 555636 143540 555688
rect 143592 555676 143598 555688
rect 201862 555676 201868 555688
rect 143592 555648 201868 555676
rect 143592 555636 143598 555648
rect 201862 555636 201868 555648
rect 201920 555636 201926 555688
rect 228634 555636 228640 555688
rect 228692 555676 228698 555688
rect 281718 555676 281724 555688
rect 228692 555648 281724 555676
rect 228692 555636 228698 555648
rect 281718 555636 281724 555648
rect 281776 555636 281782 555688
rect 59262 555568 59268 555620
rect 59320 555608 59326 555620
rect 92566 555608 92572 555620
rect 59320 555580 92572 555608
rect 59320 555568 59326 555580
rect 92566 555568 92572 555580
rect 92624 555568 92630 555620
rect 100386 555568 100392 555620
rect 100444 555608 100450 555620
rect 123478 555608 123484 555620
rect 100444 555580 123484 555608
rect 100444 555568 100450 555580
rect 123478 555568 123484 555580
rect 123536 555568 123542 555620
rect 126146 555568 126152 555620
rect 126204 555608 126210 555620
rect 200758 555608 200764 555620
rect 126204 555580 200764 555608
rect 126204 555568 126210 555580
rect 200758 555568 200764 555580
rect 200816 555568 200822 555620
rect 242894 555568 242900 555620
rect 242952 555608 242958 555620
rect 316770 555608 316776 555620
rect 242952 555580 316776 555608
rect 242952 555568 242958 555580
rect 316770 555568 316776 555580
rect 316828 555568 316834 555620
rect 64874 555500 64880 555552
rect 64932 555540 64938 555552
rect 122190 555540 122196 555552
rect 64932 555512 122196 555540
rect 64932 555500 64938 555512
rect 122190 555500 122196 555512
rect 122248 555500 122254 555552
rect 138658 555500 138664 555552
rect 138716 555540 138722 555552
rect 174906 555540 174912 555552
rect 138716 555512 174912 555540
rect 138716 555500 138722 555512
rect 174906 555500 174912 555512
rect 174964 555500 174970 555552
rect 181346 555500 181352 555552
rect 181404 555540 181410 555552
rect 281810 555540 281816 555552
rect 181404 555512 281816 555540
rect 181404 555500 181410 555512
rect 281810 555500 281816 555512
rect 281868 555500 281874 555552
rect 3510 555432 3516 555484
rect 3568 555472 3574 555484
rect 319806 555472 319812 555484
rect 3568 555444 319812 555472
rect 3568 555432 3574 555444
rect 319806 555432 319812 555444
rect 319864 555432 319870 555484
rect 171318 554208 171324 554260
rect 171376 554248 171382 554260
rect 203334 554248 203340 554260
rect 171376 554220 203340 554248
rect 171376 554208 171382 554220
rect 203334 554208 203340 554220
rect 203392 554208 203398 554260
rect 266538 554208 266544 554260
rect 266596 554248 266602 554260
rect 311158 554248 311164 554260
rect 266596 554220 311164 554248
rect 266596 554208 266602 554220
rect 311158 554208 311164 554220
rect 311216 554208 311222 554260
rect 73246 554140 73252 554192
rect 73304 554180 73310 554192
rect 108574 554180 108580 554192
rect 73304 554152 108580 554180
rect 73304 554140 73310 554152
rect 108574 554140 108580 554152
rect 108632 554140 108638 554192
rect 124306 554140 124312 554192
rect 124364 554180 124370 554192
rect 201126 554180 201132 554192
rect 124364 554152 201132 554180
rect 124364 554140 124370 554152
rect 201126 554140 201132 554152
rect 201184 554140 201190 554192
rect 229278 554140 229284 554192
rect 229336 554180 229342 554192
rect 281258 554180 281264 554192
rect 229336 554152 281264 554180
rect 229336 554140 229342 554152
rect 281258 554140 281264 554152
rect 281316 554140 281322 554192
rect 58526 554072 58532 554124
rect 58584 554112 58590 554124
rect 110414 554112 110420 554124
rect 58584 554084 110420 554112
rect 58584 554072 58590 554084
rect 110414 554072 110420 554084
rect 110472 554072 110478 554124
rect 197998 554072 198004 554124
rect 198056 554112 198062 554124
rect 283098 554112 283104 554124
rect 198056 554084 283104 554112
rect 198056 554072 198062 554084
rect 283098 554072 283104 554084
rect 283156 554072 283162 554124
rect 66714 554004 66720 554056
rect 66772 554044 66778 554056
rect 121178 554044 121184 554056
rect 66772 554016 121184 554044
rect 66772 554004 66778 554016
rect 121178 554004 121184 554016
rect 121236 554004 121242 554056
rect 138842 554004 138848 554056
rect 138900 554044 138906 554056
rect 160554 554044 160560 554056
rect 138900 554016 160560 554044
rect 138900 554004 138906 554016
rect 160554 554004 160560 554016
rect 160612 554004 160618 554056
rect 186314 554004 186320 554056
rect 186372 554044 186378 554056
rect 283190 554044 283196 554056
rect 186372 554016 283196 554044
rect 186372 554004 186378 554016
rect 283190 554004 283196 554016
rect 283248 554004 283254 554056
rect 219526 553596 219532 553648
rect 219584 553636 219590 553648
rect 219894 553636 219900 553648
rect 219584 553608 219900 553636
rect 219584 553596 219590 553608
rect 219894 553596 219900 553608
rect 219952 553596 219958 553648
rect 3510 553392 3516 553444
rect 3568 553432 3574 553444
rect 317966 553432 317972 553444
rect 3568 553404 317972 553432
rect 3568 553392 3574 553404
rect 317966 553392 317972 553404
rect 318024 553392 318030 553444
rect 226426 552916 226432 552968
rect 226484 552956 226490 552968
rect 280798 552956 280804 552968
rect 226484 552928 280804 552956
rect 226484 552916 226490 552928
rect 280798 552916 280804 552928
rect 280856 552916 280862 552968
rect 59446 552848 59452 552900
rect 59504 552888 59510 552900
rect 75914 552888 75920 552900
rect 59504 552860 75920 552888
rect 59504 552848 59510 552860
rect 75914 552848 75920 552860
rect 75972 552848 75978 552900
rect 88610 552848 88616 552900
rect 88668 552888 88674 552900
rect 103514 552888 103520 552900
rect 88668 552860 103520 552888
rect 88668 552848 88674 552860
rect 103514 552848 103520 552860
rect 103572 552848 103578 552900
rect 106918 552848 106924 552900
rect 106976 552888 106982 552900
rect 123386 552888 123392 552900
rect 106976 552860 123392 552888
rect 106976 552848 106982 552860
rect 123386 552848 123392 552860
rect 123444 552848 123450 552900
rect 128998 552848 129004 552900
rect 129056 552888 129062 552900
rect 203058 552888 203064 552900
rect 129056 552860 203064 552888
rect 129056 552848 129062 552860
rect 203058 552848 203064 552860
rect 203116 552848 203122 552900
rect 255314 552848 255320 552900
rect 255372 552888 255378 552900
rect 315298 552888 315304 552900
rect 255372 552860 315304 552888
rect 255372 552848 255378 552860
rect 315298 552848 315304 552860
rect 315356 552848 315362 552900
rect 75270 552780 75276 552832
rect 75328 552820 75334 552832
rect 96982 552820 96988 552832
rect 75328 552792 96988 552820
rect 75328 552780 75334 552792
rect 96982 552780 96988 552792
rect 97040 552780 97046 552832
rect 121454 552780 121460 552832
rect 121512 552820 121518 552832
rect 201034 552820 201040 552832
rect 121512 552792 201040 552820
rect 121512 552780 121518 552792
rect 201034 552780 201040 552792
rect 201092 552780 201098 552832
rect 247954 552780 247960 552832
rect 248012 552820 248018 552832
rect 319346 552820 319352 552832
rect 248012 552792 319352 552820
rect 248012 552780 248018 552792
rect 319346 552780 319352 552792
rect 319404 552780 319410 552832
rect 57698 552712 57704 552764
rect 57756 552752 57762 552764
rect 77386 552752 77392 552764
rect 57756 552724 77392 552752
rect 57756 552712 57762 552724
rect 77386 552712 77392 552724
rect 77444 552712 77450 552764
rect 80054 552712 80060 552764
rect 80112 552752 80118 552764
rect 120810 552752 120816 552764
rect 80112 552724 120816 552752
rect 80112 552712 80118 552724
rect 120810 552712 120816 552724
rect 120868 552712 120874 552764
rect 195974 552712 195980 552764
rect 196032 552752 196038 552764
rect 283282 552752 283288 552764
rect 196032 552724 283288 552752
rect 196032 552712 196038 552724
rect 283282 552712 283288 552724
rect 283340 552712 283346 552764
rect 69014 552644 69020 552696
rect 69072 552684 69078 552696
rect 114646 552684 114652 552696
rect 69072 552656 114652 552684
rect 69072 552644 69078 552656
rect 114646 552644 114652 552656
rect 114704 552644 114710 552696
rect 138934 552644 138940 552696
rect 138992 552684 138998 552696
rect 166258 552684 166264 552696
rect 138992 552656 166264 552684
rect 138992 552644 138998 552656
rect 166258 552644 166264 552656
rect 166316 552644 166322 552696
rect 179138 552644 179144 552696
rect 179196 552684 179202 552696
rect 271230 552684 271236 552696
rect 179196 552656 271236 552684
rect 179196 552644 179202 552656
rect 271230 552644 271236 552656
rect 271288 552644 271294 552696
rect 279510 552644 279516 552696
rect 279568 552684 279574 552696
rect 302878 552684 302884 552696
rect 279568 552656 302884 552684
rect 279568 552644 279574 552656
rect 302878 552644 302884 552656
rect 302936 552644 302942 552696
rect 192110 551556 192116 551608
rect 192168 551596 192174 551608
rect 217318 551596 217324 551608
rect 192168 551568 217324 551596
rect 192168 551556 192174 551568
rect 217318 551556 217324 551568
rect 217376 551556 217382 551608
rect 259454 551556 259460 551608
rect 259512 551596 259518 551608
rect 314010 551596 314016 551608
rect 259512 551568 314016 551596
rect 259512 551556 259518 551568
rect 314010 551556 314016 551568
rect 314068 551556 314074 551608
rect 80974 551488 80980 551540
rect 81032 551528 81038 551540
rect 122098 551528 122104 551540
rect 81032 551500 122104 551528
rect 81032 551488 81038 551500
rect 122098 551488 122104 551500
rect 122156 551488 122162 551540
rect 176654 551488 176660 551540
rect 176712 551528 176718 551540
rect 210510 551528 210516 551540
rect 176712 551500 210516 551528
rect 176712 551488 176718 551500
rect 210510 551488 210516 551500
rect 210568 551488 210574 551540
rect 253658 551488 253664 551540
rect 253716 551528 253722 551540
rect 316678 551528 316684 551540
rect 253716 551500 316684 551528
rect 253716 551488 253722 551500
rect 316678 551488 316684 551500
rect 316736 551488 316742 551540
rect 57514 551420 57520 551472
rect 57572 551460 57578 551472
rect 89806 551460 89812 551472
rect 57572 551432 89812 551460
rect 57572 551420 57578 551432
rect 89806 551420 89812 551432
rect 89864 551420 89870 551472
rect 93946 551420 93952 551472
rect 94004 551460 94010 551472
rect 114646 551460 114652 551472
rect 94004 551432 114652 551460
rect 94004 551420 94010 551432
rect 114646 551420 114652 551432
rect 114704 551420 114710 551472
rect 121546 551420 121552 551472
rect 121604 551460 121610 551472
rect 201586 551460 201592 551472
rect 121604 551432 201592 551460
rect 121604 551420 121610 551432
rect 201586 551420 201592 551432
rect 201644 551420 201650 551472
rect 211614 551420 211620 551472
rect 211672 551460 211678 551472
rect 280890 551460 280896 551472
rect 211672 551432 280896 551460
rect 211672 551420 211678 551432
rect 280890 551420 280896 551432
rect 280948 551420 280954 551472
rect 58986 551352 58992 551404
rect 59044 551392 59050 551404
rect 102502 551392 102508 551404
rect 59044 551364 102508 551392
rect 59044 551352 59050 551364
rect 102502 551352 102508 551364
rect 102560 551352 102566 551404
rect 144730 551352 144736 551404
rect 144788 551392 144794 551404
rect 156414 551392 156420 551404
rect 144788 551364 156420 551392
rect 144788 551352 144794 551364
rect 156414 551352 156420 551364
rect 156472 551352 156478 551404
rect 200206 551352 200212 551404
rect 200264 551392 200270 551404
rect 283466 551392 283472 551404
rect 200264 551364 283472 551392
rect 200264 551352 200270 551364
rect 283466 551352 283472 551364
rect 283524 551352 283530 551404
rect 65978 551284 65984 551336
rect 66036 551324 66042 551336
rect 123202 551324 123208 551336
rect 66036 551296 123208 551324
rect 66036 551284 66042 551296
rect 123202 551284 123208 551296
rect 123260 551284 123266 551336
rect 137186 551284 137192 551336
rect 137244 551324 137250 551336
rect 169110 551324 169116 551336
rect 137244 551296 169116 551324
rect 137244 551284 137250 551296
rect 169110 551284 169116 551296
rect 169168 551284 169174 551336
rect 186406 551284 186412 551336
rect 186464 551324 186470 551336
rect 281902 551324 281908 551336
rect 186464 551296 281908 551324
rect 186464 551284 186470 551296
rect 281902 551284 281908 551296
rect 281960 551284 281966 551336
rect 69106 550128 69112 550180
rect 69164 550168 69170 550180
rect 120994 550168 121000 550180
rect 69164 550140 121000 550168
rect 69164 550128 69170 550140
rect 120994 550128 121000 550140
rect 121052 550128 121058 550180
rect 193490 550128 193496 550180
rect 193548 550168 193554 550180
rect 213178 550168 213184 550180
rect 193548 550140 213184 550168
rect 193548 550128 193554 550140
rect 213178 550128 213184 550140
rect 213236 550128 213242 550180
rect 246482 550128 246488 550180
rect 246540 550168 246546 550180
rect 307018 550168 307024 550180
rect 246540 550140 307024 550168
rect 246540 550128 246546 550140
rect 307018 550128 307024 550140
rect 307076 550128 307082 550180
rect 80698 550060 80704 550112
rect 80756 550100 80762 550112
rect 109678 550100 109684 550112
rect 80756 550072 109684 550100
rect 80756 550060 80762 550072
rect 109678 550060 109684 550072
rect 109736 550060 109742 550112
rect 177758 550060 177764 550112
rect 177816 550100 177822 550112
rect 225046 550100 225052 550112
rect 177816 550072 225052 550100
rect 177816 550060 177822 550072
rect 225046 550060 225052 550072
rect 225104 550060 225110 550112
rect 245102 550060 245108 550112
rect 245160 550100 245166 550112
rect 312538 550100 312544 550112
rect 245160 550072 312544 550100
rect 245160 550060 245166 550072
rect 312538 550060 312544 550072
rect 312596 550060 312602 550112
rect 59538 549992 59544 550044
rect 59596 550032 59602 550044
rect 101030 550032 101036 550044
rect 59596 550004 101036 550032
rect 59596 549992 59602 550004
rect 101030 549992 101036 550004
rect 101088 549992 101094 550044
rect 142614 549992 142620 550044
rect 142672 550032 142678 550044
rect 202138 550032 202144 550044
rect 142672 550004 202144 550032
rect 142672 549992 142678 550004
rect 202138 549992 202144 550004
rect 202196 549992 202202 550044
rect 210326 549992 210332 550044
rect 210384 550032 210390 550044
rect 281166 550032 281172 550044
rect 210384 550004 281172 550032
rect 210384 549992 210390 550004
rect 281166 549992 281172 550004
rect 281224 549992 281230 550044
rect 70946 549924 70952 549976
rect 71004 549964 71010 549976
rect 121914 549964 121920 549976
rect 71004 549936 121920 549964
rect 71004 549924 71010 549936
rect 121914 549924 121920 549936
rect 121972 549924 121978 549976
rect 131206 549924 131212 549976
rect 131264 549964 131270 549976
rect 177298 549964 177304 549976
rect 131264 549936 177304 549964
rect 131264 549924 131270 549936
rect 177298 549924 177304 549936
rect 177356 549924 177362 549976
rect 189074 549924 189080 549976
rect 189132 549964 189138 549976
rect 262858 549964 262864 549976
rect 189132 549936 262864 549964
rect 189132 549924 189138 549936
rect 262858 549924 262864 549936
rect 262916 549924 262922 549976
rect 120258 549856 120264 549908
rect 120316 549896 120322 549908
rect 190546 549896 190552 549908
rect 120316 549868 190552 549896
rect 120316 549856 120322 549868
rect 190546 549856 190552 549868
rect 190604 549856 190610 549908
rect 197078 549856 197084 549908
rect 197136 549896 197142 549908
rect 283374 549896 283380 549908
rect 197136 549868 283380 549896
rect 197136 549856 197142 549868
rect 283374 549856 283380 549868
rect 283432 549856 283438 549908
rect 40034 549176 40040 549228
rect 40092 549216 40098 549228
rect 317506 549216 317512 549228
rect 40092 549188 317512 549216
rect 40092 549176 40098 549188
rect 317506 549176 317512 549188
rect 317564 549176 317570 549228
rect 199194 548700 199200 548752
rect 199252 548740 199258 548752
rect 215938 548740 215944 548752
rect 199252 548712 215944 548740
rect 199252 548700 199258 548712
rect 215938 548700 215944 548712
rect 215996 548700 216002 548752
rect 88426 548632 88432 548684
rect 88484 548672 88490 548684
rect 104894 548672 104900 548684
rect 88484 548644 104900 548672
rect 88484 548632 88490 548644
rect 104894 548632 104900 548644
rect 104952 548632 104958 548684
rect 189902 548632 189908 548684
rect 189960 548672 189966 548684
rect 206462 548672 206468 548684
rect 189960 548644 206468 548672
rect 189960 548632 189966 548644
rect 206462 548632 206468 548644
rect 206520 548632 206526 548684
rect 76742 548564 76748 548616
rect 76800 548604 76806 548616
rect 112438 548604 112444 548616
rect 76800 548576 112444 548604
rect 76800 548564 76806 548576
rect 112438 548564 112444 548576
rect 112496 548564 112502 548616
rect 138750 548564 138756 548616
rect 138808 548604 138814 548616
rect 153378 548604 153384 548616
rect 138808 548576 153384 548604
rect 138808 548564 138814 548576
rect 153378 548564 153384 548576
rect 153436 548564 153442 548616
rect 157886 548564 157892 548616
rect 157944 548604 157950 548616
rect 200942 548604 200948 548616
rect 157944 548576 200948 548604
rect 157944 548564 157950 548576
rect 200942 548564 200948 548576
rect 201000 548564 201006 548616
rect 205634 548564 205640 548616
rect 205692 548604 205698 548616
rect 264238 548604 264244 548616
rect 205692 548576 264244 548604
rect 205692 548564 205698 548576
rect 264238 548564 264244 548576
rect 264296 548564 264302 548616
rect 59170 548496 59176 548548
rect 59228 548536 59234 548548
rect 108206 548536 108212 548548
rect 59228 548508 108212 548536
rect 59228 548496 59234 548508
rect 108206 548496 108212 548508
rect 108264 548496 108270 548548
rect 136910 548496 136916 548548
rect 136968 548536 136974 548548
rect 202322 548536 202328 548548
rect 136968 548508 202328 548536
rect 136968 548496 136974 548508
rect 202322 548496 202328 548508
rect 202380 548496 202386 548548
rect 251542 548496 251548 548548
rect 251600 548536 251606 548548
rect 319714 548536 319720 548548
rect 251600 548508 319720 548536
rect 251600 548496 251606 548508
rect 319714 548496 319720 548508
rect 319772 548496 319778 548548
rect 283742 547476 283748 547528
rect 283800 547516 283806 547528
rect 304258 547516 304264 547528
rect 283800 547488 304264 547516
rect 283800 547476 283806 547488
rect 304258 547476 304264 547488
rect 304316 547476 304322 547528
rect 260190 547408 260196 547460
rect 260248 547448 260254 547460
rect 286502 547448 286508 547460
rect 260248 547420 286508 547448
rect 260248 547408 260254 547420
rect 286502 547408 286508 547420
rect 286560 547408 286566 547460
rect 57606 547340 57612 547392
rect 57664 547380 57670 547392
rect 91738 547380 91744 547392
rect 57664 547352 91744 547380
rect 57664 547340 57670 547352
rect 91738 547340 91744 547352
rect 91796 547340 91802 547392
rect 140498 547340 140504 547392
rect 140556 547380 140562 547392
rect 188338 547380 188344 547392
rect 140556 547352 188344 547380
rect 140556 547340 140562 547352
rect 188338 547340 188344 547352
rect 188396 547340 188402 547392
rect 190638 547340 190644 547392
rect 190696 547380 190702 547392
rect 204898 547380 204904 547392
rect 190696 547352 204904 547380
rect 190696 547340 190702 547352
rect 204898 547340 204904 547352
rect 204956 547340 204962 547392
rect 211062 547340 211068 547392
rect 211120 547380 211126 547392
rect 235994 547380 236000 547392
rect 211120 547352 236000 547380
rect 211120 547340 211126 547352
rect 235994 547340 236000 547352
rect 236052 547340 236058 547392
rect 263686 547340 263692 547392
rect 263744 547380 263750 547392
rect 309778 547380 309784 547392
rect 263744 547352 309784 547380
rect 263744 547340 263750 547352
rect 309778 547340 309784 547352
rect 309836 547340 309842 547392
rect 84562 547272 84568 547324
rect 84620 547312 84626 547324
rect 122006 547312 122012 547324
rect 84620 547284 122012 547312
rect 84620 547272 84626 547284
rect 122006 547272 122012 547284
rect 122064 547272 122070 547324
rect 124030 547272 124036 547324
rect 124088 547312 124094 547324
rect 201770 547312 201776 547324
rect 124088 547284 201776 547312
rect 124088 547272 124094 547284
rect 201770 547272 201776 547284
rect 201828 547272 201834 547324
rect 235074 547272 235080 547324
rect 235132 547312 235138 547324
rect 319622 547312 319628 547324
rect 235132 547284 319628 547312
rect 235132 547272 235138 547284
rect 319622 547272 319628 547284
rect 319680 547272 319686 547324
rect 62758 547204 62764 547256
rect 62816 547244 62822 547256
rect 105354 547244 105360 547256
rect 62816 547216 105360 547244
rect 62816 547204 62822 547216
rect 105354 547204 105360 547216
rect 105412 547204 105418 547256
rect 185578 547204 185584 547256
rect 185636 547244 185642 547256
rect 274634 547244 274640 547256
rect 185636 547216 274640 547244
rect 185636 547204 185642 547216
rect 274634 547204 274640 547216
rect 274692 547204 274698 547256
rect 282362 547204 282368 547256
rect 282420 547244 282426 547256
rect 300118 547244 300124 547256
rect 282420 547216 300124 547244
rect 282420 547204 282426 547216
rect 300118 547204 300124 547216
rect 300176 547204 300182 547256
rect 63126 547136 63132 547188
rect 63184 547176 63190 547188
rect 110506 547176 110512 547188
rect 63184 547148 110512 547176
rect 63184 547136 63190 547148
rect 110506 547136 110512 547148
rect 110564 547136 110570 547188
rect 122650 547136 122656 547188
rect 122708 547176 122714 547188
rect 137278 547176 137284 547188
rect 122708 547148 137284 547176
rect 122708 547136 122714 547148
rect 137278 547136 137284 547148
rect 137336 547136 137342 547188
rect 147858 547136 147864 547188
rect 147916 547176 147922 547188
rect 184198 547176 184204 547188
rect 147916 547148 184204 547176
rect 147916 547136 147922 547148
rect 184198 547136 184204 547148
rect 184256 547136 184262 547188
rect 187786 547136 187792 547188
rect 187844 547176 187850 547188
rect 283650 547176 283656 547188
rect 187844 547148 283656 547176
rect 187844 547136 187850 547148
rect 283650 547136 283656 547148
rect 283708 547136 283714 547188
rect 139854 546456 139860 546508
rect 139912 546496 139918 546508
rect 141878 546496 141884 546508
rect 139912 546468 141884 546496
rect 139912 546456 139918 546468
rect 141878 546456 141884 546468
rect 141936 546456 141942 546508
rect 184934 545980 184940 546032
rect 184992 546020 184998 546032
rect 216030 546020 216036 546032
rect 184992 545992 216036 546020
rect 184992 545980 184998 545992
rect 216030 545980 216036 545992
rect 216088 545980 216094 546032
rect 138290 545912 138296 545964
rect 138348 545952 138354 545964
rect 200850 545952 200856 545964
rect 138348 545924 200856 545952
rect 138348 545912 138354 545924
rect 200850 545912 200856 545924
rect 200908 545912 200914 545964
rect 206370 545912 206376 545964
rect 206428 545952 206434 545964
rect 241514 545952 241520 545964
rect 206428 545924 241520 545952
rect 206428 545912 206434 545924
rect 241514 545912 241520 545924
rect 241572 545912 241578 545964
rect 250070 545912 250076 545964
rect 250128 545952 250134 545964
rect 289078 545952 289084 545964
rect 250128 545924 289084 545952
rect 250128 545912 250134 545924
rect 289078 545912 289084 545924
rect 289136 545912 289142 545964
rect 82446 545844 82452 545896
rect 82504 545884 82510 545896
rect 116578 545884 116584 545896
rect 82504 545856 116584 545884
rect 82504 545844 82510 545856
rect 116578 545844 116584 545856
rect 116636 545844 116642 545896
rect 139026 545844 139032 545896
rect 139084 545884 139090 545896
rect 202046 545884 202052 545896
rect 139084 545856 202052 545884
rect 139084 545844 139090 545856
rect 202046 545844 202052 545856
rect 202104 545844 202110 545896
rect 217870 545844 217876 545896
rect 217928 545884 217934 545896
rect 260098 545884 260104 545896
rect 217928 545856 260104 545884
rect 217928 545844 217934 545856
rect 260098 545844 260104 545856
rect 260156 545844 260162 545896
rect 275186 545844 275192 545896
rect 275244 545884 275250 545896
rect 313918 545884 313924 545896
rect 275244 545856 313924 545884
rect 275244 545844 275250 545856
rect 313918 545844 313924 545856
rect 313976 545844 313982 545896
rect 57238 545776 57244 545828
rect 57296 545816 57302 545828
rect 103238 545816 103244 545828
rect 57296 545788 103244 545816
rect 57296 545776 57302 545788
rect 103238 545776 103244 545788
rect 103296 545776 103302 545828
rect 198550 545776 198556 545828
rect 198608 545816 198614 545828
rect 278038 545816 278044 545828
rect 198608 545788 278044 545816
rect 198608 545776 198614 545788
rect 278038 545776 278044 545788
rect 278096 545776 278102 545828
rect 71682 545708 71688 545760
rect 71740 545748 71746 545760
rect 123570 545748 123576 545760
rect 71740 545720 123576 545748
rect 71740 545708 71746 545720
rect 123570 545708 123576 545720
rect 123628 545708 123634 545760
rect 127618 545708 127624 545760
rect 127676 545748 127682 545760
rect 194686 545748 194692 545760
rect 127676 545720 194692 545748
rect 127676 545708 127682 545720
rect 194686 545708 194692 545720
rect 194744 545708 194750 545760
rect 197814 545708 197820 545760
rect 197872 545748 197878 545760
rect 210602 545748 210608 545760
rect 197872 545720 210608 545748
rect 197872 545708 197878 545720
rect 210602 545708 210608 545720
rect 210660 545708 210666 545760
rect 234338 545708 234344 545760
rect 234396 545748 234402 545760
rect 319530 545748 319536 545760
rect 234396 545720 319536 545748
rect 234396 545708 234402 545720
rect 319530 545708 319536 545720
rect 319588 545708 319594 545760
rect 288066 545232 288072 545284
rect 288124 545272 288130 545284
rect 314194 545272 314200 545284
rect 288124 545244 314200 545272
rect 288124 545232 288130 545244
rect 314194 545232 314200 545244
rect 314252 545232 314258 545284
rect 286686 545164 286692 545216
rect 286744 545204 286750 545216
rect 314010 545204 314016 545216
rect 286744 545176 314016 545204
rect 286744 545164 286750 545176
rect 314010 545164 314016 545176
rect 314068 545164 314074 545216
rect 242250 545096 242256 545148
rect 242308 545136 242314 545148
rect 316770 545136 316776 545148
rect 242308 545108 316776 545136
rect 242308 545096 242314 545108
rect 316770 545096 316776 545108
rect 316828 545096 316834 545148
rect 168374 544552 168380 544604
rect 168432 544592 168438 544604
rect 200666 544592 200672 544604
rect 168432 544564 200672 544592
rect 168432 544552 168438 544564
rect 200666 544552 200672 544564
rect 200724 544552 200730 544604
rect 270126 544552 270132 544604
rect 270184 544592 270190 544604
rect 286410 544592 286416 544604
rect 270184 544564 286416 544592
rect 270184 544552 270190 544564
rect 286410 544552 286416 544564
rect 286468 544552 286474 544604
rect 137922 544484 137928 544536
rect 137980 544524 137986 544536
rect 149790 544524 149796 544536
rect 137980 544496 149796 544524
rect 137980 544484 137986 544496
rect 149790 544484 149796 544496
rect 149848 544484 149854 544536
rect 152642 544484 152648 544536
rect 152700 544524 152706 544536
rect 201954 544524 201960 544536
rect 152700 544496 201960 544524
rect 152700 544484 152706 544496
rect 201954 544484 201960 544496
rect 202012 544484 202018 544536
rect 219158 544484 219164 544536
rect 219216 544524 219222 544536
rect 227162 544524 227168 544536
rect 219216 544496 227168 544524
rect 219216 544484 219222 544496
rect 227162 544484 227168 544496
rect 227220 544484 227226 544536
rect 267274 544484 267280 544536
rect 267332 544524 267338 544536
rect 295978 544524 295984 544536
rect 267332 544496 295984 544524
rect 267332 544484 267338 544496
rect 295978 544484 295984 544496
rect 296036 544484 296042 544536
rect 94590 544416 94596 544468
rect 94648 544456 94654 544468
rect 123294 544456 123300 544468
rect 94648 544428 123300 544456
rect 94648 544416 94654 544428
rect 123294 544416 123300 544428
rect 123352 544416 123358 544468
rect 129734 544416 129740 544468
rect 129792 544456 129798 544468
rect 202874 544456 202880 544468
rect 129792 544428 202880 544456
rect 129792 544416 129798 544428
rect 202874 544416 202880 544428
rect 202932 544416 202938 544468
rect 220722 544416 220728 544468
rect 220780 544456 220786 544468
rect 247034 544456 247040 544468
rect 220780 544428 247040 544456
rect 220780 544416 220786 544428
rect 247034 544416 247040 544428
rect 247092 544416 247098 544468
rect 271598 544416 271604 544468
rect 271656 544456 271662 544468
rect 318150 544456 318156 544468
rect 271656 544428 318156 544456
rect 271656 544416 271662 544428
rect 318150 544416 318156 544428
rect 318208 544416 318214 544468
rect 71038 544348 71044 544400
rect 71096 544388 71102 544400
rect 108942 544388 108948 544400
rect 71096 544360 108948 544388
rect 71096 544348 71102 544360
rect 108942 544348 108948 544360
rect 109000 544348 109006 544400
rect 147766 544348 147772 544400
rect 147824 544388 147830 544400
rect 166994 544388 167000 544400
rect 147824 544360 167000 544388
rect 147824 544348 147830 544360
rect 166994 544348 167000 544360
rect 167052 544348 167058 544400
rect 184198 544348 184204 544400
rect 184256 544388 184262 544400
rect 281994 544388 282000 544400
rect 184256 544360 282000 544388
rect 184256 544348 184262 544360
rect 281994 544348 282000 544360
rect 282052 544348 282058 544400
rect 69106 544008 69112 544060
rect 69164 544048 69170 544060
rect 70302 544048 70308 544060
rect 69164 544020 70308 544048
rect 69164 544008 69170 544020
rect 70302 544008 70308 544020
rect 70360 544008 70366 544060
rect 104158 544008 104164 544060
rect 104216 544008 104222 544060
rect 113266 544008 113272 544060
rect 113324 544048 113330 544060
rect 121086 544048 121092 544060
rect 113324 544020 121092 544048
rect 113324 544008 113330 544020
rect 121086 544008 121092 544020
rect 121144 544008 121150 544060
rect 121546 544008 121552 544060
rect 121604 544048 121610 544060
rect 122558 544048 122564 544060
rect 121604 544020 122564 544048
rect 121604 544008 121610 544020
rect 122558 544008 122564 544020
rect 122616 544008 122622 544060
rect 290918 544008 290924 544060
rect 290976 544048 290982 544060
rect 290976 544020 296714 544048
rect 290976 544008 290982 544020
rect 63494 543872 63500 543924
rect 63552 543912 63558 543924
rect 64506 543912 64512 543924
rect 63552 543884 64512 543912
rect 63552 543872 63558 543884
rect 64506 543872 64512 543884
rect 64564 543872 64570 543924
rect 78674 543872 78680 543924
rect 78732 543912 78738 543924
rect 79594 543912 79600 543924
rect 78732 543884 79600 543912
rect 78732 543872 78738 543884
rect 79594 543872 79600 543884
rect 79652 543872 79658 543924
rect 88426 543872 88432 543924
rect 88484 543912 88490 543924
rect 89622 543912 89628 543924
rect 88484 543884 89628 543912
rect 88484 543872 88490 543884
rect 89622 543872 89628 543884
rect 89680 543872 89686 543924
rect 89806 543872 89812 543924
rect 89864 543912 89870 543924
rect 91002 543912 91008 543924
rect 89864 543884 91008 543912
rect 89864 543872 89870 543884
rect 91002 543872 91008 543884
rect 91060 543872 91066 543924
rect 100754 543872 100760 543924
rect 100812 543912 100818 543924
rect 101766 543912 101772 543924
rect 100812 543884 101772 543912
rect 100812 543872 100818 543884
rect 101766 543872 101772 543884
rect 101824 543872 101830 543924
rect 61654 543668 61660 543720
rect 61712 543708 61718 543720
rect 64138 543708 64144 543720
rect 61712 543680 64144 543708
rect 61712 543668 61718 543680
rect 64138 543668 64144 543680
rect 64196 543668 64202 543720
rect 88978 543668 88984 543720
rect 89036 543708 89042 543720
rect 90358 543708 90364 543720
rect 89036 543680 90364 543708
rect 89036 543668 89042 543680
rect 90358 543668 90364 543680
rect 90416 543668 90422 543720
rect 104176 543708 104204 544008
rect 179506 543940 179512 543992
rect 179564 543980 179570 543992
rect 180610 543980 180616 543992
rect 179564 543952 180616 543980
rect 179564 543940 179570 543952
rect 180610 543940 180616 543952
rect 180668 543940 180674 543992
rect 293954 543940 293960 543992
rect 294012 543980 294018 543992
rect 295242 543980 295248 543992
rect 294012 543952 295248 543980
rect 294012 543940 294018 543952
rect 295242 543940 295248 543952
rect 295300 543940 295306 543992
rect 296686 543980 296714 544020
rect 314102 543980 314108 543992
rect 296686 543952 314108 543980
rect 314102 543940 314108 543952
rect 314160 543940 314166 543992
rect 106274 543872 106280 543924
rect 106332 543912 106338 543924
rect 107562 543912 107568 543924
rect 106332 543884 107568 543912
rect 106332 543872 106338 543884
rect 107562 543872 107568 543884
rect 107620 543872 107626 543924
rect 114554 543872 114560 543924
rect 114612 543912 114618 543924
rect 115382 543912 115388 543924
rect 114612 543884 115388 543912
rect 114612 543872 114618 543884
rect 115382 543872 115388 543884
rect 115440 543872 115446 543924
rect 124214 543872 124220 543924
rect 124272 543912 124278 543924
rect 125410 543912 125416 543924
rect 124272 543884 125416 543912
rect 124272 543872 124278 543884
rect 125410 543872 125416 543884
rect 125468 543872 125474 543924
rect 125594 543872 125600 543924
rect 125652 543912 125658 543924
rect 126882 543912 126888 543924
rect 125652 543884 126888 543912
rect 125652 543872 125658 543884
rect 126882 543872 126888 543884
rect 126940 543872 126946 543924
rect 136634 543872 136640 543924
rect 136692 543912 136698 543924
rect 137646 543912 137652 543924
rect 136692 543884 137652 543912
rect 136692 543872 136698 543884
rect 137646 543872 137652 543884
rect 137704 543872 137710 543924
rect 142154 543872 142160 543924
rect 142212 543912 142218 543924
rect 143350 543912 143356 543924
rect 142212 543884 143356 543912
rect 142212 543872 142218 543884
rect 143350 543872 143356 543884
rect 143408 543872 143414 543924
rect 147674 543872 147680 543924
rect 147732 543912 147738 543924
rect 148318 543912 148324 543924
rect 147732 543884 148324 543912
rect 147732 543872 147738 543884
rect 148318 543872 148324 543884
rect 148376 543872 148382 543924
rect 154574 543872 154580 543924
rect 154632 543912 154638 543924
rect 155494 543912 155500 543924
rect 154632 543884 155500 543912
rect 154632 543872 154638 543884
rect 155494 543872 155500 543884
rect 155552 543872 155558 543924
rect 158714 543872 158720 543924
rect 158772 543912 158778 543924
rect 159818 543912 159824 543924
rect 158772 543884 159824 543912
rect 158772 543872 158778 543884
rect 159818 543872 159824 543884
rect 159876 543872 159882 543924
rect 160094 543872 160100 543924
rect 160152 543912 160158 543924
rect 161290 543912 161296 543924
rect 160152 543884 161296 543912
rect 160152 543872 160158 543884
rect 161290 543872 161296 543884
rect 161348 543872 161354 543924
rect 161566 543872 161572 543924
rect 161624 543912 161630 543924
rect 162670 543912 162676 543924
rect 161624 543884 162676 543912
rect 161624 543872 161630 543884
rect 162670 543872 162676 543884
rect 162728 543872 162734 543924
rect 164326 543872 164332 543924
rect 164384 543912 164390 543924
rect 165522 543912 165528 543924
rect 164384 543884 165528 543912
rect 164384 543872 164390 543884
rect 165522 543872 165528 543884
rect 165580 543872 165586 543924
rect 186314 543872 186320 543924
rect 186372 543912 186378 543924
rect 187050 543912 187056 543924
rect 186372 543884 187056 543912
rect 186372 543872 186378 543884
rect 187050 543872 187056 543884
rect 187108 543872 187114 543924
rect 191834 543872 191840 543924
rect 191892 543912 191898 543924
rect 192754 543912 192760 543924
rect 191892 543884 192760 543912
rect 191892 543872 191898 543884
rect 192754 543872 192760 543884
rect 192812 543872 192818 543924
rect 193214 543872 193220 543924
rect 193272 543912 193278 543924
rect 194226 543912 194232 543924
rect 193272 543884 194232 543912
rect 193272 543872 193278 543884
rect 194226 543872 194232 543884
rect 194284 543872 194290 543924
rect 208394 543872 208400 543924
rect 208452 543912 208458 543924
rect 209222 543912 209228 543924
rect 208452 543884 209228 543912
rect 208452 543872 208458 543884
rect 209222 543872 209228 543884
rect 209280 543872 209286 543924
rect 212534 543872 212540 543924
rect 212592 543912 212598 543924
rect 213546 543912 213552 543924
rect 212592 543884 213552 543912
rect 212592 543872 212598 543884
rect 213546 543872 213552 543884
rect 213604 543872 213610 543924
rect 222194 543872 222200 543924
rect 222252 543912 222258 543924
rect 222838 543912 222844 543924
rect 222252 543884 222844 543912
rect 222252 543872 222258 543884
rect 222838 543872 222844 543884
rect 222896 543872 222902 543924
rect 255314 543872 255320 543924
rect 255372 543912 255378 543924
rect 256510 543912 256516 543924
rect 255372 543884 256516 543912
rect 255372 543872 255378 543884
rect 256510 543872 256516 543884
rect 256568 543872 256574 543924
rect 273254 543872 273260 543924
rect 273312 543912 273318 543924
rect 274450 543912 274456 543924
rect 273312 543884 274456 543912
rect 273312 543872 273318 543884
rect 274450 543872 274456 543884
rect 274508 543872 274514 543924
rect 285214 543872 285220 543924
rect 285272 543912 285278 543924
rect 313918 543912 313924 543924
rect 285272 543884 313924 543912
rect 285272 543872 285278 543884
rect 313918 543872 313924 543884
rect 313976 543872 313982 543924
rect 137554 543804 137560 543856
rect 137612 543844 137618 543856
rect 139762 543844 139768 543856
rect 137612 543816 139768 543844
rect 137612 543804 137618 543816
rect 139762 543804 139768 543816
rect 139820 543804 139826 543856
rect 252278 543804 252284 543856
rect 252336 543844 252342 543856
rect 317966 543844 317972 543856
rect 252336 543816 317972 543844
rect 252336 543804 252342 543816
rect 317966 543804 317972 543816
rect 318024 543804 318030 543856
rect 237926 543736 237932 543788
rect 237984 543776 237990 543788
rect 316678 543776 316684 543788
rect 237984 543748 316684 543776
rect 237984 543736 237990 543748
rect 316678 543736 316684 543748
rect 316736 543736 316742 543788
rect 106090 543708 106096 543720
rect 104176 543680 106096 543708
rect 106090 543668 106096 543680
rect 106148 543668 106154 543720
rect 108298 543668 108304 543720
rect 108356 543708 108362 543720
rect 111794 543708 111800 543720
rect 108356 543680 111800 543708
rect 108356 543668 108362 543680
rect 111794 543668 111800 543680
rect 111852 543668 111858 543720
rect 115198 543668 115204 543720
rect 115256 543708 115262 543720
rect 116118 543708 116124 543720
rect 115256 543680 116124 543708
rect 115256 543668 115262 543680
rect 116118 543668 116124 543680
rect 116176 543668 116182 543720
rect 135438 543668 135444 543720
rect 135496 543708 135502 543720
rect 137370 543708 137376 543720
rect 135496 543680 137376 543708
rect 135496 543668 135502 543680
rect 137370 543668 137376 543680
rect 137428 543668 137434 543720
rect 159358 543668 159364 543720
rect 159416 543708 159422 543720
rect 163406 543708 163412 543720
rect 159416 543680 163412 543708
rect 159416 543668 159422 543680
rect 163406 543668 163412 543680
rect 163464 543668 163470 543720
rect 165614 543668 165620 543720
rect 165672 543708 165678 543720
rect 169846 543708 169852 543720
rect 165672 543680 169852 543708
rect 165672 543668 165678 543680
rect 169846 543668 169852 543680
rect 169904 543668 169910 543720
rect 201402 543668 201408 543720
rect 201460 543708 201466 543720
rect 206278 543708 206284 543720
rect 201460 543680 206284 543708
rect 201460 543668 201466 543680
rect 206278 543668 206284 543680
rect 206336 543668 206342 543720
rect 207106 543668 207112 543720
rect 207164 543708 207170 543720
rect 209038 543708 209044 543720
rect 207164 543680 209044 543708
rect 207164 543668 207170 543680
rect 209038 543668 209044 543680
rect 209096 543668 209102 543720
rect 217226 543668 217232 543720
rect 217284 543708 217290 543720
rect 218606 543708 218612 543720
rect 217284 543680 218612 543708
rect 217284 543668 217290 543680
rect 218606 543668 218612 543680
rect 218664 543668 218670 543720
rect 219526 543668 219532 543720
rect 219584 543708 219590 543720
rect 221458 543708 221464 543720
rect 219584 543680 221464 543708
rect 219584 543668 219590 543680
rect 221458 543668 221464 543680
rect 221516 543668 221522 543720
rect 224402 543668 224408 543720
rect 224460 543708 224466 543720
rect 225782 543708 225788 543720
rect 224460 543680 225788 543708
rect 224460 543668 224466 543680
rect 225782 543668 225788 543680
rect 225840 543668 225846 543720
rect 55122 543600 55128 543652
rect 55180 543640 55186 543652
rect 67358 543640 67364 543652
rect 55180 543612 67364 543640
rect 55180 543600 55186 543612
rect 67358 543600 67364 543612
rect 67416 543600 67422 543652
rect 137830 543600 137836 543652
rect 137888 543640 137894 543652
rect 145466 543640 145472 543652
rect 137888 543612 145472 543640
rect 137888 543600 137894 543612
rect 145466 543600 145472 543612
rect 145524 543600 145530 543652
rect 164878 543600 164884 543652
rect 164936 543640 164942 543652
rect 172698 543640 172704 543652
rect 164936 543612 172704 543640
rect 164936 543600 164942 543612
rect 172698 543600 172704 543612
rect 172756 543600 172762 543652
rect 217594 543600 217600 543652
rect 217652 543640 217658 543652
rect 219250 543640 219256 543652
rect 217652 543612 219256 543640
rect 217652 543600 217658 543612
rect 219250 543600 219256 543612
rect 219308 543600 219314 543652
rect 55030 543532 55036 543584
rect 55088 543572 55094 543584
rect 88886 543572 88892 543584
rect 55088 543544 88892 543572
rect 55088 543532 55094 543544
rect 88886 543532 88892 543544
rect 88944 543532 88950 543584
rect 91094 543532 91100 543584
rect 91152 543572 91158 543584
rect 96798 543572 96804 543584
rect 91152 543544 96804 543572
rect 91152 543532 91158 543544
rect 96798 543532 96804 543544
rect 96856 543532 96862 543584
rect 110414 543532 110420 543584
rect 110472 543572 110478 543584
rect 119338 543572 119344 543584
rect 110472 543544 119344 543572
rect 110472 543532 110478 543544
rect 119338 543532 119344 543544
rect 119396 543532 119402 543584
rect 120442 543532 120448 543584
rect 120500 543572 120506 543584
rect 122650 543572 122656 543584
rect 120500 543544 122656 543572
rect 120500 543532 120506 543544
rect 122650 543532 122656 543544
rect 122708 543532 122714 543584
rect 131850 543532 131856 543584
rect 131908 543572 131914 543584
rect 133138 543572 133144 543584
rect 131908 543544 133144 543572
rect 131908 543532 131914 543544
rect 133138 543532 133144 543544
rect 133196 543532 133202 543584
rect 134978 543532 134984 543584
rect 135036 543572 135042 543584
rect 146938 543572 146944 543584
rect 135036 543544 146944 543572
rect 135036 543532 135042 543544
rect 146938 543532 146944 543544
rect 146996 543532 147002 543584
rect 57790 543464 57796 543516
rect 57848 543504 57854 543516
rect 93210 543504 93216 543516
rect 57848 543476 93216 543504
rect 57848 543464 57854 543476
rect 93210 543464 93216 543476
rect 93268 543464 93274 543516
rect 118234 543464 118240 543516
rect 118292 543504 118298 543516
rect 126238 543504 126244 543516
rect 118292 543476 126244 543504
rect 118292 543464 118298 543476
rect 126238 543464 126244 543476
rect 126296 543464 126302 543516
rect 136358 543464 136364 543516
rect 136416 543504 136422 543516
rect 156966 543504 156972 543516
rect 136416 543476 156972 543504
rect 136416 543464 136422 543476
rect 156966 543464 156972 543476
rect 157024 543464 157030 543516
rect 58710 543396 58716 543448
rect 58768 543436 58774 543448
rect 95326 543436 95332 543448
rect 58768 543408 95332 543436
rect 58768 543396 58774 543408
rect 95326 543396 95332 543408
rect 95384 543396 95390 543448
rect 96062 543396 96068 543448
rect 96120 543436 96126 543448
rect 106918 543436 106924 543448
rect 96120 543408 106924 543436
rect 96120 543396 96126 543408
rect 106918 543396 106924 543408
rect 106976 543396 106982 543448
rect 114002 543396 114008 543448
rect 114060 543436 114066 543448
rect 124490 543436 124496 543448
rect 114060 543408 124496 543436
rect 114060 543396 114066 543408
rect 124490 543396 124496 543408
rect 124548 543396 124554 543448
rect 134886 543396 134892 543448
rect 134944 543436 134950 543448
rect 157702 543436 157708 543448
rect 134944 543408 157708 543436
rect 134944 543396 134950 543408
rect 157702 543396 157708 543408
rect 157760 543396 157766 543448
rect 164142 543396 164148 543448
rect 164200 543436 164206 543448
rect 173986 543436 173992 543448
rect 164200 543408 173992 543436
rect 164200 543396 164206 543408
rect 173986 543396 173992 543408
rect 174044 543396 174050 543448
rect 199930 543396 199936 543448
rect 199988 543436 199994 543448
rect 210418 543436 210424 543448
rect 199988 543408 210424 543436
rect 199988 543396 199994 543408
rect 210418 543396 210424 543408
rect 210476 543396 210482 543448
rect 56502 543328 56508 543380
rect 56560 543368 56566 543380
rect 83918 543368 83924 543380
rect 56560 543340 83924 543368
rect 56560 543328 56566 543340
rect 83918 543328 83924 543340
rect 83976 543328 83982 543380
rect 85298 543328 85304 543380
rect 85356 543368 85362 543380
rect 122282 543368 122288 543380
rect 85356 543340 122288 543368
rect 85356 543328 85362 543340
rect 122282 543328 122288 543340
rect 122340 543328 122346 543380
rect 136450 543328 136456 543380
rect 136508 543368 136514 543380
rect 164878 543368 164884 543380
rect 136508 543340 164884 543368
rect 136508 543328 136514 543340
rect 164878 543328 164884 543340
rect 164936 543328 164942 543380
rect 195606 543328 195612 543380
rect 195664 543368 195670 543380
rect 206462 543368 206468 543380
rect 195664 543340 206468 543368
rect 195664 543328 195670 543340
rect 206462 543328 206468 543340
rect 206520 543328 206526 543380
rect 257246 543328 257252 543380
rect 257304 543368 257310 543380
rect 300578 543368 300584 543380
rect 257304 543340 300584 543368
rect 257304 543328 257310 543340
rect 300578 543328 300584 543340
rect 300636 543328 300642 543380
rect 56318 543260 56324 543312
rect 56376 543300 56382 543312
rect 99650 543300 99656 543312
rect 56376 543272 99656 543300
rect 56376 543260 56382 543272
rect 99650 543260 99656 543272
rect 99708 543260 99714 543312
rect 106826 543260 106832 543312
rect 106884 543300 106890 543312
rect 124398 543300 124404 543312
rect 106884 543272 124404 543300
rect 106884 543260 106890 543272
rect 124398 543260 124404 543272
rect 124456 543260 124462 543312
rect 128262 543260 128268 543312
rect 128320 543300 128326 543312
rect 157978 543300 157984 543312
rect 128320 543272 157984 543300
rect 128320 543260 128326 543272
rect 157978 543260 157984 543272
rect 158036 543260 158042 543312
rect 160738 543260 160744 543312
rect 160796 543300 160802 543312
rect 167730 543300 167736 543312
rect 160796 543272 167736 543300
rect 160796 543260 160802 543272
rect 167730 543260 167736 543272
rect 167788 543260 167794 543312
rect 170582 543260 170588 543312
rect 170640 543300 170646 543312
rect 199378 543300 199384 543312
rect 170640 543272 199384 543300
rect 170640 543260 170646 543272
rect 199378 543260 199384 543272
rect 199436 543260 199442 543312
rect 252922 543260 252928 543312
rect 252980 543300 252986 543312
rect 300210 543300 300216 543312
rect 252980 543272 300216 543300
rect 252980 543260 252986 543272
rect 300210 543260 300216 543272
rect 300268 543260 300274 543312
rect 54938 543192 54944 543244
rect 54996 543232 55002 543244
rect 98914 543232 98920 543244
rect 54996 543204 98920 543232
rect 54996 543192 55002 543204
rect 98914 543192 98920 543204
rect 98972 543192 98978 543244
rect 103974 543192 103980 543244
rect 104032 543232 104038 543244
rect 124766 543232 124772 543244
rect 104032 543204 124772 543232
rect 104032 543192 104038 543204
rect 124766 543192 124772 543204
rect 124824 543192 124830 543244
rect 138566 543192 138572 543244
rect 138624 543232 138630 543244
rect 175550 543232 175556 543244
rect 138624 543204 175556 543232
rect 138624 543192 138630 543204
rect 175550 543192 175556 543204
rect 175608 543192 175614 543244
rect 181990 543192 181996 543244
rect 182048 543232 182054 543244
rect 197998 543232 198004 543244
rect 182048 543204 198004 543232
rect 182048 543192 182054 543204
rect 197998 543192 198004 543204
rect 198056 543192 198062 543244
rect 202138 543192 202144 543244
rect 202196 543232 202202 543244
rect 216122 543232 216128 543244
rect 202196 543204 216128 543232
rect 202196 543192 202202 543204
rect 216122 543192 216128 543204
rect 216180 543192 216186 543244
rect 217962 543192 217968 543244
rect 218020 543232 218026 543244
rect 230014 543232 230020 543244
rect 218020 543204 230020 543232
rect 218020 543192 218026 543204
rect 230014 543192 230020 543204
rect 230072 543192 230078 543244
rect 231486 543192 231492 543244
rect 231544 543232 231550 543244
rect 238754 543232 238760 543244
rect 231544 543204 238760 543232
rect 231544 543192 231550 543204
rect 238754 543192 238760 543204
rect 238812 543192 238818 543244
rect 276566 543192 276572 543244
rect 276624 543232 276630 543244
rect 318334 543232 318340 543244
rect 276624 543204 318340 543232
rect 276624 543192 276630 543204
rect 318334 543192 318340 543204
rect 318392 543192 318398 543244
rect 56410 543124 56416 543176
rect 56468 543164 56474 543176
rect 73798 543164 73804 543176
rect 56468 543136 73804 543164
rect 56468 543124 56474 543136
rect 73798 543124 73804 543136
rect 73856 543124 73862 543176
rect 78122 543124 78128 543176
rect 78180 543164 78186 543176
rect 121914 543164 121920 543176
rect 78180 543136 121920 543164
rect 78180 543124 78186 543136
rect 121914 543124 121920 543136
rect 121972 543124 121978 543176
rect 135070 543124 135076 543176
rect 135128 543164 135134 543176
rect 171962 543164 171968 543176
rect 135128 543136 171968 543164
rect 135128 543124 135134 543136
rect 171962 543124 171968 543136
rect 172020 543124 172026 543176
rect 176286 543124 176292 543176
rect 176344 543164 176350 543176
rect 214558 543164 214564 543176
rect 176344 543136 214564 543164
rect 176344 543124 176350 543136
rect 214558 543124 214564 543136
rect 214616 543124 214622 543176
rect 216398 543124 216404 543176
rect 216456 543164 216462 543176
rect 255958 543164 255964 543176
rect 216456 543136 255964 543164
rect 216456 543124 216462 543136
rect 255958 543124 255964 543136
rect 256016 543124 256022 543176
rect 257982 543124 257988 543176
rect 258040 543164 258046 543176
rect 280982 543164 280988 543176
rect 258040 543136 280988 543164
rect 258040 543124 258046 543136
rect 280982 543124 280988 543136
rect 281040 543124 281046 543176
rect 298094 543124 298100 543176
rect 298152 543164 298158 543176
rect 317046 543164 317052 543176
rect 298152 543136 317052 543164
rect 298152 543124 298158 543136
rect 317046 543124 317052 543136
rect 317104 543124 317110 543176
rect 58802 543056 58808 543108
rect 58860 543096 58866 543108
rect 116854 543096 116860 543108
rect 58860 543068 116860 543096
rect 58860 543056 58866 543068
rect 116854 543056 116860 543068
rect 116912 543056 116918 543108
rect 135162 543056 135168 543108
rect 135220 543096 135226 543108
rect 151262 543096 151268 543108
rect 135220 543068 151268 543096
rect 135220 543056 135226 543068
rect 151262 543056 151268 543068
rect 151320 543056 151326 543108
rect 154114 543056 154120 543108
rect 154172 543096 154178 543108
rect 199470 543096 199476 543108
rect 154172 543068 199476 543096
rect 154172 543056 154178 543068
rect 199470 543056 199476 543068
rect 199528 543056 199534 543108
rect 203518 543056 203524 543108
rect 203576 543096 203582 543108
rect 211798 543096 211804 543108
rect 203576 543068 211804 543096
rect 203576 543056 203582 543068
rect 211798 543056 211804 543068
rect 211856 543056 211862 543108
rect 220078 543056 220084 543108
rect 220136 543096 220142 543108
rect 232866 543096 232872 543108
rect 220136 543068 232872 543096
rect 220136 543056 220142 543068
rect 232866 543056 232872 543068
rect 232924 543056 232930 543108
rect 239398 543056 239404 543108
rect 239456 543096 239462 543108
rect 281074 543096 281080 543108
rect 239456 543068 281080 543096
rect 239456 543056 239462 543068
rect 281074 543056 281080 543068
rect 281132 543056 281138 543108
rect 295978 543056 295984 543108
rect 296036 543096 296042 543108
rect 304258 543096 304264 543108
rect 296036 543068 304264 543096
rect 296036 543056 296042 543068
rect 304258 543056 304264 543068
rect 304316 543056 304322 543108
rect 58618 542988 58624 543040
rect 58676 543028 58682 543040
rect 117590 543028 117596 543040
rect 58676 543000 117596 543028
rect 58676 542988 58682 543000
rect 117590 542988 117596 543000
rect 117648 542988 117654 543040
rect 118970 542988 118976 543040
rect 119028 543028 119034 543040
rect 134794 543028 134800 543040
rect 119028 543000 134800 543028
rect 119028 542988 119034 543000
rect 134794 542988 134800 543000
rect 134852 542988 134858 543040
rect 146202 542988 146208 543040
rect 146260 543028 146266 543040
rect 201494 543028 201500 543040
rect 146260 543000 201500 543028
rect 146260 542988 146266 543000
rect 201494 542988 201500 543000
rect 201552 542988 201558 543040
rect 202782 542988 202788 543040
rect 202840 543028 202846 543040
rect 211062 543028 211068 543040
rect 202840 543000 211068 543028
rect 202840 542988 202846 543000
rect 211062 542988 211068 543000
rect 211120 542988 211126 543040
rect 218698 542988 218704 543040
rect 218756 543028 218762 543040
rect 233602 543028 233608 543040
rect 218756 543000 233608 543028
rect 218756 542988 218762 543000
rect 233602 542988 233608 543000
rect 233660 542988 233666 543040
rect 240778 542988 240784 543040
rect 240836 543028 240842 543040
rect 284938 543028 284944 543040
rect 240836 543000 284944 543028
rect 240836 542988 240842 543000
rect 284938 542988 284944 543000
rect 284996 542988 285002 543040
rect 299566 542988 299572 543040
rect 299624 543028 299630 543040
rect 319438 543028 319444 543040
rect 299624 543000 319444 543028
rect 299624 542988 299630 543000
rect 319438 542988 319444 543000
rect 319496 542988 319502 543040
rect 280154 542920 280160 542972
rect 280212 542960 280218 542972
rect 301682 542960 301688 542972
rect 280212 542932 301688 542960
rect 280212 542920 280218 542932
rect 301682 542920 301688 542932
rect 301740 542920 301746 542972
rect 278038 542852 278044 542904
rect 278096 542892 278102 542904
rect 300394 542892 300400 542904
rect 278096 542864 300400 542892
rect 278096 542852 278102 542864
rect 300394 542852 300400 542864
rect 300452 542852 300458 542904
rect 277302 542784 277308 542836
rect 277360 542824 277366 542836
rect 301958 542824 301964 542836
rect 277360 542796 301964 542824
rect 277360 542784 277366 542796
rect 301958 542784 301964 542796
rect 302016 542784 302022 542836
rect 275922 542716 275928 542768
rect 275980 542756 275986 542768
rect 301866 542756 301872 542768
rect 275980 542728 301872 542756
rect 275980 542716 275986 542728
rect 301866 542716 301872 542728
rect 301924 542716 301930 542768
rect 270862 542648 270868 542700
rect 270920 542688 270926 542700
rect 300302 542688 300308 542700
rect 270920 542660 300308 542688
rect 270920 542648 270926 542660
rect 300302 542648 300308 542660
rect 300360 542648 300366 542700
rect 273714 542580 273720 542632
rect 273772 542620 273778 542632
rect 304350 542620 304356 542632
rect 273772 542592 304356 542620
rect 273772 542580 273778 542592
rect 304350 542580 304356 542592
rect 304408 542580 304414 542632
rect 285950 542512 285956 542564
rect 286008 542552 286014 542564
rect 300118 542552 300124 542564
rect 286008 542524 300124 542552
rect 286008 542512 286014 542524
rect 300118 542512 300124 542524
rect 300176 542512 300182 542564
rect 281626 542444 281632 542496
rect 281684 542484 281690 542496
rect 302878 542484 302884 542496
rect 281684 542456 302884 542484
rect 281684 542444 281690 542456
rect 302878 542444 302884 542456
rect 302936 542444 302942 542496
rect 237190 542376 237196 542428
rect 237248 542416 237254 542428
rect 282914 542416 282920 542428
rect 237248 542388 282920 542416
rect 237248 542376 237254 542388
rect 282914 542376 282920 542388
rect 282972 542376 282978 542428
rect 284478 542376 284484 542428
rect 284536 542416 284542 542428
rect 301406 542416 301412 542428
rect 284536 542388 301412 542416
rect 284536 542376 284542 542388
rect 301406 542376 301412 542388
rect 301464 542376 301470 542428
rect 236454 541832 236460 541884
rect 236512 541872 236518 541884
rect 304442 541872 304448 541884
rect 236512 541844 304448 541872
rect 236512 541832 236518 541844
rect 304442 541832 304448 541844
rect 304500 541832 304506 541884
rect 235810 541764 235816 541816
rect 235868 541804 235874 541816
rect 319438 541804 319444 541816
rect 235868 541776 319444 541804
rect 235868 541764 235874 541776
rect 319438 541764 319444 541776
rect 319496 541764 319502 541816
rect 268746 541696 268752 541748
rect 268804 541736 268810 541748
rect 301774 541736 301780 541748
rect 268804 541708 301780 541736
rect 268804 541696 268810 541708
rect 301774 541696 301780 541708
rect 301832 541696 301838 541748
rect 263042 541628 263048 541680
rect 263100 541668 263106 541680
rect 302050 541668 302056 541680
rect 263100 541640 302056 541668
rect 263100 541628 263106 541640
rect 302050 541628 302056 541640
rect 302108 541628 302114 541680
rect 260834 541560 260840 541612
rect 260892 541600 260898 541612
rect 317138 541600 317144 541612
rect 260892 541572 317144 541600
rect 260892 541560 260898 541572
rect 317138 541560 317144 541572
rect 317196 541560 317202 541612
rect 243630 541492 243636 541544
rect 243688 541532 243694 541544
rect 300670 541532 300676 541544
rect 243688 541504 300676 541532
rect 243688 541492 243694 541504
rect 300670 541492 300676 541504
rect 300728 541492 300734 541544
rect 244366 541424 244372 541476
rect 244424 541464 244430 541476
rect 303062 541464 303068 541476
rect 244424 541436 303068 541464
rect 244424 541424 244430 541436
rect 303062 541424 303068 541436
rect 303120 541424 303126 541476
rect 255866 541356 255872 541408
rect 255924 541396 255930 541408
rect 318150 541396 318156 541408
rect 255924 541368 318156 541396
rect 255924 541356 255930 541368
rect 318150 541356 318156 541368
rect 318208 541356 318214 541408
rect 240042 541288 240048 541340
rect 240100 541328 240106 541340
rect 303154 541328 303160 541340
rect 240100 541300 303160 541328
rect 240100 541288 240106 541300
rect 303154 541288 303160 541300
rect 303212 541288 303218 541340
rect 254394 541220 254400 541272
rect 254452 541260 254458 541272
rect 319714 541260 319720 541272
rect 254452 541232 319720 541260
rect 254452 541220 254458 541232
rect 319714 541220 319720 541232
rect 319772 541220 319778 541272
rect 283098 541152 283104 541204
rect 283156 541192 283162 541204
rect 316954 541192 316960 541204
rect 283156 541164 316960 541192
rect 283156 541152 283162 541164
rect 316954 541152 316960 541164
rect 317012 541152 317018 541204
rect 249426 541084 249432 541136
rect 249484 541124 249490 541136
rect 317966 541124 317972 541136
rect 249484 541096 317972 541124
rect 249484 541084 249490 541096
rect 317966 541084 317972 541096
rect 318024 541084 318030 541136
rect 247218 541016 247224 541068
rect 247276 541056 247282 541068
rect 319622 541056 319628 541068
rect 247276 541028 319628 541056
rect 247276 541016 247282 541028
rect 319622 541016 319628 541028
rect 319680 541016 319686 541068
rect 272334 540948 272340 541000
rect 272392 540988 272398 541000
rect 300486 540988 300492 541000
rect 272392 540960 300492 540988
rect 272392 540948 272398 540960
rect 300486 540948 300492 540960
rect 300544 540948 300550 541000
rect 293770 540608 293776 540660
rect 293828 540648 293834 540660
rect 293828 540620 296714 540648
rect 293828 540608 293834 540620
rect 296686 540580 296714 540620
rect 314286 540580 314292 540592
rect 296686 540552 314292 540580
rect 314286 540540 314292 540552
rect 314344 540540 314350 540592
rect 287330 540472 287336 540524
rect 287388 540512 287394 540524
rect 314378 540512 314384 540524
rect 287388 540484 314384 540512
rect 287388 540472 287394 540484
rect 314378 540472 314384 540484
rect 314436 540472 314442 540524
rect 278774 540404 278780 540456
rect 278832 540444 278838 540456
rect 301498 540444 301504 540456
rect 278832 540416 301504 540444
rect 278832 540404 278838 540416
rect 301498 540404 301504 540416
rect 301556 540404 301562 540456
rect 265894 540336 265900 540388
rect 265952 540376 265958 540388
rect 307018 540376 307024 540388
rect 265952 540348 307024 540376
rect 265952 540336 265958 540348
rect 307018 540336 307024 540348
rect 307076 540336 307082 540388
rect 265158 540268 265164 540320
rect 265216 540308 265222 540320
rect 312538 540308 312544 540320
rect 265216 540280 312544 540308
rect 265216 540268 265222 540280
rect 312538 540268 312544 540280
rect 312596 540268 312602 540320
rect 273070 540200 273076 540252
rect 273128 540240 273134 540252
rect 319806 540240 319812 540252
rect 273128 540212 319812 540240
rect 273128 540200 273134 540212
rect 319806 540200 319812 540212
rect 319864 540200 319870 540252
rect 262306 540132 262312 540184
rect 262364 540172 262370 540184
rect 318426 540172 318432 540184
rect 262364 540144 318432 540172
rect 262364 540132 262370 540144
rect 318426 540132 318432 540144
rect 318484 540132 318490 540184
rect 3602 540064 3608 540116
rect 3660 540104 3666 540116
rect 319346 540104 319352 540116
rect 3660 540076 319352 540104
rect 3660 540064 3666 540076
rect 319346 540064 319352 540076
rect 319404 540064 319410 540116
rect 301498 539520 301504 539572
rect 301556 539560 301562 539572
rect 318058 539560 318064 539572
rect 301556 539532 318064 539560
rect 301556 539520 301562 539532
rect 318058 539520 318064 539532
rect 318116 539520 318122 539572
rect 304442 535372 304448 535424
rect 304500 535412 304506 535424
rect 317598 535412 317604 535424
rect 304500 535384 317604 535412
rect 304500 535372 304506 535384
rect 317598 535372 317604 535384
rect 317656 535372 317662 535424
rect 302234 532176 302240 532228
rect 302292 532216 302298 532228
rect 304442 532216 304448 532228
rect 302292 532188 304448 532216
rect 302292 532176 302298 532188
rect 304442 532176 304448 532188
rect 304500 532176 304506 532228
rect 300670 529864 300676 529916
rect 300728 529904 300734 529916
rect 317598 529904 317604 529916
rect 300728 529876 317604 529904
rect 300728 529864 300734 529876
rect 317598 529864 317604 529876
rect 317656 529864 317662 529916
rect 303154 525716 303160 525768
rect 303212 525756 303218 525768
rect 317598 525756 317604 525768
rect 303212 525728 317604 525756
rect 303212 525716 303218 525728
rect 317598 525716 317604 525728
rect 317656 525716 317662 525768
rect 431218 525376 431224 525428
rect 431276 525416 431282 525428
rect 431402 525416 431408 525428
rect 431276 525388 431408 525416
rect 431276 525376 431282 525388
rect 431402 525376 431408 525388
rect 431460 525376 431466 525428
rect 430942 525240 430948 525292
rect 431000 525280 431006 525292
rect 431218 525280 431224 525292
rect 431000 525252 431224 525280
rect 431000 525240 431006 525252
rect 431218 525240 431224 525252
rect 431276 525240 431282 525292
rect 430574 524968 430580 525020
rect 430632 525008 430638 525020
rect 430850 525008 430856 525020
rect 430632 524980 430856 525008
rect 430632 524968 430638 524980
rect 430850 524968 430856 524980
rect 430908 524968 430914 525020
rect 319254 523676 319260 523728
rect 319312 523716 319318 523728
rect 319622 523716 319628 523728
rect 319312 523688 319628 523716
rect 319312 523676 319318 523688
rect 319622 523676 319628 523688
rect 319680 523676 319686 523728
rect 314194 520208 314200 520260
rect 314252 520248 314258 520260
rect 511994 520248 512000 520260
rect 314252 520220 512000 520248
rect 314252 520208 314258 520220
rect 511994 520208 512000 520220
rect 512052 520208 512058 520260
rect 302970 520140 302976 520192
rect 303028 520180 303034 520192
rect 457622 520180 457628 520192
rect 303028 520152 457628 520180
rect 303028 520140 303034 520152
rect 457622 520140 457628 520152
rect 457680 520140 457686 520192
rect 317230 520072 317236 520124
rect 317288 520112 317294 520124
rect 457530 520112 457536 520124
rect 317288 520084 457536 520112
rect 317288 520072 317294 520084
rect 457530 520072 457536 520084
rect 457588 520072 457594 520124
rect 300302 520004 300308 520056
rect 300360 520044 300366 520056
rect 430942 520044 430948 520056
rect 300360 520016 430948 520044
rect 300360 520004 300366 520016
rect 430942 520004 430948 520016
rect 431000 520004 431006 520056
rect 300394 519936 300400 519988
rect 300452 519976 300458 519988
rect 430850 519976 430856 519988
rect 300452 519948 430856 519976
rect 300452 519936 300458 519948
rect 430850 519936 430856 519948
rect 430908 519936 430914 519988
rect 300578 519868 300584 519920
rect 300636 519908 300642 519920
rect 431310 519908 431316 519920
rect 300636 519880 431316 519908
rect 300636 519868 300642 519880
rect 431310 519868 431316 519880
rect 431368 519868 431374 519920
rect 301958 519800 301964 519852
rect 302016 519840 302022 519852
rect 431218 519840 431224 519852
rect 302016 519812 431224 519840
rect 302016 519800 302022 519812
rect 431218 519800 431224 519812
rect 431276 519800 431282 519852
rect 301682 519732 301688 519784
rect 301740 519772 301746 519784
rect 430574 519772 430580 519784
rect 301740 519744 430580 519772
rect 301740 519732 301746 519744
rect 430574 519732 430580 519744
rect 430632 519732 430638 519784
rect 319530 519664 319536 519716
rect 319588 519704 319594 519716
rect 431402 519704 431408 519716
rect 319588 519676 431408 519704
rect 319588 519664 319594 519676
rect 431402 519664 431408 519676
rect 431460 519664 431466 519716
rect 301866 519188 301872 519240
rect 301924 519228 301930 519240
rect 351270 519228 351276 519240
rect 301924 519200 351276 519228
rect 301924 519188 301930 519200
rect 351270 519188 351276 519200
rect 351328 519188 351334 519240
rect 305638 519120 305644 519172
rect 305696 519160 305702 519172
rect 369302 519160 369308 519172
rect 305696 519132 369308 519160
rect 305696 519120 305702 519132
rect 369302 519120 369308 519132
rect 369360 519120 369366 519172
rect 304350 519052 304356 519104
rect 304408 519092 304414 519104
rect 396902 519092 396908 519104
rect 304408 519064 396908 519092
rect 304408 519052 304414 519064
rect 396902 519052 396908 519064
rect 396960 519052 396966 519104
rect 318334 518984 318340 519036
rect 318392 519024 318398 519036
rect 414934 519024 414940 519036
rect 318392 518996 414940 519024
rect 318392 518984 318398 518996
rect 414934 518984 414940 518996
rect 414992 518984 414998 519036
rect 320082 518956 320088 518968
rect 319640 518928 320088 518956
rect 312538 518848 312544 518900
rect 312596 518888 312602 518900
rect 319640 518888 319668 518928
rect 320082 518916 320088 518928
rect 320140 518916 320146 518968
rect 324866 518916 324872 518968
rect 324924 518956 324930 518968
rect 429194 518956 429200 518968
rect 324924 518928 429200 518956
rect 324924 518916 324930 518928
rect 429194 518916 429200 518928
rect 429252 518916 429258 518968
rect 312596 518860 319668 518888
rect 312596 518848 312602 518860
rect 319714 518848 319720 518900
rect 319772 518888 319778 518900
rect 346670 518888 346676 518900
rect 319772 518860 346676 518888
rect 319772 518848 319778 518860
rect 346670 518848 346676 518860
rect 346728 518848 346734 518900
rect 319438 518780 319444 518832
rect 319496 518820 319502 518832
rect 333238 518820 333244 518832
rect 319496 518792 333244 518820
rect 319496 518780 319502 518792
rect 333238 518780 333244 518792
rect 333296 518780 333302 518832
rect 318426 518712 318432 518764
rect 318484 518752 318490 518764
rect 328730 518752 328736 518764
rect 318484 518724 328736 518752
rect 318484 518712 318490 518724
rect 328730 518712 328736 518724
rect 328788 518712 328794 518764
rect 318058 518644 318064 518696
rect 318116 518684 318122 518696
rect 423950 518684 423956 518696
rect 318116 518656 423956 518684
rect 318116 518644 318122 518656
rect 423950 518644 423956 518656
rect 424008 518644 424014 518696
rect 302050 518576 302056 518628
rect 302108 518616 302114 518628
rect 401594 518616 401600 518628
rect 302108 518588 401600 518616
rect 302108 518576 302114 518588
rect 401594 518576 401600 518588
rect 401652 518576 401658 518628
rect 318150 518508 318156 518560
rect 318208 518548 318214 518560
rect 406010 518548 406016 518560
rect 318208 518520 406016 518548
rect 318208 518508 318214 518520
rect 406010 518508 406016 518520
rect 406068 518508 406074 518560
rect 301774 518440 301780 518492
rect 301832 518480 301838 518492
rect 387886 518480 387892 518492
rect 301832 518452 387892 518480
rect 301832 518440 301838 518452
rect 387886 518440 387892 518452
rect 387944 518440 387950 518492
rect 307018 518372 307024 518424
rect 307076 518412 307082 518424
rect 383654 518412 383660 518424
rect 307076 518384 383660 518412
rect 307076 518372 307082 518384
rect 383654 518372 383660 518384
rect 383712 518372 383718 518424
rect 319806 518304 319812 518356
rect 319864 518344 319870 518356
rect 364702 518344 364708 518356
rect 319864 518316 364708 518344
rect 319864 518304 319870 518316
rect 364702 518304 364708 518316
rect 364760 518304 364766 518356
rect 319254 518236 319260 518288
rect 319312 518276 319318 518288
rect 360286 518276 360292 518288
rect 319312 518248 360292 518276
rect 319312 518236 319318 518248
rect 360286 518236 360292 518248
rect 360344 518236 360350 518288
rect 317138 518168 317144 518220
rect 317196 518208 317202 518220
rect 342254 518208 342260 518220
rect 317196 518180 342260 518208
rect 317196 518168 317202 518180
rect 342254 518168 342260 518180
rect 342312 518168 342318 518220
rect 300210 518100 300216 518152
rect 300268 518140 300274 518152
rect 431126 518140 431132 518152
rect 300268 518112 431132 518140
rect 300268 518100 300274 518112
rect 431126 518100 431132 518112
rect 431184 518100 431190 518152
rect 303062 518032 303068 518084
rect 303120 518072 303126 518084
rect 419534 518072 419540 518084
rect 303120 518044 419540 518072
rect 303120 518032 303126 518044
rect 419534 518032 419540 518044
rect 419592 518032 419598 518084
rect 300486 517964 300492 518016
rect 300544 518004 300550 518016
rect 410518 518004 410524 518016
rect 300544 517976 410524 518004
rect 300544 517964 300550 517976
rect 410518 517964 410524 517976
rect 410576 517964 410582 518016
rect 304258 517420 304264 517472
rect 304316 517460 304322 517472
rect 505094 517460 505100 517472
rect 304316 517432 505100 517460
rect 304316 517420 304322 517432
rect 505094 517420 505100 517432
rect 505152 517420 505158 517472
rect 318242 517352 318248 517404
rect 318300 517392 318306 517404
rect 512178 517392 512184 517404
rect 318300 517364 512184 517392
rect 318300 517352 318306 517364
rect 512178 517352 512184 517364
rect 512236 517352 512242 517404
rect 300118 517284 300124 517336
rect 300176 517324 300182 517336
rect 483014 517324 483020 517336
rect 300176 517296 483020 517324
rect 300176 517284 300182 517296
rect 483014 517284 483020 517296
rect 483072 517284 483078 517336
rect 317046 517216 317052 517268
rect 317104 517256 317110 517268
rect 457438 517256 457444 517268
rect 317104 517228 457444 517256
rect 317104 517216 317110 517228
rect 457438 517216 457444 517228
rect 457496 517216 457502 517268
rect 301498 517148 301504 517200
rect 301556 517188 301562 517200
rect 430758 517188 430764 517200
rect 301556 517160 430764 517188
rect 301556 517148 301562 517160
rect 430758 517148 430764 517160
rect 430816 517148 430822 517200
rect 302786 517080 302792 517132
rect 302844 517120 302850 517132
rect 431034 517120 431040 517132
rect 302844 517092 431040 517120
rect 302844 517080 302850 517092
rect 431034 517080 431040 517092
rect 431092 517080 431098 517132
rect 302878 516128 302884 516180
rect 302936 516168 302942 516180
rect 519538 516168 519544 516180
rect 302936 516140 519544 516168
rect 302936 516128 302942 516140
rect 519538 516128 519544 516140
rect 519596 516128 519602 516180
rect 314010 516060 314016 516112
rect 314068 516100 314074 516112
rect 512086 516100 512092 516112
rect 314068 516072 512092 516100
rect 314068 516060 314074 516072
rect 512086 516060 512092 516072
rect 512144 516060 512150 516112
rect 314102 515992 314108 516044
rect 314160 516032 314166 516044
rect 489914 516032 489920 516044
rect 314160 516004 489920 516032
rect 314160 515992 314166 516004
rect 489914 515992 489920 516004
rect 489972 515992 489978 516044
rect 314378 515924 314384 515976
rect 314436 515964 314442 515976
rect 474734 515964 474740 515976
rect 314436 515936 474740 515964
rect 314436 515924 314442 515936
rect 474734 515924 474740 515936
rect 474792 515924 474798 515976
rect 313918 515856 313924 515908
rect 313976 515896 313982 515908
rect 466454 515896 466460 515908
rect 313976 515868 466460 515896
rect 313976 515856 313982 515868
rect 466454 515856 466460 515868
rect 466512 515856 466518 515908
rect 314286 515788 314292 515840
rect 314344 515828 314350 515840
rect 459554 515828 459560 515840
rect 314344 515800 459560 515828
rect 314344 515788 314350 515800
rect 459554 515788 459560 515800
rect 459612 515788 459618 515840
rect 316770 515720 316776 515772
rect 316828 515760 316834 515772
rect 429562 515760 429568 515772
rect 316828 515732 429568 515760
rect 316828 515720 316834 515732
rect 429562 515720 429568 515732
rect 429620 515720 429626 515772
rect 316954 515652 316960 515704
rect 317012 515692 317018 515704
rect 429470 515692 429476 515704
rect 317012 515664 429476 515692
rect 317012 515652 317018 515664
rect 429470 515652 429476 515664
rect 429528 515652 429534 515704
rect 304442 515380 304448 515432
rect 304500 515420 304506 515432
rect 580258 515420 580264 515432
rect 304500 515392 580264 515420
rect 304500 515380 304506 515392
rect 580258 515380 580264 515392
rect 580316 515380 580322 515432
rect 316678 514700 316684 514752
rect 316736 514740 316742 514752
rect 428366 514740 428372 514752
rect 316736 514712 428372 514740
rect 316736 514700 316742 514712
rect 428366 514700 428372 514712
rect 428424 514700 428430 514752
rect 316862 514632 316868 514684
rect 316920 514672 316926 514684
rect 427814 514672 427820 514684
rect 316920 514644 427820 514672
rect 316920 514632 316926 514644
rect 427814 514632 427820 514644
rect 427872 514632 427878 514684
rect 498194 511912 498200 511964
rect 498252 511952 498258 511964
rect 580166 511952 580172 511964
rect 498252 511924 580172 511952
rect 498252 511912 498258 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 41322 509872 41328 509924
rect 41380 509912 41386 509924
rect 57698 509912 57704 509924
rect 41380 509884 57704 509912
rect 41380 509872 41386 509884
rect 57698 509872 57704 509884
rect 57756 509872 57762 509924
rect 302878 487160 302884 487212
rect 302936 487200 302942 487212
rect 520918 487200 520924 487212
rect 302936 487172 520924 487200
rect 302936 487160 302942 487172
rect 520918 487160 520924 487172
rect 520976 487160 520982 487212
rect 189074 480020 189080 480072
rect 189132 480060 189138 480072
rect 189350 480060 189356 480072
rect 189132 480032 189356 480060
rect 189132 480020 189138 480032
rect 189350 480020 189356 480032
rect 189408 480020 189414 480072
rect 160110 479816 160116 479868
rect 160168 479856 160174 479868
rect 160278 479856 160284 479868
rect 160168 479828 160284 479856
rect 160168 479816 160174 479828
rect 160278 479816 160284 479828
rect 160336 479816 160342 479868
rect 197554 479816 197560 479868
rect 197612 479856 197618 479868
rect 198274 479856 198280 479868
rect 197612 479828 198280 479856
rect 197612 479816 197618 479828
rect 198274 479816 198280 479828
rect 198332 479816 198338 479868
rect 50798 479136 50804 479188
rect 50856 479176 50862 479188
rect 84378 479176 84384 479188
rect 50856 479148 84384 479176
rect 50856 479136 50862 479148
rect 84378 479136 84384 479148
rect 84436 479136 84442 479188
rect 51994 479068 52000 479120
rect 52052 479108 52058 479120
rect 99374 479108 99380 479120
rect 52052 479080 99380 479108
rect 52052 479068 52058 479080
rect 99374 479068 99380 479080
rect 99432 479068 99438 479120
rect 50338 479000 50344 479052
rect 50396 479040 50402 479052
rect 98914 479040 98920 479052
rect 50396 479012 98920 479040
rect 50396 479000 50402 479012
rect 98914 479000 98920 479012
rect 98972 479000 98978 479052
rect 140774 479000 140780 479052
rect 140832 479040 140838 479052
rect 199102 479040 199108 479052
rect 140832 479012 199108 479040
rect 140832 479000 140838 479012
rect 199102 479000 199108 479012
rect 199160 479000 199166 479052
rect 51718 478932 51724 478984
rect 51776 478972 51782 478984
rect 100202 478972 100208 478984
rect 51776 478944 100208 478972
rect 51776 478932 51782 478944
rect 100202 478932 100208 478944
rect 100260 478932 100266 478984
rect 109034 478932 109040 478984
rect 109092 478972 109098 478984
rect 206094 478972 206100 478984
rect 109092 478944 206100 478972
rect 109092 478932 109098 478944
rect 206094 478932 206100 478944
rect 206152 478932 206158 478984
rect 45370 478864 45376 478916
rect 45428 478904 45434 478916
rect 105078 478904 105084 478916
rect 45428 478876 105084 478904
rect 45428 478864 45434 478876
rect 105078 478864 105084 478876
rect 105136 478864 105142 478916
rect 109494 478864 109500 478916
rect 109552 478904 109558 478916
rect 207106 478904 207112 478916
rect 109552 478876 207112 478904
rect 109552 478864 109558 478876
rect 207106 478864 207112 478876
rect 207164 478864 207170 478916
rect 53742 478796 53748 478848
rect 53800 478836 53806 478848
rect 74258 478836 74264 478848
rect 53800 478808 74264 478836
rect 53800 478796 53806 478808
rect 74258 478796 74264 478808
rect 74316 478796 74322 478848
rect 75362 478796 75368 478848
rect 75420 478836 75426 478848
rect 107286 478836 107292 478848
rect 75420 478808 107292 478836
rect 75420 478796 75426 478808
rect 107286 478796 107292 478808
rect 107344 478796 107350 478848
rect 149514 478796 149520 478848
rect 149572 478836 149578 478848
rect 208394 478836 208400 478848
rect 149572 478808 208400 478836
rect 149572 478796 149578 478808
rect 208394 478796 208400 478808
rect 208452 478796 208458 478848
rect 59998 478728 60004 478780
rect 60056 478768 60062 478780
rect 91830 478768 91836 478780
rect 60056 478740 91836 478768
rect 60056 478728 60062 478740
rect 91830 478728 91836 478740
rect 91888 478728 91894 478780
rect 152182 478728 152188 478780
rect 152240 478768 152246 478780
rect 210234 478768 210240 478780
rect 152240 478740 210240 478768
rect 152240 478728 152246 478740
rect 210234 478728 210240 478740
rect 210292 478728 210298 478780
rect 52178 478660 52184 478712
rect 52236 478700 52242 478712
rect 84838 478700 84844 478712
rect 52236 478672 84844 478700
rect 52236 478660 52242 478672
rect 84838 478660 84844 478672
rect 84896 478660 84902 478712
rect 154390 478660 154396 478712
rect 154448 478700 154454 478712
rect 211338 478700 211344 478712
rect 154448 478672 211344 478700
rect 154448 478660 154454 478672
rect 211338 478660 211344 478672
rect 211396 478660 211402 478712
rect 238938 478660 238944 478712
rect 238996 478700 239002 478712
rect 356698 478700 356704 478712
rect 238996 478672 356704 478700
rect 238996 478660 239002 478672
rect 356698 478660 356704 478672
rect 356756 478660 356762 478712
rect 50706 478592 50712 478644
rect 50764 478632 50770 478644
rect 68922 478632 68928 478644
rect 50764 478604 68928 478632
rect 50764 478592 50770 478604
rect 68922 478592 68928 478604
rect 68980 478592 68986 478644
rect 71314 478592 71320 478644
rect 71372 478632 71378 478644
rect 106366 478632 106372 478644
rect 71372 478604 106372 478632
rect 71372 478592 71378 478604
rect 106366 478592 106372 478604
rect 106424 478592 106430 478644
rect 153102 478592 153108 478644
rect 153160 478632 153166 478644
rect 205634 478632 205640 478644
rect 153160 478604 205640 478632
rect 153160 478592 153166 478604
rect 205634 478592 205640 478604
rect 205692 478592 205698 478644
rect 239858 478592 239864 478644
rect 239916 478632 239922 478644
rect 362310 478632 362316 478644
rect 239916 478604 362316 478632
rect 239916 478592 239922 478604
rect 362310 478592 362316 478604
rect 362368 478592 362374 478644
rect 68278 478524 68284 478576
rect 68336 478564 68342 478576
rect 104618 478564 104624 478576
rect 68336 478536 104624 478564
rect 68336 478524 68342 478536
rect 104618 478524 104624 478536
rect 104676 478524 104682 478576
rect 149146 478524 149152 478576
rect 149204 478564 149210 478576
rect 200758 478564 200764 478576
rect 149204 478536 200764 478564
rect 149204 478524 149210 478536
rect 200758 478524 200764 478536
rect 200816 478524 200822 478576
rect 240226 478524 240232 478576
rect 240284 478564 240290 478576
rect 365162 478564 365168 478576
rect 240284 478536 365168 478564
rect 240284 478524 240290 478536
rect 365162 478524 365168 478536
rect 365220 478524 365226 478576
rect 68370 478456 68376 478508
rect 68428 478496 68434 478508
rect 105538 478496 105544 478508
rect 68428 478468 105544 478496
rect 68428 478456 68434 478468
rect 105538 478456 105544 478468
rect 105596 478456 105602 478508
rect 151262 478456 151268 478508
rect 151320 478496 151326 478508
rect 201586 478496 201592 478508
rect 151320 478468 201592 478496
rect 151320 478456 151326 478468
rect 201586 478456 201592 478468
rect 201644 478456 201650 478508
rect 232314 478456 232320 478508
rect 232372 478496 232378 478508
rect 360838 478496 360844 478508
rect 232372 478468 360844 478496
rect 232372 478456 232378 478468
rect 360838 478456 360844 478468
rect 360896 478456 360902 478508
rect 54754 478388 54760 478440
rect 54812 478428 54818 478440
rect 102410 478428 102416 478440
rect 54812 478400 102416 478428
rect 54812 478388 54818 478400
rect 102410 478388 102416 478400
rect 102468 478388 102474 478440
rect 157886 478388 157892 478440
rect 157944 478428 157950 478440
rect 205634 478428 205640 478440
rect 157944 478400 205640 478428
rect 157944 478388 157950 478400
rect 205634 478388 205640 478400
rect 205692 478388 205698 478440
rect 235442 478388 235448 478440
rect 235500 478428 235506 478440
rect 366450 478428 366456 478440
rect 235500 478400 366456 478428
rect 235500 478388 235506 478400
rect 366450 478388 366456 478400
rect 366508 478388 366514 478440
rect 48038 478320 48044 478372
rect 48096 478360 48102 478372
rect 97534 478360 97540 478372
rect 48096 478332 97540 478360
rect 48096 478320 48102 478332
rect 97534 478320 97540 478332
rect 97592 478320 97598 478372
rect 153470 478320 153476 478372
rect 153528 478360 153534 478372
rect 200482 478360 200488 478372
rect 153528 478332 200488 478360
rect 153528 478320 153534 478332
rect 200482 478320 200488 478332
rect 200540 478320 200546 478372
rect 209406 478320 209412 478372
rect 209464 478360 209470 478372
rect 216674 478360 216680 478372
rect 209464 478332 216680 478360
rect 209464 478320 209470 478332
rect 216674 478320 216680 478332
rect 216732 478320 216738 478372
rect 224402 478320 224408 478372
rect 224460 478360 224466 478372
rect 358170 478360 358176 478372
rect 224460 478332 358176 478360
rect 224460 478320 224466 478332
rect 358170 478320 358176 478332
rect 358228 478320 358234 478372
rect 51902 478252 51908 478304
rect 51960 478292 51966 478304
rect 99742 478292 99748 478304
rect 51960 478264 99748 478292
rect 51960 478252 51966 478264
rect 99742 478252 99748 478264
rect 99800 478252 99806 478304
rect 138934 478252 138940 478304
rect 138992 478292 138998 478304
rect 193858 478292 193864 478304
rect 138992 478264 193864 478292
rect 138992 478252 138998 478264
rect 193858 478252 193864 478264
rect 193916 478252 193922 478304
rect 209590 478252 209596 478304
rect 209648 478292 209654 478304
rect 221734 478292 221740 478304
rect 209648 478264 221740 478292
rect 209648 478252 209654 478264
rect 221734 478252 221740 478264
rect 221792 478252 221798 478304
rect 230566 478252 230572 478304
rect 230624 478292 230630 478304
rect 366358 478292 366364 478304
rect 230624 478264 366364 478292
rect 230624 478252 230630 478264
rect 366358 478252 366364 478264
rect 366416 478252 366422 478304
rect 47946 478184 47952 478236
rect 48004 478224 48010 478236
rect 97166 478224 97172 478236
rect 48004 478196 97172 478224
rect 48004 478184 48010 478196
rect 97166 478184 97172 478196
rect 97224 478184 97230 478236
rect 109862 478184 109868 478236
rect 109920 478224 109926 478236
rect 169018 478224 169024 478236
rect 109920 478196 169024 478224
rect 109920 478184 109926 478196
rect 169018 478184 169024 478196
rect 169076 478184 169082 478236
rect 200206 478184 200212 478236
rect 200264 478224 200270 478236
rect 212258 478224 212264 478236
rect 200264 478196 212264 478224
rect 200264 478184 200270 478196
rect 212258 478184 212264 478196
rect 212316 478184 212322 478236
rect 225322 478184 225328 478236
rect 225380 478224 225386 478236
rect 362218 478224 362224 478236
rect 225380 478196 362224 478224
rect 225380 478184 225386 478196
rect 362218 478184 362224 478196
rect 362276 478184 362282 478236
rect 55122 478116 55128 478168
rect 55180 478156 55186 478168
rect 89622 478156 89628 478168
rect 55180 478128 89628 478156
rect 55180 478116 55186 478128
rect 89622 478116 89628 478128
rect 89680 478116 89686 478168
rect 95326 478116 95332 478168
rect 95384 478156 95390 478168
rect 182818 478156 182824 478168
rect 95384 478128 182824 478156
rect 95384 478116 95390 478128
rect 182818 478116 182824 478128
rect 182876 478116 182882 478168
rect 186498 478116 186504 478168
rect 186556 478156 186562 478168
rect 198182 478156 198188 478168
rect 186556 478128 198188 478156
rect 186556 478116 186562 478128
rect 198182 478116 198188 478128
rect 198240 478116 198246 478168
rect 201954 478116 201960 478168
rect 202012 478156 202018 478168
rect 217318 478156 217324 478168
rect 202012 478128 217324 478156
rect 202012 478116 202018 478128
rect 217318 478116 217324 478128
rect 217376 478116 217382 478168
rect 225690 478116 225696 478168
rect 225748 478156 225754 478168
rect 373258 478156 373264 478168
rect 225748 478128 373264 478156
rect 225748 478116 225754 478128
rect 373258 478116 373264 478128
rect 373316 478116 373322 478168
rect 64138 478048 64144 478100
rect 64196 478088 64202 478100
rect 69658 478088 69664 478100
rect 64196 478060 69664 478088
rect 64196 478048 64202 478060
rect 69658 478048 69664 478060
rect 69716 478048 69722 478100
rect 75270 478048 75276 478100
rect 75328 478088 75334 478100
rect 102870 478088 102876 478100
rect 75328 478060 102876 478088
rect 75328 478048 75334 478060
rect 102870 478048 102876 478060
rect 102928 478048 102934 478100
rect 150434 478048 150440 478100
rect 150492 478088 150498 478100
rect 197446 478088 197452 478100
rect 150492 478060 197452 478088
rect 150492 478048 150498 478060
rect 197446 478048 197452 478060
rect 197504 478048 197510 478100
rect 56502 477980 56508 478032
rect 56560 478020 56566 478032
rect 81710 478020 81716 478032
rect 56560 477992 81716 478020
rect 56560 477980 56566 477992
rect 81710 477980 81716 477992
rect 81768 477980 81774 478032
rect 156598 477980 156604 478032
rect 156656 478020 156662 478032
rect 197354 478020 197360 478032
rect 156656 477992 197360 478020
rect 156656 477980 156662 477992
rect 197354 477980 197360 477992
rect 197412 477980 197418 478032
rect 50890 477912 50896 477964
rect 50948 477952 50954 477964
rect 75822 477952 75828 477964
rect 50948 477924 75828 477952
rect 50948 477912 50954 477924
rect 75822 477912 75828 477924
rect 75880 477912 75886 477964
rect 139394 477912 139400 477964
rect 139452 477952 139458 477964
rect 178586 477952 178592 477964
rect 139452 477924 178592 477952
rect 139452 477912 139458 477924
rect 178586 477912 178592 477924
rect 178644 477912 178650 477964
rect 58434 477844 58440 477896
rect 58492 477884 58498 477896
rect 81250 477884 81256 477896
rect 58492 477856 81256 477884
rect 58492 477844 58498 477856
rect 81250 477844 81256 477856
rect 81308 477844 81314 477896
rect 168926 477844 168932 477896
rect 168984 477884 168990 477896
rect 206370 477884 206376 477896
rect 168984 477856 206376 477884
rect 168984 477844 168990 477856
rect 206370 477844 206376 477856
rect 206428 477844 206434 477896
rect 194870 477572 194876 477624
rect 194928 477612 194934 477624
rect 196986 477612 196992 477624
rect 194928 477584 196992 477612
rect 194928 477572 194934 477584
rect 196986 477572 196992 477584
rect 197044 477572 197050 477624
rect 202414 477572 202420 477624
rect 202472 477612 202478 477624
rect 209498 477612 209504 477624
rect 202472 477584 209504 477612
rect 202472 477572 202478 477584
rect 209498 477572 209504 477584
rect 209556 477572 209562 477624
rect 195790 477504 195796 477556
rect 195848 477544 195854 477556
rect 196894 477544 196900 477556
rect 195848 477516 196900 477544
rect 195848 477504 195854 477516
rect 196894 477504 196900 477516
rect 196952 477504 196958 477556
rect 208578 477504 208584 477556
rect 208636 477544 208642 477556
rect 210786 477544 210792 477556
rect 208636 477516 210792 477544
rect 208636 477504 208642 477516
rect 210786 477504 210792 477516
rect 210844 477504 210850 477556
rect 211154 477504 211160 477556
rect 211212 477544 211218 477556
rect 214558 477544 214564 477556
rect 211212 477516 214564 477544
rect 211212 477504 211218 477516
rect 214558 477504 214564 477516
rect 214616 477504 214622 477556
rect 220170 477504 220176 477556
rect 220228 477544 220234 477556
rect 222654 477544 222660 477556
rect 220228 477516 222660 477544
rect 220228 477504 220234 477516
rect 222654 477504 222660 477516
rect 222712 477504 222718 477556
rect 297082 477368 297088 477420
rect 297140 477408 297146 477420
rect 372522 477408 372528 477420
rect 297140 477380 372528 477408
rect 297140 477368 297146 477380
rect 372522 477368 372528 477380
rect 372580 477368 372586 477420
rect 290918 477300 290924 477352
rect 290976 477340 290982 477352
rect 365622 477340 365628 477352
rect 290976 477312 365628 477340
rect 290976 477300 290982 477312
rect 365622 477300 365628 477312
rect 365680 477300 365686 477352
rect 283006 477232 283012 477284
rect 283064 477272 283070 477284
rect 359734 477272 359740 477284
rect 283064 477244 359740 477272
rect 283064 477232 283070 477244
rect 359734 477232 359740 477244
rect 359792 477232 359798 477284
rect 282546 477164 282552 477216
rect 282604 477204 282610 477216
rect 363506 477204 363512 477216
rect 282604 477176 363512 477204
rect 282604 477164 282610 477176
rect 363506 477164 363512 477176
rect 363564 477164 363570 477216
rect 261846 477096 261852 477148
rect 261904 477136 261910 477148
rect 374178 477136 374184 477148
rect 261904 477108 374184 477136
rect 261904 477096 261910 477108
rect 374178 477096 374184 477108
rect 374236 477096 374242 477148
rect 256602 477028 256608 477080
rect 256660 477068 256666 477080
rect 376386 477068 376392 477080
rect 256660 477040 376392 477068
rect 256660 477028 256666 477040
rect 376386 477028 376392 477040
rect 376444 477028 376450 477080
rect 242894 476960 242900 477012
rect 242952 477000 242958 477012
rect 368014 477000 368020 477012
rect 242952 476972 368020 477000
rect 242952 476960 242958 476972
rect 368014 476960 368020 476972
rect 368072 476960 368078 477012
rect 45462 476892 45468 476944
rect 45520 476932 45526 476944
rect 117866 476932 117872 476944
rect 45520 476904 117872 476932
rect 45520 476892 45526 476904
rect 117866 476892 117872 476904
rect 117924 476892 117930 476944
rect 177758 476892 177764 476944
rect 177816 476932 177822 476944
rect 211982 476932 211988 476944
rect 177816 476904 211988 476932
rect 177816 476892 177822 476904
rect 211982 476892 211988 476904
rect 212040 476892 212046 476944
rect 247310 476892 247316 476944
rect 247368 476932 247374 476944
rect 374730 476932 374736 476944
rect 247368 476904 374736 476932
rect 247368 476892 247374 476904
rect 374730 476892 374736 476904
rect 374788 476892 374794 476944
rect 60550 476824 60556 476876
rect 60608 476864 60614 476876
rect 120718 476864 120724 476876
rect 60608 476836 120724 476864
rect 60608 476824 60614 476836
rect 120718 476824 120724 476836
rect 120776 476824 120782 476876
rect 120828 476836 125594 476864
rect 3602 476756 3608 476808
rect 3660 476796 3666 476808
rect 120828 476796 120856 476836
rect 3660 476768 120856 476796
rect 125566 476796 125594 476836
rect 159634 476824 159640 476876
rect 159692 476864 159698 476876
rect 218698 476864 218704 476876
rect 159692 476836 218704 476864
rect 159692 476824 159698 476836
rect 218698 476824 218704 476836
rect 218756 476824 218762 476876
rect 236730 476824 236736 476876
rect 236788 476864 236794 476876
rect 364978 476864 364984 476876
rect 236788 476836 364984 476864
rect 236788 476824 236794 476836
rect 364978 476824 364984 476836
rect 365036 476824 365042 476876
rect 429378 476796 429384 476808
rect 125566 476768 429384 476796
rect 3660 476756 3666 476768
rect 429378 476756 429384 476768
rect 429436 476756 429442 476808
rect 120718 476688 120724 476740
rect 120776 476728 120782 476740
rect 120776 476700 128354 476728
rect 120776 476688 120782 476700
rect 128326 476660 128354 476700
rect 133138 476660 133144 476672
rect 128326 476632 133144 476660
rect 133138 476620 133144 476632
rect 133196 476620 133202 476672
rect 70394 476076 70400 476128
rect 70452 476116 70458 476128
rect 70854 476116 70860 476128
rect 70452 476088 70860 476116
rect 70452 476076 70458 476088
rect 70854 476076 70860 476088
rect 70912 476076 70918 476128
rect 85758 476076 85764 476128
rect 85816 476116 85822 476128
rect 85942 476116 85948 476128
rect 85816 476088 85948 476116
rect 85816 476076 85822 476088
rect 85942 476076 85948 476088
rect 86000 476076 86006 476128
rect 47762 476008 47768 476060
rect 47820 476048 47826 476060
rect 111702 476048 111708 476060
rect 47820 476020 111708 476048
rect 47820 476008 47826 476020
rect 111702 476008 111708 476020
rect 111760 476008 111766 476060
rect 46658 475940 46664 475992
rect 46716 475980 46722 475992
rect 111242 475980 111248 475992
rect 46716 475952 111248 475980
rect 46716 475940 46722 475952
rect 111242 475940 111248 475952
rect 111300 475940 111306 475992
rect 294046 475940 294052 475992
rect 294104 475980 294110 475992
rect 294230 475980 294236 475992
rect 294104 475952 294236 475980
rect 294104 475940 294110 475952
rect 294230 475940 294236 475952
rect 294288 475940 294294 475992
rect 49234 475872 49240 475924
rect 49292 475912 49298 475924
rect 115198 475912 115204 475924
rect 49292 475884 115204 475912
rect 49292 475872 49298 475884
rect 115198 475872 115204 475884
rect 115256 475872 115262 475924
rect 274726 475872 274732 475924
rect 274784 475912 274790 475924
rect 274910 475912 274916 475924
rect 274784 475884 274916 475912
rect 274784 475872 274790 475884
rect 274910 475872 274916 475884
rect 274968 475872 274974 475924
rect 291838 475872 291844 475924
rect 291896 475912 291902 475924
rect 373902 475912 373908 475924
rect 291896 475884 373908 475912
rect 291896 475872 291902 475884
rect 373902 475872 373908 475884
rect 373960 475872 373966 475924
rect 46382 475804 46388 475856
rect 46440 475844 46446 475856
rect 112530 475844 112536 475856
rect 46440 475816 112536 475844
rect 46440 475804 46446 475816
rect 112530 475804 112536 475816
rect 112588 475804 112594 475856
rect 267550 475804 267556 475856
rect 267608 475844 267614 475856
rect 359458 475844 359464 475856
rect 267608 475816 359464 475844
rect 267608 475804 267614 475816
rect 359458 475804 359464 475816
rect 359516 475804 359522 475856
rect 46474 475736 46480 475788
rect 46532 475776 46538 475788
rect 112070 475776 112076 475788
rect 46532 475748 112076 475776
rect 46532 475736 46538 475748
rect 112070 475736 112076 475748
rect 112128 475736 112134 475788
rect 267090 475736 267096 475788
rect 267148 475776 267154 475788
rect 359550 475776 359556 475788
rect 267148 475748 359556 475776
rect 267148 475736 267154 475748
rect 359550 475736 359556 475748
rect 359608 475736 359614 475788
rect 50246 475668 50252 475720
rect 50304 475708 50310 475720
rect 116026 475708 116032 475720
rect 50304 475680 116032 475708
rect 50304 475668 50310 475680
rect 116026 475668 116032 475680
rect 116084 475668 116090 475720
rect 136358 475668 136364 475720
rect 136416 475708 136422 475720
rect 141878 475708 141884 475720
rect 136416 475680 141884 475708
rect 136416 475668 136422 475680
rect 141878 475668 141884 475680
rect 141936 475668 141942 475720
rect 171134 475668 171140 475720
rect 171192 475708 171198 475720
rect 171318 475708 171324 475720
rect 171192 475680 171324 475708
rect 171192 475668 171198 475680
rect 171318 475668 171324 475680
rect 171376 475668 171382 475720
rect 184290 475668 184296 475720
rect 184348 475708 184354 475720
rect 216122 475708 216128 475720
rect 184348 475680 216128 475708
rect 184348 475668 184354 475680
rect 216122 475668 216128 475680
rect 216180 475668 216186 475720
rect 273254 475668 273260 475720
rect 273312 475708 273318 475720
rect 369762 475708 369768 475720
rect 273312 475680 369768 475708
rect 273312 475668 273318 475680
rect 369762 475668 369768 475680
rect 369820 475668 369826 475720
rect 48130 475600 48136 475652
rect 48188 475640 48194 475652
rect 115658 475640 115664 475652
rect 48188 475612 115664 475640
rect 48188 475600 48194 475612
rect 115658 475600 115664 475612
rect 115716 475600 115722 475652
rect 138106 475600 138112 475652
rect 138164 475640 138170 475652
rect 200482 475640 200488 475652
rect 138164 475612 200488 475640
rect 138164 475600 138170 475612
rect 200482 475600 200488 475612
rect 200540 475600 200546 475652
rect 219526 475600 219532 475652
rect 219584 475600 219590 475652
rect 272886 475600 272892 475652
rect 272944 475640 272950 475652
rect 372430 475640 372436 475652
rect 272944 475612 372436 475640
rect 272944 475600 272950 475612
rect 372430 475600 372436 475612
rect 372488 475600 372494 475652
rect 47854 475532 47860 475584
rect 47912 475572 47918 475584
rect 119614 475572 119620 475584
rect 47912 475544 119620 475572
rect 47912 475532 47918 475544
rect 119614 475532 119620 475544
rect 119672 475532 119678 475584
rect 136726 475532 136732 475584
rect 136784 475572 136790 475584
rect 199378 475572 199384 475584
rect 136784 475544 199384 475572
rect 136784 475532 136790 475544
rect 199378 475532 199384 475544
rect 199436 475532 199442 475584
rect 57146 475464 57152 475516
rect 57204 475504 57210 475516
rect 132402 475504 132408 475516
rect 57204 475476 132408 475504
rect 57204 475464 57210 475476
rect 132402 475464 132408 475476
rect 132460 475464 132466 475516
rect 137646 475464 137652 475516
rect 137704 475504 137710 475516
rect 137704 475476 141832 475504
rect 137704 475464 137710 475476
rect 57330 475396 57336 475448
rect 57388 475436 57394 475448
rect 135898 475436 135904 475448
rect 57388 475408 135904 475436
rect 57388 475396 57394 475408
rect 135898 475396 135904 475408
rect 135956 475396 135962 475448
rect 140774 475396 140780 475448
rect 140832 475436 140838 475448
rect 141694 475436 141700 475448
rect 140832 475408 141700 475436
rect 140832 475396 140838 475408
rect 141694 475396 141700 475408
rect 141752 475396 141758 475448
rect 141804 475436 141832 475476
rect 141878 475464 141884 475516
rect 141936 475504 141942 475516
rect 201678 475504 201684 475516
rect 141936 475476 201684 475504
rect 141936 475464 141942 475476
rect 201678 475464 201684 475476
rect 201736 475464 201742 475516
rect 212534 475504 212540 475516
rect 212460 475476 212540 475504
rect 204438 475436 204444 475448
rect 141804 475408 204444 475436
rect 204438 475396 204444 475408
rect 204496 475396 204502 475448
rect 62114 475328 62120 475380
rect 62172 475368 62178 475380
rect 62942 475368 62948 475380
rect 62172 475340 62948 475368
rect 62172 475328 62178 475340
rect 62942 475328 62948 475340
rect 63000 475328 63006 475380
rect 63494 475328 63500 475380
rect 63552 475368 63558 475380
rect 64230 475368 64236 475380
rect 63552 475340 64236 475368
rect 63552 475328 63558 475340
rect 64230 475328 64236 475340
rect 64288 475328 64294 475380
rect 64322 475328 64328 475380
rect 64380 475368 64386 475380
rect 64380 475340 186314 475368
rect 64380 475328 64386 475340
rect 49142 475260 49148 475312
rect 49200 475300 49206 475312
rect 97994 475300 98000 475312
rect 49200 475272 98000 475300
rect 49200 475260 49206 475272
rect 97994 475260 98000 475272
rect 98052 475260 98058 475312
rect 100846 475260 100852 475312
rect 100904 475300 100910 475312
rect 101214 475300 101220 475312
rect 100904 475272 101220 475300
rect 100904 475260 100910 475272
rect 101214 475260 101220 475272
rect 101272 475260 101278 475312
rect 103606 475260 103612 475312
rect 103664 475300 103670 475312
rect 103790 475300 103796 475312
rect 103664 475272 103796 475300
rect 103664 475260 103670 475272
rect 103790 475260 103796 475272
rect 103848 475260 103854 475312
rect 107654 475260 107660 475312
rect 107712 475300 107718 475312
rect 107838 475300 107844 475312
rect 107712 475272 107844 475300
rect 107712 475260 107718 475272
rect 107838 475260 107844 475272
rect 107896 475260 107902 475312
rect 133966 475260 133972 475312
rect 134024 475300 134030 475312
rect 134702 475300 134708 475312
rect 134024 475272 134708 475300
rect 134024 475260 134030 475272
rect 134702 475260 134708 475272
rect 134760 475260 134766 475312
rect 139394 475260 139400 475312
rect 139452 475300 139458 475312
rect 140038 475300 140044 475312
rect 139452 475272 140044 475300
rect 139452 475260 139458 475272
rect 140038 475260 140044 475272
rect 140096 475260 140102 475312
rect 140866 475260 140872 475312
rect 140924 475300 140930 475312
rect 141326 475300 141332 475312
rect 140924 475272 141332 475300
rect 140924 475260 140930 475272
rect 141326 475260 141332 475272
rect 141384 475260 141390 475312
rect 142246 475260 142252 475312
rect 142304 475300 142310 475312
rect 142614 475300 142620 475312
rect 142304 475272 142620 475300
rect 142304 475260 142310 475272
rect 142614 475260 142620 475272
rect 142672 475260 142678 475312
rect 143534 475260 143540 475312
rect 143592 475300 143598 475312
rect 143902 475300 143908 475312
rect 143592 475272 143908 475300
rect 143592 475260 143598 475272
rect 143902 475260 143908 475272
rect 143960 475260 143966 475312
rect 150434 475260 150440 475312
rect 150492 475300 150498 475312
rect 151446 475300 151452 475312
rect 150492 475272 151452 475300
rect 150492 475260 150498 475272
rect 151446 475260 151452 475272
rect 151504 475260 151510 475312
rect 160094 475260 160100 475312
rect 160152 475300 160158 475312
rect 160646 475300 160652 475312
rect 160152 475272 160652 475300
rect 160152 475260 160158 475272
rect 160646 475260 160652 475272
rect 160704 475260 160710 475312
rect 161566 475260 161572 475312
rect 161624 475300 161630 475312
rect 161934 475300 161940 475312
rect 161624 475272 161940 475300
rect 161624 475260 161630 475272
rect 161934 475260 161940 475272
rect 161992 475260 161998 475312
rect 165614 475260 165620 475312
rect 165672 475300 165678 475312
rect 166350 475300 166356 475312
rect 165672 475272 166356 475300
rect 165672 475260 165678 475272
rect 166350 475260 166356 475272
rect 166408 475260 166414 475312
rect 166994 475260 167000 475312
rect 167052 475300 167058 475312
rect 167730 475300 167736 475312
rect 167052 475272 167736 475300
rect 167052 475260 167058 475272
rect 167730 475260 167736 475272
rect 167788 475260 167794 475312
rect 178126 475260 178132 475312
rect 178184 475300 178190 475312
rect 178678 475300 178684 475312
rect 178184 475272 178684 475300
rect 178184 475260 178190 475272
rect 178678 475260 178684 475272
rect 178736 475260 178742 475312
rect 179414 475260 179420 475312
rect 179472 475300 179478 475312
rect 180058 475300 180064 475312
rect 179472 475272 180064 475300
rect 179472 475260 179478 475272
rect 180058 475260 180064 475272
rect 180116 475260 180122 475312
rect 180886 475260 180892 475312
rect 180944 475300 180950 475312
rect 181438 475300 181444 475312
rect 180944 475272 181444 475300
rect 180944 475260 180950 475272
rect 181438 475260 181444 475272
rect 181496 475260 181502 475312
rect 182358 475260 182364 475312
rect 182416 475300 182422 475312
rect 182726 475300 182732 475312
rect 182416 475272 182732 475300
rect 182416 475260 182422 475272
rect 182726 475260 182732 475272
rect 182784 475260 182790 475312
rect 183554 475260 183560 475312
rect 183612 475300 183618 475312
rect 184382 475300 184388 475312
rect 183612 475272 184388 475300
rect 183612 475260 183618 475272
rect 184382 475260 184388 475272
rect 184440 475260 184446 475312
rect 185026 475260 185032 475312
rect 185084 475300 185090 475312
rect 185854 475300 185860 475312
rect 185084 475272 185860 475300
rect 185084 475260 185090 475272
rect 185854 475260 185860 475272
rect 185912 475260 185918 475312
rect 51810 475192 51816 475244
rect 51868 475232 51874 475244
rect 98454 475232 98460 475244
rect 51868 475204 98460 475232
rect 51868 475192 51874 475204
rect 98454 475192 98460 475204
rect 98512 475192 98518 475244
rect 100754 475192 100760 475244
rect 100812 475232 100818 475244
rect 101582 475232 101588 475244
rect 100812 475204 101588 475232
rect 100812 475192 100818 475204
rect 101582 475192 101588 475204
rect 101640 475192 101646 475244
rect 142154 475192 142160 475244
rect 142212 475232 142218 475244
rect 142982 475232 142988 475244
rect 142212 475204 142988 475232
rect 142212 475192 142218 475204
rect 142982 475192 142988 475204
rect 143040 475192 143046 475244
rect 161474 475192 161480 475244
rect 161532 475232 161538 475244
rect 161750 475232 161756 475244
rect 161532 475204 161756 475232
rect 161532 475192 161538 475204
rect 161750 475192 161756 475204
rect 161808 475192 161814 475244
rect 180794 475192 180800 475244
rect 180852 475232 180858 475244
rect 181070 475232 181076 475244
rect 180852 475204 181076 475232
rect 180852 475192 180858 475204
rect 181070 475192 181076 475204
rect 181128 475192 181134 475244
rect 182174 475192 182180 475244
rect 182232 475232 182238 475244
rect 182542 475232 182548 475244
rect 182232 475204 182548 475232
rect 182232 475192 182238 475204
rect 182542 475192 182548 475204
rect 182600 475192 182606 475244
rect 186286 475232 186314 475340
rect 205726 475328 205732 475380
rect 205784 475368 205790 475380
rect 206462 475368 206468 475380
rect 205784 475340 206468 475368
rect 205784 475328 205790 475340
rect 206462 475328 206468 475340
rect 206520 475328 206526 475380
rect 207198 475328 207204 475380
rect 207256 475368 207262 475380
rect 207750 475368 207756 475380
rect 207256 475340 207756 475368
rect 207256 475328 207262 475340
rect 207750 475328 207756 475340
rect 207808 475328 207814 475380
rect 209774 475328 209780 475380
rect 209832 475368 209838 475380
rect 209958 475368 209964 475380
rect 209832 475340 209964 475368
rect 209832 475328 209838 475340
rect 209958 475328 209964 475340
rect 210016 475328 210022 475380
rect 212460 475300 212488 475476
rect 212534 475464 212540 475476
rect 212592 475464 212598 475516
rect 219544 475448 219572 475600
rect 253014 475532 253020 475584
rect 253072 475572 253078 475584
rect 365438 475572 365444 475584
rect 253072 475544 365444 475572
rect 253072 475532 253078 475544
rect 365438 475532 365444 475544
rect 365496 475532 365502 475584
rect 243354 475464 243360 475516
rect 243412 475504 243418 475516
rect 369210 475504 369216 475516
rect 243412 475476 369216 475504
rect 243412 475464 243418 475476
rect 369210 475464 369216 475476
rect 369268 475464 369274 475516
rect 219526 475396 219532 475448
rect 219584 475396 219590 475448
rect 247770 475396 247776 475448
rect 247828 475436 247834 475448
rect 376202 475436 376208 475448
rect 247828 475408 376208 475436
rect 247828 475396 247834 475408
rect 376202 475396 376208 475408
rect 376260 475396 376266 475448
rect 212534 475328 212540 475380
rect 212592 475368 212598 475380
rect 213086 475368 213092 475380
rect 212592 475340 213092 475368
rect 212592 475328 212598 475340
rect 213086 475328 213092 475340
rect 213144 475328 213150 475380
rect 213914 475328 213920 475380
rect 213972 475368 213978 475380
rect 214926 475368 214932 475380
rect 213972 475340 214932 475368
rect 213972 475328 213978 475340
rect 214926 475328 214932 475340
rect 214984 475328 214990 475380
rect 215294 475328 215300 475380
rect 215352 475368 215358 475380
rect 216214 475368 216220 475380
rect 215352 475340 216220 475368
rect 215352 475328 215358 475340
rect 216214 475328 216220 475340
rect 216272 475328 216278 475380
rect 218054 475328 218060 475380
rect 218112 475368 218118 475380
rect 218790 475368 218796 475380
rect 218112 475340 218796 475368
rect 218112 475328 218118 475340
rect 218790 475328 218796 475340
rect 218848 475328 218854 475380
rect 222194 475328 222200 475380
rect 222252 475368 222258 475380
rect 374638 475368 374644 475380
rect 222252 475340 374644 475368
rect 222252 475328 222258 475340
rect 374638 475328 374644 475340
rect 374696 475328 374702 475380
rect 212718 475300 212724 475312
rect 212460 475272 212724 475300
rect 212718 475260 212724 475272
rect 212776 475260 212782 475312
rect 244274 475260 244280 475312
rect 244332 475300 244338 475312
rect 244550 475300 244556 475312
rect 244332 475272 244556 475300
rect 244332 475260 244338 475272
rect 244550 475260 244556 475272
rect 244608 475260 244614 475312
rect 245654 475260 245660 475312
rect 245712 475300 245718 475312
rect 246574 475300 246580 475312
rect 245712 475272 246580 475300
rect 245712 475260 245718 475272
rect 246574 475260 246580 475272
rect 246632 475260 246638 475312
rect 248506 475260 248512 475312
rect 248564 475300 248570 475312
rect 249150 475300 249156 475312
rect 248564 475272 249156 475300
rect 248564 475260 248570 475272
rect 249150 475260 249156 475272
rect 249208 475260 249214 475312
rect 251174 475260 251180 475312
rect 251232 475300 251238 475312
rect 251358 475300 251364 475312
rect 251232 475272 251364 475300
rect 251232 475260 251238 475272
rect 251358 475260 251364 475272
rect 251416 475260 251422 475312
rect 252554 475260 252560 475312
rect 252612 475300 252618 475312
rect 253198 475300 253204 475312
rect 252612 475272 253204 475300
rect 252612 475260 252618 475272
rect 253198 475260 253204 475272
rect 253256 475260 253262 475312
rect 259454 475260 259460 475312
rect 259512 475300 259518 475312
rect 260190 475300 260196 475312
rect 259512 475272 260196 475300
rect 259512 475260 259518 475272
rect 260190 475260 260196 475272
rect 260248 475260 260254 475312
rect 262214 475260 262220 475312
rect 262272 475300 262278 475312
rect 262398 475300 262404 475312
rect 262272 475272 262404 475300
rect 262272 475260 262278 475272
rect 262398 475260 262404 475272
rect 262456 475260 262462 475312
rect 276106 475260 276112 475312
rect 276164 475300 276170 475312
rect 276566 475300 276572 475312
rect 276164 475272 276572 475300
rect 276164 475260 276170 475272
rect 276566 475260 276572 475272
rect 276624 475260 276630 475312
rect 277486 475260 277492 475312
rect 277544 475300 277550 475312
rect 277854 475300 277860 475312
rect 277544 475272 277860 475300
rect 277544 475260 277550 475272
rect 277854 475260 277860 475272
rect 277912 475260 277918 475312
rect 284294 475260 284300 475312
rect 284352 475300 284358 475312
rect 284846 475300 284852 475312
rect 284352 475272 284852 475300
rect 284352 475260 284358 475272
rect 284846 475260 284852 475272
rect 284904 475260 284910 475312
rect 285674 475260 285680 475312
rect 285732 475300 285738 475312
rect 286686 475300 286692 475312
rect 285732 475272 286692 475300
rect 285732 475260 285738 475272
rect 286686 475260 286692 475272
rect 286744 475260 286750 475312
rect 291194 475260 291200 475312
rect 291252 475300 291258 475312
rect 291930 475300 291936 475312
rect 291252 475272 291936 475300
rect 291252 475260 291258 475272
rect 291930 475260 291936 475272
rect 291988 475260 291994 475312
rect 296714 475260 296720 475312
rect 296772 475300 296778 475312
rect 297726 475300 297732 475312
rect 296772 475272 297732 475300
rect 296772 475260 296778 475272
rect 297726 475260 297732 475272
rect 297784 475260 297790 475312
rect 199194 475232 199200 475244
rect 186286 475204 199200 475232
rect 199194 475192 199200 475204
rect 199252 475192 199258 475244
rect 276014 475192 276020 475244
rect 276072 475232 276078 475244
rect 276934 475232 276940 475244
rect 276072 475204 276940 475232
rect 276072 475192 276078 475204
rect 276934 475192 276940 475204
rect 276992 475192 276998 475244
rect 277394 475192 277400 475244
rect 277452 475232 277458 475244
rect 278222 475232 278228 475244
rect 277452 475204 278228 475232
rect 277452 475192 277458 475204
rect 278222 475192 278228 475204
rect 278280 475192 278286 475244
rect 54662 475124 54668 475176
rect 54720 475164 54726 475176
rect 96706 475164 96712 475176
rect 54720 475136 96712 475164
rect 54720 475124 54726 475136
rect 96706 475124 96712 475136
rect 96764 475124 96770 475176
rect 182266 475124 182272 475176
rect 182324 475164 182330 475176
rect 183094 475164 183100 475176
rect 182324 475136 183100 475164
rect 182324 475124 182330 475136
rect 183094 475124 183100 475136
rect 183152 475124 183158 475176
rect 205634 475124 205640 475176
rect 205692 475164 205698 475176
rect 205910 475164 205916 475176
rect 205692 475136 205916 475164
rect 205692 475124 205698 475136
rect 205910 475124 205916 475136
rect 205968 475124 205974 475176
rect 62758 475056 62764 475108
rect 62816 475096 62822 475108
rect 64322 475096 64328 475108
rect 62816 475068 64328 475096
rect 62816 475056 62822 475068
rect 64322 475056 64328 475068
rect 64380 475056 64386 475108
rect 64966 475056 64972 475108
rect 65024 475096 65030 475108
rect 65518 475096 65524 475108
rect 65024 475068 65524 475096
rect 65024 475056 65030 475068
rect 65518 475056 65524 475068
rect 65576 475056 65582 475108
rect 66254 475056 66260 475108
rect 66312 475096 66318 475108
rect 66806 475096 66812 475108
rect 66312 475068 66812 475096
rect 66312 475056 66318 475068
rect 66806 475056 66812 475068
rect 66864 475056 66870 475108
rect 71866 475056 71872 475108
rect 71924 475096 71930 475108
rect 72602 475096 72608 475108
rect 71924 475068 72608 475096
rect 71924 475056 71930 475068
rect 72602 475056 72608 475068
rect 72660 475056 72666 475108
rect 78674 475056 78680 475108
rect 78732 475096 78738 475108
rect 79686 475096 79692 475108
rect 78732 475068 79692 475096
rect 78732 475056 78738 475068
rect 79686 475056 79692 475068
rect 79744 475056 79750 475108
rect 82814 475056 82820 475108
rect 82872 475096 82878 475108
rect 83550 475096 83556 475108
rect 82872 475068 83556 475096
rect 82872 475056 82878 475068
rect 83550 475056 83556 475068
rect 83608 475056 83614 475108
rect 85666 475056 85672 475108
rect 85724 475096 85730 475108
rect 86310 475096 86316 475108
rect 85724 475068 86316 475096
rect 85724 475056 85730 475068
rect 86310 475056 86316 475068
rect 86368 475056 86374 475108
rect 87046 475056 87052 475108
rect 87104 475096 87110 475108
rect 87230 475096 87236 475108
rect 87104 475068 87236 475096
rect 87104 475056 87110 475068
rect 87230 475056 87236 475068
rect 87288 475056 87294 475108
rect 88426 475056 88432 475108
rect 88484 475096 88490 475108
rect 88886 475096 88892 475108
rect 88484 475068 88892 475096
rect 88484 475056 88490 475068
rect 88886 475056 88892 475068
rect 88944 475056 88950 475108
rect 89806 475056 89812 475108
rect 89864 475096 89870 475108
rect 90726 475096 90732 475108
rect 89864 475068 90732 475096
rect 89864 475056 89870 475068
rect 90726 475056 90732 475068
rect 90784 475056 90790 475108
rect 92474 475056 92480 475108
rect 92532 475096 92538 475108
rect 92934 475096 92940 475108
rect 92532 475068 92940 475096
rect 92532 475056 92538 475068
rect 92934 475056 92940 475068
rect 92992 475056 92998 475108
rect 86954 474988 86960 475040
rect 87012 475028 87018 475040
rect 87598 475028 87604 475040
rect 87012 475000 87604 475028
rect 87012 474988 87018 475000
rect 87598 474988 87604 475000
rect 87656 474988 87662 475040
rect 88518 474988 88524 475040
rect 88576 475028 88582 475040
rect 88702 475028 88708 475040
rect 88576 475000 88708 475028
rect 88576 474988 88582 475000
rect 88702 474988 88708 475000
rect 88760 474988 88766 475040
rect 92566 474988 92572 475040
rect 92624 475028 92630 475040
rect 93302 475028 93308 475040
rect 92624 475000 93308 475028
rect 92624 474988 92630 475000
rect 93302 474988 93308 475000
rect 93360 474988 93366 475040
rect 293586 474648 293592 474700
rect 293644 474688 293650 474700
rect 379330 474688 379336 474700
rect 293644 474660 379336 474688
rect 293644 474648 293650 474660
rect 379330 474648 379336 474660
rect 379388 474648 379394 474700
rect 282086 474580 282092 474632
rect 282144 474620 282150 474632
rect 379974 474620 379980 474632
rect 282144 474592 379980 474620
rect 282144 474580 282150 474592
rect 379974 474580 379980 474592
rect 380032 474580 380038 474632
rect 275922 474512 275928 474564
rect 275980 474552 275986 474564
rect 373718 474552 373724 474564
rect 275980 474524 373724 474552
rect 275980 474512 275986 474524
rect 373718 474512 373724 474524
rect 373776 474512 373782 474564
rect 260926 474444 260932 474496
rect 260984 474484 260990 474496
rect 362494 474484 362500 474496
rect 260984 474456 362500 474484
rect 260984 474444 260990 474456
rect 362494 474444 362500 474456
rect 362552 474444 362558 474496
rect 254762 474376 254768 474428
rect 254820 474416 254826 474428
rect 366818 474416 366824 474428
rect 254820 474388 366824 474416
rect 254820 474376 254826 474388
rect 366818 474376 366824 474388
rect 366876 474376 366882 474428
rect 255222 474308 255228 474360
rect 255280 474348 255286 474360
rect 369118 474348 369124 474360
rect 255280 474320 369124 474348
rect 255280 474308 255286 474320
rect 369118 474308 369124 474320
rect 369176 474308 369182 474360
rect 252186 474240 252192 474292
rect 252244 474280 252250 474292
rect 366910 474280 366916 474292
rect 252244 474252 366916 474280
rect 252244 474240 252250 474252
rect 366910 474240 366916 474252
rect 366968 474240 366974 474292
rect 242434 474172 242440 474224
rect 242492 474212 242498 474224
rect 370590 474212 370596 474224
rect 242492 474184 370596 474212
rect 242492 474172 242498 474184
rect 370590 474172 370596 474184
rect 370648 474172 370654 474224
rect 204990 474104 204996 474156
rect 205048 474144 205054 474156
rect 217318 474144 217324 474156
rect 205048 474116 217324 474144
rect 205048 474104 205054 474116
rect 217318 474104 217324 474116
rect 217376 474104 217382 474156
rect 228818 474104 228824 474156
rect 228876 474144 228882 474156
rect 363598 474144 363604 474156
rect 228876 474116 363604 474144
rect 228876 474104 228882 474116
rect 363598 474104 363604 474116
rect 363656 474104 363662 474156
rect 96246 474076 96252 474088
rect 84166 474048 96252 474076
rect 58802 473968 58808 474020
rect 58860 474008 58866 474020
rect 84166 474008 84194 474048
rect 96246 474036 96252 474048
rect 96304 474036 96310 474088
rect 176010 474036 176016 474088
rect 176068 474076 176074 474088
rect 210602 474076 210608 474088
rect 176068 474048 210608 474076
rect 176068 474036 176074 474048
rect 210602 474036 210608 474048
rect 210660 474036 210666 474088
rect 238110 474036 238116 474088
rect 238168 474076 238174 474088
rect 376294 474076 376300 474088
rect 238168 474048 376300 474076
rect 238168 474036 238174 474048
rect 376294 474036 376300 474048
rect 376352 474036 376358 474088
rect 58860 473980 84194 474008
rect 58860 473968 58866 473980
rect 166258 473968 166264 474020
rect 166316 474008 166322 474020
rect 215938 474008 215944 474020
rect 166316 473980 215944 474008
rect 166316 473968 166322 473980
rect 215938 473968 215944 473980
rect 215996 473968 216002 474020
rect 228358 473968 228364 474020
rect 228416 474008 228422 474020
rect 367830 474008 367836 474020
rect 228416 473980 367836 474008
rect 228416 473968 228422 473980
rect 367830 473968 367836 473980
rect 367888 473968 367894 474020
rect 295334 473900 295340 473952
rect 295392 473940 295398 473952
rect 375466 473940 375472 473952
rect 295392 473912 375472 473940
rect 295392 473900 295398 473912
rect 375466 473900 375472 473912
rect 375524 473900 375530 473952
rect 81526 473560 81532 473612
rect 81584 473600 81590 473612
rect 82262 473600 82268 473612
rect 81584 473572 82268 473600
rect 81584 473560 81590 473572
rect 82262 473560 82268 473572
rect 82320 473560 82326 473612
rect 46842 473288 46848 473340
rect 46900 473328 46906 473340
rect 116486 473328 116492 473340
rect 46900 473300 116492 473328
rect 46900 473288 46906 473300
rect 116486 473288 116492 473300
rect 116544 473288 116550 473340
rect 58618 473220 58624 473272
rect 58676 473260 58682 473272
rect 130562 473260 130568 473272
rect 58676 473232 130568 473260
rect 58676 473220 58682 473232
rect 130562 473220 130568 473232
rect 130620 473220 130626 473272
rect 59722 473152 59728 473204
rect 59780 473192 59786 473204
rect 132586 473192 132592 473204
rect 59780 473164 132592 473192
rect 59780 473152 59786 473164
rect 132586 473152 132592 473164
rect 132644 473152 132650 473204
rect 43990 473084 43996 473136
rect 44048 473124 44054 473136
rect 118234 473124 118240 473136
rect 44048 473096 118240 473124
rect 44048 473084 44054 473096
rect 118234 473084 118240 473096
rect 118292 473084 118298 473136
rect 298554 473084 298560 473136
rect 298612 473124 298618 473136
rect 373994 473124 374000 473136
rect 298612 473096 374000 473124
rect 298612 473084 298618 473096
rect 373994 473084 374000 473096
rect 374052 473084 374058 473136
rect 49050 473016 49056 473068
rect 49108 473056 49114 473068
rect 131022 473056 131028 473068
rect 49108 473028 131028 473056
rect 49108 473016 49114 473028
rect 131022 473016 131028 473028
rect 131080 473016 131086 473068
rect 275462 473016 275468 473068
rect 275520 473056 275526 473068
rect 356882 473056 356888 473068
rect 275520 473028 356888 473056
rect 275520 473016 275526 473028
rect 356882 473016 356888 473028
rect 356940 473016 356946 473068
rect 50154 472948 50160 473000
rect 50212 472988 50218 473000
rect 131482 472988 131488 473000
rect 50212 472960 131488 472988
rect 50212 472948 50218 472960
rect 131482 472948 131488 472960
rect 131540 472948 131546 473000
rect 295794 472948 295800 473000
rect 295852 472988 295858 473000
rect 377766 472988 377772 473000
rect 295852 472960 377772 472988
rect 295852 472948 295858 472960
rect 377766 472948 377772 472960
rect 377824 472948 377830 473000
rect 52270 472880 52276 472932
rect 52328 472920 52334 472932
rect 134150 472920 134156 472932
rect 52328 472892 134156 472920
rect 52328 472880 52334 472892
rect 134150 472880 134156 472892
rect 134208 472880 134214 472932
rect 279234 472880 279240 472932
rect 279292 472920 279298 472932
rect 364886 472920 364892 472932
rect 279292 472892 364892 472920
rect 279292 472880 279298 472892
rect 364886 472880 364892 472892
rect 364944 472880 364950 472932
rect 47578 472812 47584 472864
rect 47636 472852 47642 472864
rect 129734 472852 129740 472864
rect 47636 472824 129740 472852
rect 47636 472812 47642 472824
rect 129734 472812 129740 472824
rect 129792 472812 129798 472864
rect 280798 472812 280804 472864
rect 280856 472852 280862 472864
rect 369670 472852 369676 472864
rect 280856 472824 369676 472852
rect 280856 472812 280862 472824
rect 369670 472812 369676 472824
rect 369728 472812 369734 472864
rect 46106 472744 46112 472796
rect 46164 472784 46170 472796
rect 129274 472784 129280 472796
rect 46164 472756 129280 472784
rect 46164 472744 46170 472756
rect 129274 472744 129280 472756
rect 129332 472744 129338 472796
rect 258810 472744 258816 472796
rect 258868 472784 258874 472796
rect 372246 472784 372252 472796
rect 258868 472756 372252 472784
rect 258868 472744 258874 472756
rect 372246 472744 372252 472756
rect 372304 472744 372310 472796
rect 42334 472676 42340 472728
rect 42392 472716 42398 472728
rect 131942 472716 131948 472728
rect 42392 472688 131948 472716
rect 42392 472676 42398 472688
rect 131942 472676 131948 472688
rect 132000 472676 132006 472728
rect 238478 472676 238484 472728
rect 238536 472716 238542 472728
rect 358078 472716 358084 472728
rect 238536 472688 358084 472716
rect 238536 472676 238542 472688
rect 358078 472676 358084 472688
rect 358136 472676 358142 472728
rect 43254 472608 43260 472660
rect 43312 472648 43318 472660
rect 132494 472648 132500 472660
rect 43312 472620 132500 472648
rect 43312 472608 43318 472620
rect 132494 472608 132500 472620
rect 132552 472608 132558 472660
rect 175550 472608 175556 472660
rect 175608 472648 175614 472660
rect 213178 472648 213184 472660
rect 175608 472620 213184 472648
rect 175608 472608 175614 472620
rect 213178 472608 213184 472620
rect 213236 472608 213242 472660
rect 239398 472608 239404 472660
rect 239456 472648 239462 472660
rect 378778 472648 378784 472660
rect 239456 472620 378784 472648
rect 239456 472608 239462 472620
rect 378778 472608 378784 472620
rect 378836 472608 378842 472660
rect 47670 472540 47676 472592
rect 47728 472580 47734 472592
rect 116946 472580 116952 472592
rect 47728 472552 116952 472580
rect 47728 472540 47734 472552
rect 116946 472540 116952 472552
rect 117004 472540 117010 472592
rect 54570 472472 54576 472524
rect 54628 472512 54634 472524
rect 117406 472512 117412 472524
rect 54628 472484 117412 472512
rect 54628 472472 54634 472484
rect 117406 472472 117412 472484
rect 117464 472472 117470 472524
rect 172514 472472 172520 472524
rect 172572 472512 172578 472524
rect 173526 472512 173532 472524
rect 172572 472484 173532 472512
rect 172572 472472 172578 472484
rect 173526 472472 173532 472484
rect 173584 472472 173590 472524
rect 57882 472404 57888 472456
rect 57940 472444 57946 472456
rect 114278 472444 114284 472456
rect 57940 472416 114284 472444
rect 57940 472404 57946 472416
rect 114278 472404 114284 472416
rect 114336 472404 114342 472456
rect 296162 471928 296168 471980
rect 296220 471968 296226 471980
rect 373810 471968 373816 471980
rect 296220 471940 373816 471968
rect 296220 471928 296226 471940
rect 373810 471928 373816 471940
rect 373868 471928 373874 471980
rect 288710 471860 288716 471912
rect 288768 471900 288774 471912
rect 375190 471900 375196 471912
rect 288768 471872 375196 471900
rect 288768 471860 288774 471872
rect 375190 471860 375196 471872
rect 375248 471860 375254 471912
rect 270678 471792 270684 471844
rect 270736 471832 270742 471844
rect 358446 471832 358452 471844
rect 270736 471804 358452 471832
rect 270736 471792 270742 471804
rect 358446 471792 358452 471804
rect 358504 471792 358510 471844
rect 272426 471724 272432 471776
rect 272484 471764 272490 471776
rect 360746 471764 360752 471776
rect 272484 471736 360752 471764
rect 272484 471724 272490 471736
rect 360746 471724 360752 471736
rect 360804 471724 360810 471776
rect 266262 471656 266268 471708
rect 266320 471696 266326 471708
rect 356790 471696 356796 471708
rect 266320 471668 356796 471696
rect 266320 471656 266326 471668
rect 356790 471656 356796 471668
rect 356848 471656 356854 471708
rect 265802 471588 265808 471640
rect 265860 471628 265866 471640
rect 361022 471628 361028 471640
rect 265860 471600 361028 471628
rect 265860 471588 265866 471600
rect 361022 471588 361028 471600
rect 361080 471588 361086 471640
rect 257430 471520 257436 471572
rect 257488 471560 257494 471572
rect 358354 471560 358360 471572
rect 257488 471532 358360 471560
rect 257488 471520 257494 471532
rect 358354 471520 358360 471532
rect 358412 471520 358418 471572
rect 259638 471452 259644 471504
rect 259696 471492 259702 471504
rect 369486 471492 369492 471504
rect 259696 471464 369492 471492
rect 259696 471452 259702 471464
rect 369486 471452 369492 471464
rect 369544 471452 369550 471504
rect 253934 471384 253940 471436
rect 253992 471424 253998 471436
rect 369578 471424 369584 471436
rect 253992 471396 369584 471424
rect 253992 471384 253998 471396
rect 369578 471384 369584 471396
rect 369636 471384 369642 471436
rect 193214 471316 193220 471368
rect 193272 471356 193278 471368
rect 194134 471356 194140 471368
rect 193272 471328 194140 471356
rect 193272 471316 193278 471328
rect 194134 471316 194140 471328
rect 194192 471316 194198 471368
rect 198734 471316 198740 471368
rect 198792 471356 198798 471368
rect 199010 471356 199016 471368
rect 198792 471328 199016 471356
rect 198792 471316 198798 471328
rect 199010 471316 199016 471328
rect 199068 471316 199074 471368
rect 244458 471316 244464 471368
rect 244516 471356 244522 471368
rect 371970 471356 371976 471368
rect 244516 471328 371976 471356
rect 244516 471316 244522 471328
rect 371970 471316 371976 471328
rect 372028 471316 372034 471368
rect 57698 471248 57704 471300
rect 57756 471288 57762 471300
rect 113910 471288 113916 471300
rect 57756 471260 113916 471288
rect 57756 471248 57762 471260
rect 113910 471248 113916 471260
rect 113968 471248 113974 471300
rect 169386 471248 169392 471300
rect 169444 471288 169450 471300
rect 207658 471288 207664 471300
rect 169444 471260 207664 471288
rect 169444 471248 169450 471260
rect 207658 471248 207664 471260
rect 207716 471248 207722 471300
rect 226794 471248 226800 471300
rect 226852 471288 226858 471300
rect 376110 471288 376116 471300
rect 226852 471260 376116 471288
rect 226852 471248 226858 471260
rect 376110 471248 376116 471260
rect 376168 471248 376174 471300
rect 190454 471180 190460 471232
rect 190512 471220 190518 471232
rect 190638 471220 190644 471232
rect 190512 471192 190644 471220
rect 190512 471180 190518 471192
rect 190638 471180 190644 471192
rect 190696 471180 190702 471232
rect 191834 471180 191840 471232
rect 191892 471220 191898 471232
rect 192846 471220 192852 471232
rect 191892 471192 192852 471220
rect 191892 471180 191898 471192
rect 192846 471180 192852 471192
rect 192904 471180 192910 471232
rect 193306 471180 193312 471232
rect 193364 471220 193370 471232
rect 193766 471220 193772 471232
rect 193364 471192 193772 471220
rect 193364 471180 193370 471192
rect 193766 471180 193772 471192
rect 193824 471180 193830 471232
rect 198826 471180 198832 471232
rect 198884 471220 198890 471232
rect 199470 471220 199476 471232
rect 198884 471192 199476 471220
rect 198884 471180 198890 471192
rect 199470 471180 199476 471192
rect 199528 471180 199534 471232
rect 202874 471180 202880 471232
rect 202932 471220 202938 471232
rect 203150 471220 203156 471232
rect 202932 471192 203156 471220
rect 202932 471180 202938 471192
rect 203150 471180 203156 471192
rect 203208 471180 203214 471232
rect 204346 471180 204352 471232
rect 204404 471220 204410 471232
rect 205174 471220 205180 471232
rect 204404 471192 205180 471220
rect 204404 471180 204410 471192
rect 205174 471180 205180 471192
rect 205232 471180 205238 471232
rect 267734 471180 267740 471232
rect 267792 471220 267798 471232
rect 268102 471220 268108 471232
rect 267792 471192 268108 471220
rect 267792 471180 267798 471192
rect 268102 471180 268108 471192
rect 268160 471180 268166 471232
rect 203150 471044 203156 471096
rect 203208 471084 203214 471096
rect 203886 471084 203892 471096
rect 203208 471056 203892 471084
rect 203208 471044 203214 471056
rect 203886 471044 203892 471056
rect 203944 471044 203950 471096
rect 43622 470500 43628 470552
rect 43680 470540 43686 470552
rect 120166 470540 120172 470552
rect 43680 470512 120172 470540
rect 43680 470500 43686 470512
rect 120166 470500 120172 470512
rect 120224 470500 120230 470552
rect 43806 470432 43812 470484
rect 43864 470472 43870 470484
rect 121730 470472 121736 470484
rect 43864 470444 121736 470472
rect 43864 470432 43870 470444
rect 121730 470432 121736 470444
rect 121788 470432 121794 470484
rect 56042 470364 56048 470416
rect 56100 470404 56106 470416
rect 133966 470404 133972 470416
rect 56100 470376 133972 470404
rect 56100 470364 56106 470376
rect 133966 470364 133972 470376
rect 134024 470364 134030 470416
rect 42702 470296 42708 470348
rect 42760 470336 42766 470348
rect 121914 470336 121920 470348
rect 42760 470308 121920 470336
rect 42760 470296 42766 470308
rect 121914 470296 121920 470308
rect 121972 470296 121978 470348
rect 278866 470296 278872 470348
rect 278924 470336 278930 470348
rect 356974 470336 356980 470348
rect 278924 470308 356980 470336
rect 278924 470296 278930 470308
rect 356974 470296 356980 470308
rect 357032 470296 357038 470348
rect 45186 470228 45192 470280
rect 45244 470268 45250 470280
rect 124950 470268 124956 470280
rect 45244 470240 124956 470268
rect 45244 470228 45250 470240
rect 124950 470228 124956 470240
rect 125008 470228 125014 470280
rect 285950 470228 285956 470280
rect 286008 470268 286014 470280
rect 379146 470268 379152 470280
rect 286008 470240 379152 470268
rect 286008 470228 286014 470240
rect 379146 470228 379152 470240
rect 379204 470228 379210 470280
rect 43530 470160 43536 470212
rect 43588 470200 43594 470212
rect 122834 470200 122840 470212
rect 43588 470172 122840 470200
rect 43588 470160 43594 470172
rect 122834 470160 122840 470172
rect 122892 470160 122898 470212
rect 269942 470160 269948 470212
rect 270000 470200 270006 470212
rect 371786 470200 371792 470212
rect 270000 470172 371792 470200
rect 270000 470160 270006 470172
rect 371786 470160 371792 470172
rect 371844 470160 371850 470212
rect 43714 470092 43720 470144
rect 43772 470132 43778 470144
rect 124490 470132 124496 470144
rect 43772 470104 124496 470132
rect 43772 470092 43778 470104
rect 124490 470092 124496 470104
rect 124548 470092 124554 470144
rect 258166 470092 258172 470144
rect 258224 470132 258230 470144
rect 364058 470132 364064 470144
rect 258224 470104 364064 470132
rect 258224 470092 258230 470104
rect 364058 470092 364064 470104
rect 364116 470092 364122 470144
rect 42242 470024 42248 470076
rect 42300 470064 42306 470076
rect 123662 470064 123668 470076
rect 42300 470036 123668 470064
rect 42300 470024 42306 470036
rect 123662 470024 123668 470036
rect 123720 470024 123726 470076
rect 252646 470024 252652 470076
rect 252704 470064 252710 470076
rect 376478 470064 376484 470076
rect 252704 470036 376484 470064
rect 252704 470024 252710 470036
rect 376478 470024 376484 470036
rect 376536 470024 376542 470076
rect 42518 469956 42524 470008
rect 42576 469996 42582 470008
rect 124214 469996 124220 470008
rect 42576 469968 124220 469996
rect 42576 469956 42582 469968
rect 124214 469956 124220 469968
rect 124272 469956 124278 470008
rect 187142 469956 187148 470008
rect 187200 469996 187206 470008
rect 209222 469996 209228 470008
rect 187200 469968 209228 469996
rect 187200 469956 187206 469968
rect 209222 469956 209228 469968
rect 209280 469956 209286 470008
rect 245838 469956 245844 470008
rect 245896 469996 245902 470008
rect 370682 469996 370688 470008
rect 245896 469968 370688 469996
rect 245896 469956 245902 469968
rect 370682 469956 370688 469968
rect 370740 469956 370746 470008
rect 48958 469888 48964 469940
rect 49016 469928 49022 469940
rect 132678 469928 132684 469940
rect 49016 469900 132684 469928
rect 49016 469888 49022 469900
rect 132678 469888 132684 469900
rect 132736 469888 132742 469940
rect 176746 469888 176752 469940
rect 176804 469928 176810 469940
rect 204990 469928 204996 469940
rect 176804 469900 204996 469928
rect 176804 469888 176810 469900
rect 204990 469888 204996 469900
rect 205048 469888 205054 469940
rect 205910 469888 205916 469940
rect 205968 469928 205974 469940
rect 217594 469928 217600 469940
rect 205968 469900 217600 469928
rect 205968 469888 205974 469900
rect 217594 469888 217600 469900
rect 217652 469888 217658 469940
rect 242894 469888 242900 469940
rect 242952 469928 242958 469940
rect 374822 469928 374828 469940
rect 242952 469900 374828 469928
rect 242952 469888 242958 469900
rect 374822 469888 374828 469900
rect 374880 469888 374886 469940
rect 44726 469820 44732 469872
rect 44784 469860 44790 469872
rect 143626 469860 143632 469872
rect 44784 469832 143632 469860
rect 44784 469820 44790 469832
rect 143626 469820 143632 469832
rect 143684 469820 143690 469872
rect 165706 469820 165712 469872
rect 165764 469860 165770 469872
rect 211798 469860 211804 469872
rect 165764 469832 211804 469860
rect 165764 469820 165770 469832
rect 211798 469820 211804 469832
rect 211856 469820 211862 469872
rect 229186 469820 229192 469872
rect 229244 469860 229250 469872
rect 367922 469860 367928 469872
rect 229244 469832 367928 469860
rect 229244 469820 229250 469832
rect 367922 469820 367928 469832
rect 367980 469820 367986 469872
rect 53650 469752 53656 469804
rect 53708 469792 53714 469804
rect 127158 469792 127164 469804
rect 53708 469764 127164 469792
rect 53708 469752 53714 469764
rect 127158 469752 127164 469764
rect 127216 469752 127222 469804
rect 57054 469684 57060 469736
rect 57112 469724 57118 469736
rect 128446 469724 128452 469736
rect 57112 469696 128452 469724
rect 57112 469684 57118 469696
rect 128446 469684 128452 469696
rect 128504 469684 128510 469736
rect 58526 469616 58532 469668
rect 58584 469656 58590 469668
rect 128538 469656 128544 469668
rect 58584 469628 128544 469656
rect 58584 469616 58590 469628
rect 128538 469616 128544 469628
rect 128596 469616 128602 469668
rect 40954 469072 40960 469124
rect 41012 469112 41018 469124
rect 62114 469112 62120 469124
rect 41012 469084 62120 469112
rect 41012 469072 41018 469084
rect 62114 469072 62120 469084
rect 62172 469072 62178 469124
rect 289906 469072 289912 469124
rect 289964 469112 289970 469124
rect 362678 469112 362684 469124
rect 289964 469084 362684 469112
rect 289964 469072 289970 469084
rect 362678 469072 362684 469084
rect 362736 469072 362742 469124
rect 40862 469004 40868 469056
rect 40920 469044 40926 469056
rect 62206 469044 62212 469056
rect 40920 469016 62212 469044
rect 40920 469004 40926 469016
rect 62206 469004 62212 469016
rect 62264 469004 62270 469056
rect 274726 469004 274732 469056
rect 274784 469044 274790 469056
rect 363414 469044 363420 469056
rect 274784 469016 363420 469044
rect 274784 469004 274790 469016
rect 363414 469004 363420 469016
rect 363472 469004 363478 469056
rect 45094 468936 45100 468988
rect 45152 468976 45158 468988
rect 71038 468976 71044 468988
rect 45152 468948 71044 468976
rect 45152 468936 45158 468948
rect 71038 468936 71044 468948
rect 71096 468936 71102 468988
rect 178218 468936 178224 468988
rect 178276 468976 178282 468988
rect 202322 468976 202328 468988
rect 178276 468948 202328 468976
rect 178276 468936 178282 468948
rect 202322 468936 202328 468948
rect 202380 468936 202386 468988
rect 271230 468936 271236 468988
rect 271288 468976 271294 468988
rect 361298 468976 361304 468988
rect 271288 468948 361304 468976
rect 271288 468936 271294 468948
rect 361298 468936 361304 468948
rect 361356 468936 361362 468988
rect 44082 468868 44088 468920
rect 44140 468908 44146 468920
rect 70578 468908 70584 468920
rect 44140 468880 70584 468908
rect 44140 468868 44146 468880
rect 70578 468868 70584 468880
rect 70636 468868 70642 468920
rect 178678 468868 178684 468920
rect 178736 468908 178742 468920
rect 205910 468908 205916 468920
rect 178736 468880 205916 468908
rect 178736 468868 178742 468880
rect 205910 468868 205916 468880
rect 205968 468868 205974 468920
rect 273346 468868 273352 468920
rect 273404 468908 273410 468920
rect 368382 468908 368388 468920
rect 273404 468880 368388 468908
rect 273404 468868 273410 468880
rect 368382 468868 368388 468880
rect 368440 468868 368446 468920
rect 46566 468800 46572 468852
rect 46624 468840 46630 468852
rect 75270 468840 75276 468852
rect 46624 468812 75276 468840
rect 46624 468800 46630 468812
rect 75270 468800 75276 468812
rect 75328 468800 75334 468852
rect 161750 468800 161756 468852
rect 161808 468840 161814 468852
rect 210418 468840 210424 468852
rect 161808 468812 210424 468840
rect 161808 468800 161814 468812
rect 210418 468800 210424 468812
rect 210476 468800 210482 468852
rect 263778 468800 263784 468852
rect 263836 468840 263842 468852
rect 362586 468840 362592 468852
rect 263836 468812 362592 468840
rect 263836 468800 263842 468812
rect 362586 468800 362592 468812
rect 362644 468800 362650 468852
rect 41046 468732 41052 468784
rect 41104 468772 41110 468784
rect 93946 468772 93952 468784
rect 41104 468744 93952 468772
rect 41104 468732 41110 468744
rect 93946 468732 93952 468744
rect 94004 468732 94010 468784
rect 162946 468732 162952 468784
rect 163004 468772 163010 468784
rect 216030 468772 216036 468784
rect 163004 468744 216036 468772
rect 163004 468732 163010 468744
rect 216030 468732 216036 468744
rect 216088 468732 216094 468784
rect 262398 468732 262404 468784
rect 262456 468772 262462 468784
rect 368198 468772 368204 468784
rect 262456 468744 368204 468772
rect 262456 468732 262462 468744
rect 368198 468732 368204 468744
rect 368256 468732 368262 468784
rect 45002 468664 45008 468716
rect 45060 468704 45066 468716
rect 104986 468704 104992 468716
rect 45060 468676 104992 468704
rect 45060 468664 45066 468676
rect 104986 468664 104992 468676
rect 105044 468664 105050 468716
rect 139486 468664 139492 468716
rect 139544 468704 139550 468716
rect 207474 468704 207480 468716
rect 139544 468676 207480 468704
rect 139544 468664 139550 468676
rect 207474 468664 207480 468676
rect 207532 468664 207538 468716
rect 259546 468664 259552 468716
rect 259604 468704 259610 468716
rect 370866 468704 370872 468716
rect 259604 468676 370872 468704
rect 259604 468664 259610 468676
rect 370866 468664 370872 468676
rect 370924 468664 370930 468716
rect 44910 468596 44916 468648
rect 44968 468636 44974 468648
rect 106366 468636 106372 468648
rect 44968 468608 106372 468636
rect 44968 468596 44974 468608
rect 106366 468596 106372 468608
rect 106424 468596 106430 468648
rect 127710 468596 127716 468648
rect 127768 468636 127774 468648
rect 197630 468636 197636 468648
rect 127768 468608 197636 468636
rect 127768 468596 127774 468608
rect 197630 468596 197636 468608
rect 197688 468596 197694 468648
rect 245746 468596 245752 468648
rect 245804 468636 245810 468648
rect 365254 468636 365260 468648
rect 245804 468608 365260 468636
rect 245804 468596 245810 468608
rect 365254 468596 365260 468608
rect 365312 468596 365318 468648
rect 59354 468528 59360 468580
rect 59412 468568 59418 468580
rect 179598 468568 179604 468580
rect 59412 468540 179604 468568
rect 59412 468528 59418 468540
rect 179598 468528 179604 468540
rect 179656 468528 179662 468580
rect 187878 468528 187884 468580
rect 187936 468568 187942 468580
rect 209406 468568 209412 468580
rect 187936 468540 209412 468568
rect 187936 468528 187942 468540
rect 209406 468528 209412 468540
rect 209464 468528 209470 468580
rect 241606 468528 241612 468580
rect 241664 468568 241670 468580
rect 366542 468568 366548 468580
rect 241664 468540 366548 468568
rect 241664 468528 241670 468540
rect 366542 468528 366548 468540
rect 366600 468528 366606 468580
rect 15838 468460 15844 468512
rect 15896 468500 15902 468512
rect 378134 468500 378140 468512
rect 15896 468472 378140 468500
rect 15896 468460 15902 468472
rect 378134 468460 378140 468472
rect 378192 468460 378198 468512
rect 285858 467712 285864 467764
rect 285916 467752 285922 467764
rect 357066 467752 357072 467764
rect 285916 467724 357072 467752
rect 285916 467712 285922 467724
rect 357066 467712 357072 467724
rect 357124 467712 357130 467764
rect 294138 467644 294144 467696
rect 294196 467684 294202 467696
rect 376570 467684 376576 467696
rect 294196 467656 376576 467684
rect 294196 467644 294202 467656
rect 376570 467644 376576 467656
rect 376628 467644 376634 467696
rect 265066 467576 265072 467628
rect 265124 467616 265130 467628
rect 365530 467616 365536 467628
rect 265124 467588 365536 467616
rect 265124 467576 265130 467588
rect 365530 467576 365536 467588
rect 365588 467576 365594 467628
rect 269206 467508 269212 467560
rect 269264 467548 269270 467560
rect 375926 467548 375932 467560
rect 269264 467520 375932 467548
rect 269264 467508 269270 467520
rect 375926 467508 375932 467520
rect 375984 467508 375990 467560
rect 268654 467440 268660 467492
rect 268712 467480 268718 467492
rect 375282 467480 375288 467492
rect 268712 467452 375288 467480
rect 268712 467440 268718 467452
rect 375282 467440 375288 467452
rect 375340 467440 375346 467492
rect 253934 467372 253940 467424
rect 253992 467412 253998 467424
rect 364150 467412 364156 467424
rect 253992 467384 364156 467412
rect 253992 467372 253998 467384
rect 364150 467372 364156 467384
rect 364208 467372 364214 467424
rect 187970 467304 187976 467356
rect 188028 467344 188034 467356
rect 200758 467344 200764 467356
rect 188028 467316 200764 467344
rect 188028 467304 188034 467316
rect 200758 467304 200764 467316
rect 200816 467304 200822 467356
rect 207290 467304 207296 467356
rect 207348 467344 207354 467356
rect 217686 467344 217692 467356
rect 207348 467316 217692 467344
rect 207348 467304 207354 467316
rect 217686 467304 217692 467316
rect 217744 467304 217750 467356
rect 258074 467304 258080 467356
rect 258132 467344 258138 467356
rect 373442 467344 373448 467356
rect 258132 467316 373448 467344
rect 258132 467304 258138 467316
rect 373442 467304 373448 467316
rect 373500 467304 373506 467356
rect 185118 467236 185124 467288
rect 185176 467276 185182 467288
rect 214650 467276 214656 467288
rect 185176 467248 214656 467276
rect 185176 467236 185182 467248
rect 214650 467236 214656 467248
rect 214708 467236 214714 467288
rect 244458 467236 244464 467288
rect 244516 467276 244522 467288
rect 360930 467276 360936 467288
rect 244516 467248 360936 467276
rect 244516 467236 244522 467248
rect 360930 467236 360936 467248
rect 360988 467236 360994 467288
rect 176654 467168 176660 467220
rect 176712 467208 176718 467220
rect 207842 467208 207848 467220
rect 176712 467180 207848 467208
rect 176712 467168 176718 467180
rect 207842 467168 207848 467180
rect 207900 467168 207906 467220
rect 237374 467168 237380 467220
rect 237432 467208 237438 467220
rect 358262 467208 358268 467220
rect 237432 467180 358268 467208
rect 237432 467168 237438 467180
rect 358262 467168 358268 467180
rect 358320 467168 358326 467220
rect 57514 467100 57520 467152
rect 57572 467140 57578 467152
rect 114738 467140 114744 467152
rect 57572 467112 114744 467140
rect 57572 467100 57578 467112
rect 114738 467100 114744 467112
rect 114796 467100 114802 467152
rect 171410 467100 171416 467152
rect 171468 467140 171474 467152
rect 209038 467140 209044 467152
rect 171468 467112 209044 467140
rect 171468 467100 171474 467112
rect 209038 467100 209044 467112
rect 209096 467100 209102 467152
rect 227714 467100 227720 467152
rect 227772 467140 227778 467152
rect 370498 467140 370504 467152
rect 227772 467112 370504 467140
rect 227772 467100 227778 467112
rect 370498 467100 370504 467112
rect 370556 467100 370562 467152
rect 44818 466352 44824 466404
rect 44876 466392 44882 466404
rect 68370 466392 68376 466404
rect 44876 466364 68376 466392
rect 44876 466352 44882 466364
rect 68370 466352 68376 466364
rect 68428 466352 68434 466404
rect 182450 466352 182456 466404
rect 182508 466392 182514 466404
rect 206554 466392 206560 466404
rect 182508 466364 206560 466392
rect 182508 466352 182514 466364
rect 206554 466352 206560 466364
rect 206612 466352 206618 466404
rect 52086 466284 52092 466336
rect 52144 466324 52150 466336
rect 82814 466324 82820 466336
rect 52144 466296 82820 466324
rect 52144 466284 52150 466296
rect 82814 466284 82820 466296
rect 82872 466284 82878 466336
rect 190638 466284 190644 466336
rect 190696 466324 190702 466336
rect 214834 466324 214840 466336
rect 190696 466296 214840 466324
rect 190696 466284 190702 466296
rect 214834 466284 214840 466296
rect 214892 466284 214898 466336
rect 50522 466216 50528 466268
rect 50580 466256 50586 466268
rect 82906 466256 82912 466268
rect 50580 466228 82912 466256
rect 50580 466216 50586 466228
rect 82906 466216 82912 466228
rect 82964 466216 82970 466268
rect 191926 466216 191932 466268
rect 191984 466256 191990 466268
rect 216306 466256 216312 466268
rect 191984 466228 216312 466256
rect 191984 466216 191990 466228
rect 216306 466216 216312 466228
rect 216364 466216 216370 466268
rect 289814 466216 289820 466268
rect 289872 466256 289878 466268
rect 361390 466256 361396 466268
rect 289872 466228 361396 466256
rect 289872 466216 289878 466228
rect 361390 466216 361396 466228
rect 361448 466216 361454 466268
rect 42426 466148 42432 466200
rect 42484 466188 42490 466200
rect 75178 466188 75184 466200
rect 42484 466160 75184 466188
rect 42484 466148 42490 466160
rect 75178 466148 75184 466160
rect 75236 466148 75242 466200
rect 182358 466148 182364 466200
rect 182416 466188 182422 466200
rect 207934 466188 207940 466200
rect 182416 466160 207940 466188
rect 182416 466148 182422 466160
rect 207934 466148 207940 466160
rect 207992 466148 207998 466200
rect 299474 466148 299480 466200
rect 299532 466188 299538 466200
rect 371234 466188 371240 466200
rect 299532 466160 371240 466188
rect 299532 466148 299538 466160
rect 371234 466148 371240 466160
rect 371292 466148 371298 466200
rect 48222 466080 48228 466132
rect 48280 466120 48286 466132
rect 81526 466120 81532 466132
rect 48280 466092 81532 466120
rect 48280 466080 48286 466092
rect 81526 466080 81532 466092
rect 81584 466080 81590 466132
rect 174078 466080 174084 466132
rect 174136 466120 174142 466132
rect 200850 466120 200856 466132
rect 174136 466092 200856 466120
rect 174136 466080 174142 466092
rect 200850 466080 200856 466092
rect 200908 466080 200914 466132
rect 296806 466080 296812 466132
rect 296864 466120 296870 466132
rect 369026 466120 369032 466132
rect 296864 466092 369032 466120
rect 296864 466080 296870 466092
rect 369026 466080 369032 466092
rect 369084 466080 369090 466132
rect 49418 466012 49424 466064
rect 49476 466052 49482 466064
rect 82998 466052 83004 466064
rect 49476 466024 83004 466052
rect 49476 466012 49482 466024
rect 82998 466012 83004 466024
rect 83056 466012 83062 466064
rect 192018 466012 192024 466064
rect 192076 466052 192082 466064
rect 219158 466052 219164 466064
rect 192076 466024 219164 466052
rect 192076 466012 192082 466024
rect 219158 466012 219164 466024
rect 219216 466012 219222 466064
rect 298186 466012 298192 466064
rect 298244 466052 298250 466064
rect 373166 466052 373172 466064
rect 298244 466024 373172 466052
rect 298244 466012 298250 466024
rect 373166 466012 373172 466024
rect 373224 466012 373230 466064
rect 59814 465944 59820 465996
rect 59872 465984 59878 465996
rect 102226 465984 102232 465996
rect 59872 465956 102232 465984
rect 59872 465944 59878 465956
rect 102226 465944 102232 465956
rect 102284 465944 102290 465996
rect 139394 465944 139400 465996
rect 139452 465984 139458 465996
rect 197078 465984 197084 465996
rect 139452 465956 197084 465984
rect 139452 465944 139458 465956
rect 197078 465944 197084 465956
rect 197136 465944 197142 465996
rect 288526 465944 288532 465996
rect 288584 465984 288590 465996
rect 371050 465984 371056 465996
rect 288584 465956 371056 465984
rect 288584 465944 288590 465956
rect 371050 465944 371056 465956
rect 371108 465944 371114 465996
rect 57238 465876 57244 465928
rect 57296 465916 57302 465928
rect 103606 465916 103612 465928
rect 57296 465888 103612 465916
rect 57296 465876 57302 465888
rect 103606 465876 103612 465888
rect 103664 465876 103670 465928
rect 140958 465876 140964 465928
rect 141016 465916 141022 465928
rect 200574 465916 200580 465928
rect 141016 465888 200580 465916
rect 141016 465876 141022 465888
rect 200574 465876 200580 465888
rect 200632 465876 200638 465928
rect 240226 465876 240232 465928
rect 240284 465916 240290 465928
rect 366634 465916 366640 465928
rect 240284 465888 366640 465916
rect 240284 465876 240290 465888
rect 366634 465876 366640 465888
rect 366692 465876 366698 465928
rect 53190 465808 53196 465860
rect 53248 465848 53254 465860
rect 100846 465848 100852 465860
rect 53248 465820 100852 465848
rect 53248 465808 53254 465820
rect 100846 465808 100852 465820
rect 100904 465808 100910 465860
rect 140774 465808 140780 465860
rect 140832 465848 140838 465860
rect 201770 465848 201776 465860
rect 140832 465820 201776 465848
rect 140832 465808 140838 465820
rect 201770 465808 201776 465820
rect 201828 465808 201834 465860
rect 241514 465808 241520 465860
rect 241572 465848 241578 465860
rect 369302 465848 369308 465860
rect 241572 465820 369308 465848
rect 241572 465808 241578 465820
rect 369302 465808 369308 465820
rect 369360 465808 369366 465860
rect 58710 465740 58716 465792
rect 58768 465780 58774 465792
rect 110598 465780 110604 465792
rect 58768 465752 110604 465780
rect 58768 465740 58774 465752
rect 110598 465740 110604 465752
rect 110656 465740 110662 465792
rect 140866 465740 140872 465792
rect 140924 465780 140930 465792
rect 204530 465780 204536 465792
rect 140924 465752 204536 465780
rect 140924 465740 140930 465752
rect 204530 465740 204536 465752
rect 204588 465740 204594 465792
rect 226334 465740 226340 465792
rect 226392 465780 226398 465792
rect 363690 465780 363696 465792
rect 226392 465752 363696 465780
rect 226392 465740 226398 465752
rect 363690 465740 363696 465752
rect 363748 465740 363754 465792
rect 53098 465672 53104 465724
rect 53156 465712 53162 465724
rect 100938 465712 100944 465724
rect 53156 465684 100944 465712
rect 53156 465672 53162 465684
rect 100938 465672 100944 465684
rect 100996 465672 101002 465724
rect 107838 465672 107844 465724
rect 107896 465712 107902 465724
rect 202966 465712 202972 465724
rect 107896 465684 202972 465712
rect 107896 465672 107902 465684
rect 202966 465672 202972 465684
rect 203024 465672 203030 465724
rect 226426 465672 226432 465724
rect 226484 465712 226490 465724
rect 371878 465712 371884 465724
rect 226484 465684 371884 465712
rect 226484 465672 226490 465684
rect 371878 465672 371884 465684
rect 371936 465672 371942 465724
rect 40770 465604 40776 465656
rect 40828 465644 40834 465656
rect 60826 465644 60832 465656
rect 40828 465616 60832 465644
rect 40828 465604 40834 465616
rect 60826 465604 60832 465616
rect 60884 465604 60890 465656
rect 183646 465604 183652 465656
rect 183704 465644 183710 465656
rect 205174 465644 205180 465656
rect 183704 465616 205180 465644
rect 183704 465604 183710 465616
rect 205174 465604 205180 465616
rect 205232 465604 205238 465656
rect 46290 465536 46296 465588
rect 46348 465576 46354 465588
rect 64966 465576 64972 465588
rect 46348 465548 64972 465576
rect 46348 465536 46354 465548
rect 64966 465536 64972 465548
rect 65024 465536 65030 465588
rect 182266 465536 182272 465588
rect 182324 465576 182330 465588
rect 202414 465576 202420 465588
rect 182324 465548 202420 465576
rect 182324 465536 182330 465548
rect 202414 465536 202420 465548
rect 202472 465536 202478 465588
rect 47486 465468 47492 465520
rect 47544 465508 47550 465520
rect 65058 465508 65064 465520
rect 47544 465480 65064 465508
rect 47544 465468 47550 465480
rect 65058 465468 65064 465480
rect 65116 465468 65122 465520
rect 192110 465468 192116 465520
rect 192168 465508 192174 465520
rect 208026 465508 208032 465520
rect 192168 465480 208032 465508
rect 192168 465468 192174 465480
rect 208026 465468 208032 465480
rect 208084 465468 208090 465520
rect 294046 464856 294052 464908
rect 294104 464896 294110 464908
rect 358538 464896 358544 464908
rect 294104 464868 358544 464896
rect 294104 464856 294110 464868
rect 358538 464856 358544 464868
rect 358596 464856 358602 464908
rect 292666 464788 292672 464840
rect 292724 464828 292730 464840
rect 367646 464828 367652 464840
rect 292724 464800 367652 464828
rect 292724 464788 292730 464800
rect 367646 464788 367652 464800
rect 367704 464788 367710 464840
rect 283006 464720 283012 464772
rect 283064 464760 283070 464772
rect 357986 464760 357992 464772
rect 283064 464732 357992 464760
rect 283064 464720 283070 464732
rect 357986 464720 357992 464732
rect 358044 464720 358050 464772
rect 284386 464652 284392 464704
rect 284444 464692 284450 464704
rect 359918 464692 359924 464704
rect 284444 464664 359924 464692
rect 284444 464652 284450 464664
rect 359918 464652 359924 464664
rect 359976 464652 359982 464704
rect 284478 464584 284484 464636
rect 284536 464624 284542 464636
rect 360562 464624 360568 464636
rect 284536 464596 360568 464624
rect 284536 464584 284542 464596
rect 360562 464584 360568 464596
rect 360620 464584 360626 464636
rect 293954 464516 293960 464568
rect 294012 464556 294018 464568
rect 377858 464556 377864 464568
rect 294012 464528 377864 464556
rect 294012 464516 294018 464528
rect 377858 464516 377864 464528
rect 377916 464516 377922 464568
rect 291286 464448 291292 464500
rect 291344 464488 291350 464500
rect 378042 464488 378048 464500
rect 291344 464460 378048 464488
rect 291344 464448 291350 464460
rect 378042 464448 378048 464460
rect 378100 464448 378106 464500
rect 285766 464380 285772 464432
rect 285824 464420 285830 464432
rect 377490 464420 377496 464432
rect 285824 464392 377496 464420
rect 285824 464380 285830 464392
rect 377490 464380 377496 464392
rect 377548 464380 377554 464432
rect 57606 464312 57612 464364
rect 57664 464352 57670 464364
rect 111978 464352 111984 464364
rect 57664 464324 111984 464352
rect 57664 464312 57670 464324
rect 111978 464312 111984 464324
rect 112036 464312 112042 464364
rect 158714 464312 158720 464364
rect 158772 464352 158778 464364
rect 203518 464352 203524 464364
rect 158772 464324 203524 464352
rect 158772 464312 158778 464324
rect 203518 464312 203524 464324
rect 203576 464312 203582 464364
rect 284294 464312 284300 464364
rect 284352 464352 284358 464364
rect 377398 464352 377404 464364
rect 284352 464324 377404 464352
rect 284352 464312 284358 464324
rect 377398 464312 377404 464324
rect 377456 464312 377462 464364
rect 55858 463632 55864 463684
rect 55916 463672 55922 463684
rect 87138 463672 87144 463684
rect 55916 463644 87144 463672
rect 55916 463632 55922 463644
rect 87138 463632 87144 463644
rect 87196 463632 87202 463684
rect 185026 463632 185032 463684
rect 185084 463672 185090 463684
rect 212074 463672 212080 463684
rect 185084 463644 212080 463672
rect 185084 463632 185090 463644
rect 212074 463632 212080 463644
rect 212132 463632 212138 463684
rect 282914 463632 282920 463684
rect 282972 463672 282978 463684
rect 359826 463672 359832 463684
rect 282972 463644 359832 463672
rect 282972 463632 282978 463644
rect 359826 463632 359832 463644
rect 359884 463632 359890 463684
rect 55030 463564 55036 463616
rect 55088 463604 55094 463616
rect 86954 463604 86960 463616
rect 55088 463576 86960 463604
rect 55088 463564 55094 463576
rect 86954 463564 86960 463576
rect 87012 463564 87018 463616
rect 190454 463564 190460 463616
rect 190512 463604 190518 463616
rect 217502 463604 217508 463616
rect 190512 463576 217508 463604
rect 190512 463564 190518 463576
rect 217502 463564 217508 463576
rect 217560 463564 217566 463616
rect 277578 463564 277584 463616
rect 277636 463604 277642 463616
rect 360654 463604 360660 463616
rect 277636 463576 360660 463604
rect 277636 463564 277642 463576
rect 360654 463564 360660 463576
rect 360712 463564 360718 463616
rect 48866 463496 48872 463548
rect 48924 463536 48930 463548
rect 81618 463536 81624 463548
rect 48924 463508 81624 463536
rect 48924 463496 48930 463508
rect 81618 463496 81624 463508
rect 81676 463496 81682 463548
rect 186314 463496 186320 463548
rect 186372 463536 186378 463548
rect 213454 463536 213460 463548
rect 186372 463508 213460 463536
rect 186372 463496 186378 463508
rect 213454 463496 213460 463508
rect 213512 463496 213518 463548
rect 276198 463496 276204 463548
rect 276256 463536 276262 463548
rect 364794 463536 364800 463548
rect 276256 463508 364800 463536
rect 276256 463496 276262 463508
rect 364794 463496 364800 463508
rect 364852 463496 364858 463548
rect 56226 463428 56232 463480
rect 56284 463468 56290 463480
rect 88426 463468 88432 463480
rect 56284 463440 88432 463468
rect 56284 463428 56290 463440
rect 88426 463428 88432 463440
rect 88484 463428 88490 463480
rect 180978 463428 180984 463480
rect 181036 463468 181042 463480
rect 210694 463468 210700 463480
rect 181036 463440 210700 463468
rect 181036 463428 181042 463440
rect 210694 463428 210700 463440
rect 210752 463428 210758 463480
rect 277394 463428 277400 463480
rect 277452 463468 277458 463480
rect 367554 463468 367560 463480
rect 277452 463440 367560 463468
rect 277452 463428 277458 463440
rect 367554 463428 367560 463440
rect 367612 463428 367618 463480
rect 56134 463360 56140 463412
rect 56192 463400 56198 463412
rect 88610 463400 88616 463412
rect 56192 463372 88616 463400
rect 56192 463360 56198 463372
rect 88610 463360 88616 463372
rect 88668 463360 88674 463412
rect 180886 463360 180892 463412
rect 180944 463400 180950 463412
rect 212166 463400 212172 463412
rect 180944 463372 212172 463400
rect 180944 463360 180950 463372
rect 212166 463360 212172 463372
rect 212224 463360 212230 463412
rect 273254 463360 273260 463412
rect 273312 463400 273318 463412
rect 366174 463400 366180 463412
rect 273312 463372 366180 463400
rect 273312 463360 273318 463372
rect 366174 463360 366180 463372
rect 366232 463360 366238 463412
rect 52914 463292 52920 463344
rect 52972 463332 52978 463344
rect 85666 463332 85672 463344
rect 52972 463304 85672 463332
rect 52972 463292 52978 463304
rect 85666 463292 85672 463304
rect 85724 463292 85730 463344
rect 175274 463292 175280 463344
rect 175332 463332 175338 463344
rect 206646 463332 206652 463344
rect 175332 463304 206652 463332
rect 175332 463292 175338 463304
rect 206646 463292 206652 463304
rect 206704 463292 206710 463344
rect 267826 463292 267832 463344
rect 267884 463332 267890 463344
rect 362862 463332 362868 463344
rect 267884 463304 362868 463332
rect 267884 463292 267890 463304
rect 362862 463292 362868 463304
rect 362920 463292 362926 463344
rect 56410 463224 56416 463276
rect 56468 463264 56474 463276
rect 89714 463264 89720 463276
rect 56468 463236 89720 463264
rect 56468 463224 56474 463236
rect 89714 463224 89720 463236
rect 89772 463224 89778 463276
rect 168374 463224 168380 463276
rect 168432 463264 168438 463276
rect 209130 463264 209136 463276
rect 168432 463236 209136 463264
rect 168432 463224 168438 463236
rect 209130 463224 209136 463236
rect 209188 463224 209194 463276
rect 274634 463224 274640 463276
rect 274692 463264 274698 463276
rect 370406 463264 370412 463276
rect 274692 463236 370412 463264
rect 274692 463224 274698 463236
rect 370406 463224 370412 463236
rect 370464 463224 370470 463276
rect 54846 463156 54852 463208
rect 54904 463196 54910 463208
rect 88518 463196 88524 463208
rect 54904 463168 88524 463196
rect 54904 463156 54910 463168
rect 88518 463156 88524 463168
rect 88576 463156 88582 463208
rect 160094 463156 160100 463208
rect 160152 463196 160158 463208
rect 202138 463196 202144 463208
rect 160152 463168 202144 463196
rect 160152 463156 160158 463168
rect 202138 463156 202144 463168
rect 202196 463156 202202 463208
rect 267734 463156 267740 463208
rect 267792 463196 267798 463208
rect 367002 463196 367008 463208
rect 267792 463168 367008 463196
rect 267792 463156 267798 463168
rect 367002 463156 367008 463168
rect 367060 463156 367066 463208
rect 57422 463088 57428 463140
rect 57480 463128 57486 463140
rect 113358 463128 113364 463140
rect 57480 463100 113364 463128
rect 57480 463088 57486 463100
rect 113358 463088 113364 463100
rect 113416 463088 113422 463140
rect 142338 463088 142344 463140
rect 142396 463128 142402 463140
rect 208486 463128 208492 463140
rect 142396 463100 208492 463128
rect 142396 463088 142402 463100
rect 208486 463088 208492 463100
rect 208544 463088 208550 463140
rect 249978 463088 249984 463140
rect 250036 463128 250042 463140
rect 370774 463128 370780 463140
rect 250036 463100 370780 463128
rect 250036 463088 250042 463100
rect 370774 463088 370780 463100
rect 370832 463088 370838 463140
rect 53282 463020 53288 463072
rect 53340 463060 53346 463072
rect 87046 463060 87052 463072
rect 53340 463032 87052 463060
rect 53340 463020 53346 463032
rect 87046 463020 87052 463032
rect 87104 463020 87110 463072
rect 109034 463020 109040 463072
rect 109092 463060 109098 463072
rect 200390 463060 200396 463072
rect 109092 463032 200396 463060
rect 109092 463020 109098 463032
rect 200390 463020 200396 463032
rect 200448 463020 200454 463072
rect 248598 463020 248604 463072
rect 248656 463060 248662 463072
rect 372062 463060 372068 463072
rect 248656 463032 372068 463060
rect 248656 463020 248662 463032
rect 372062 463020 372068 463032
rect 372120 463020 372126 463072
rect 53374 462952 53380 463004
rect 53432 462992 53438 463004
rect 92566 462992 92572 463004
rect 53432 462964 92572 462992
rect 53432 462952 53438 462964
rect 92566 462952 92572 462964
rect 92624 462952 92630 463004
rect 107654 462952 107660 463004
rect 107712 462992 107718 463004
rect 200298 462992 200304 463004
rect 107712 462964 200304 462992
rect 107712 462952 107718 462964
rect 200298 462952 200304 462964
rect 200356 462952 200362 463004
rect 240134 462952 240140 463004
rect 240192 462992 240198 463004
rect 363782 462992 363788 463004
rect 240192 462964 363788 462992
rect 240192 462952 240198 462964
rect 363782 462952 363788 462964
rect 363840 462952 363846 463004
rect 54938 462884 54944 462936
rect 54996 462924 55002 462936
rect 85574 462924 85580 462936
rect 54996 462896 85580 462924
rect 54996 462884 55002 462896
rect 85574 462884 85580 462896
rect 85632 462884 85638 462936
rect 190546 462884 190552 462936
rect 190604 462924 190610 462936
rect 203794 462924 203800 462936
rect 190604 462896 203800 462924
rect 190604 462884 190610 462896
rect 203794 462884 203800 462896
rect 203852 462884 203858 462936
rect 40586 462816 40592 462868
rect 40644 462856 40650 462868
rect 60734 462856 60740 462868
rect 40644 462828 60740 462856
rect 40644 462816 40650 462828
rect 60734 462816 60740 462828
rect 60792 462816 60798 462868
rect 189258 462816 189264 462868
rect 189316 462856 189322 462868
rect 199378 462856 199384 462868
rect 189316 462828 199384 462856
rect 189316 462816 189322 462828
rect 199378 462816 199384 462828
rect 199436 462816 199442 462868
rect 46198 462748 46204 462800
rect 46256 462788 46262 462800
rect 64874 462788 64880 462800
rect 46256 462760 64880 462788
rect 46256 462748 46262 462760
rect 64874 462748 64880 462760
rect 64932 462748 64938 462800
rect 193398 462544 193404 462596
rect 193456 462584 193462 462596
rect 202506 462584 202512 462596
rect 193456 462556 202512 462584
rect 193456 462544 193462 462556
rect 202506 462544 202512 462556
rect 202564 462544 202570 462596
rect 133138 462272 133144 462324
rect 133196 462312 133202 462324
rect 178310 462312 178316 462324
rect 133196 462284 178316 462312
rect 133196 462272 133202 462284
rect 178310 462272 178316 462284
rect 178368 462272 178374 462324
rect 287146 462204 287152 462256
rect 287204 462244 287210 462256
rect 362770 462244 362776 462256
rect 287204 462216 362776 462244
rect 287204 462204 287210 462216
rect 362770 462204 362776 462216
rect 362828 462204 362834 462256
rect 298094 462136 298100 462188
rect 298152 462176 298158 462188
rect 375742 462176 375748 462188
rect 298152 462148 375748 462176
rect 298152 462136 298158 462148
rect 375742 462136 375748 462148
rect 375800 462136 375806 462188
rect 280154 462068 280160 462120
rect 280212 462108 280218 462120
rect 363322 462108 363328 462120
rect 280212 462080 363328 462108
rect 280212 462068 280218 462080
rect 363322 462068 363328 462080
rect 363380 462068 363386 462120
rect 260834 462000 260840 462052
rect 260892 462040 260898 462052
rect 361114 462040 361120 462052
rect 260892 462012 361120 462040
rect 260892 462000 260898 462012
rect 361114 462000 361120 462012
rect 361172 462000 361178 462052
rect 269114 461932 269120 461984
rect 269172 461972 269178 461984
rect 370314 461972 370320 461984
rect 269172 461944 370320 461972
rect 269172 461932 269178 461944
rect 370314 461932 370320 461944
rect 370372 461932 370378 461984
rect 191834 461864 191840 461916
rect 191892 461904 191898 461916
rect 205358 461904 205364 461916
rect 191892 461876 205364 461904
rect 191892 461864 191898 461876
rect 205358 461864 205364 461876
rect 205416 461864 205422 461916
rect 263594 461864 263600 461916
rect 263652 461904 263658 461916
rect 372338 461904 372344 461916
rect 263652 461876 372344 461904
rect 263652 461864 263658 461876
rect 372338 461864 372344 461876
rect 372396 461864 372402 461916
rect 511258 461864 511264 461916
rect 511316 461904 511322 461916
rect 517514 461904 517520 461916
rect 511316 461876 517520 461904
rect 511316 461864 511322 461876
rect 517514 461864 517520 461876
rect 517572 461864 517578 461916
rect 182174 461796 182180 461848
rect 182232 461836 182238 461848
rect 203610 461836 203616 461848
rect 182232 461808 203616 461836
rect 182232 461796 182238 461808
rect 203610 461796 203616 461808
rect 203668 461796 203674 461848
rect 264974 461796 264980 461848
rect 265032 461836 265038 461848
rect 375098 461836 375104 461848
rect 265032 461808 375104 461836
rect 265032 461796 265038 461808
rect 375098 461796 375104 461808
rect 375156 461796 375162 461848
rect 179598 461728 179604 461780
rect 179656 461768 179662 461780
rect 201586 461768 201592 461780
rect 179656 461740 201592 461768
rect 179656 461728 179662 461740
rect 201586 461728 201592 461740
rect 201644 461728 201650 461780
rect 262306 461728 262312 461780
rect 262364 461768 262370 461780
rect 373534 461768 373540 461780
rect 262364 461740 373540 461768
rect 262364 461728 262370 461740
rect 373534 461728 373540 461740
rect 373592 461728 373598 461780
rect 179506 461660 179512 461712
rect 179564 461700 179570 461712
rect 206738 461700 206744 461712
rect 179564 461672 206744 461700
rect 179564 461660 179570 461672
rect 206738 461660 206744 461672
rect 206796 461660 206802 461712
rect 251266 461660 251272 461712
rect 251324 461700 251330 461712
rect 365346 461700 365352 461712
rect 251324 461672 365352 461700
rect 251324 461660 251330 461672
rect 365346 461660 365352 461672
rect 365404 461660 365410 461712
rect 161566 461592 161572 461644
rect 161624 461632 161630 461644
rect 213270 461632 213276 461644
rect 161624 461604 213276 461632
rect 161624 461592 161630 461604
rect 213270 461592 213276 461604
rect 213328 461592 213334 461644
rect 252554 461592 252560 461644
rect 252612 461632 252618 461644
rect 375006 461632 375012 461644
rect 252612 461604 375012 461632
rect 252612 461592 252618 461604
rect 375006 461592 375012 461604
rect 375064 461592 375070 461644
rect 178310 461048 178316 461100
rect 178368 461088 178374 461100
rect 210050 461088 210056 461100
rect 178368 461060 210056 461088
rect 178368 461048 178374 461060
rect 210050 461048 210056 461060
rect 210108 461048 210114 461100
rect 338298 461048 338304 461100
rect 338356 461088 338362 461100
rect 357434 461088 357440 461100
rect 338356 461060 357440 461088
rect 338356 461048 338362 461060
rect 357434 461048 357440 461060
rect 357492 461088 357498 461100
rect 498378 461088 498384 461100
rect 357492 461060 498384 461088
rect 357492 461048 357498 461060
rect 498378 461048 498384 461060
rect 498436 461048 498442 461100
rect 201586 460980 201592 461032
rect 201644 461020 201650 461032
rect 339770 461020 339776 461032
rect 201644 460992 339776 461020
rect 201644 460980 201650 460992
rect 339770 460980 339776 460992
rect 339828 461020 339834 461032
rect 358814 461020 358820 461032
rect 339828 460992 358820 461020
rect 339828 460980 339834 460992
rect 358814 460980 358820 460992
rect 358872 461020 358878 461032
rect 499850 461020 499856 461032
rect 358872 460992 499856 461020
rect 358872 460980 358878 460992
rect 499850 460980 499856 460992
rect 499908 461020 499914 461032
rect 517606 461020 517612 461032
rect 499908 460992 517612 461020
rect 499908 460980 499914 460992
rect 517606 460980 517612 460992
rect 517664 460980 517670 461032
rect 190914 460912 190920 460964
rect 190972 460952 190978 460964
rect 207014 460952 207020 460964
rect 190972 460924 207020 460952
rect 190972 460912 190978 460924
rect 207014 460912 207020 460924
rect 207072 460912 207078 460964
rect 210050 460912 210056 460964
rect 210108 460952 210114 460964
rect 338298 460952 338304 460964
rect 210108 460924 338304 460952
rect 210108 460912 210114 460924
rect 338298 460912 338304 460924
rect 338356 460912 338362 460964
rect 350994 460912 351000 460964
rect 351052 460952 351058 460964
rect 367738 460952 367744 460964
rect 351052 460924 367744 460952
rect 351052 460912 351058 460924
rect 367738 460912 367744 460924
rect 367796 460912 367802 460964
rect 498378 460912 498384 460964
rect 498436 460952 498442 460964
rect 517698 460952 517704 460964
rect 498436 460924 517704 460952
rect 498436 460912 498442 460924
rect 517698 460912 517704 460924
rect 517756 460912 517762 460964
rect 48682 460844 48688 460896
rect 48740 460884 48746 460896
rect 78766 460884 78772 460896
rect 48740 460856 78772 460884
rect 48740 460844 48746 460856
rect 78766 460844 78772 460856
rect 78824 460844 78830 460896
rect 157334 460844 157340 460896
rect 157392 460884 157398 460896
rect 218330 460884 218336 460896
rect 157392 460856 218336 460884
rect 157392 460844 157398 460856
rect 218330 460844 218336 460856
rect 218388 460844 218394 460896
rect 285674 460844 285680 460896
rect 285732 460884 285738 460896
rect 377122 460884 377128 460896
rect 285732 460856 377128 460884
rect 285732 460844 285738 460856
rect 377122 460844 377128 460856
rect 377180 460844 377186 460896
rect 53374 460776 53380 460828
rect 53432 460816 53438 460828
rect 78674 460816 78680 460828
rect 53432 460788 78680 460816
rect 53432 460776 53438 460788
rect 78674 460776 78680 460788
rect 78732 460776 78738 460828
rect 193858 460776 193864 460828
rect 193916 460816 193922 460828
rect 203334 460816 203340 460828
rect 193916 460788 203340 460816
rect 193916 460776 193922 460788
rect 203334 460776 203340 460788
rect 203392 460776 203398 460828
rect 287054 460776 287060 460828
rect 287112 460816 287118 460828
rect 379422 460816 379428 460828
rect 287112 460788 379428 460816
rect 287112 460776 287118 460788
rect 379422 460776 379428 460788
rect 379480 460776 379486 460828
rect 51626 460708 51632 460760
rect 51684 460748 51690 460760
rect 76098 460748 76104 460760
rect 51684 460720 76104 460748
rect 51684 460708 51690 460720
rect 76098 460708 76104 460720
rect 76156 460708 76162 460760
rect 189166 460708 189172 460760
rect 189224 460748 189230 460760
rect 202598 460748 202604 460760
rect 189224 460720 202604 460748
rect 189224 460708 189230 460720
rect 202598 460708 202604 460720
rect 202656 460708 202662 460760
rect 266354 460708 266360 460760
rect 266412 460748 266418 460760
rect 368290 460748 368296 460760
rect 266412 460720 368296 460748
rect 266412 460708 266418 460720
rect 368290 460708 368296 460720
rect 368348 460708 368354 460760
rect 52362 460640 52368 460692
rect 52420 460680 52426 460692
rect 76006 460680 76012 460692
rect 52420 460652 76012 460680
rect 52420 460640 52426 460652
rect 76006 460640 76012 460652
rect 76064 460640 76070 460692
rect 193306 460640 193312 460692
rect 193364 460680 193370 460692
rect 208854 460680 208860 460692
rect 193364 460652 208860 460680
rect 193364 460640 193370 460652
rect 208854 460640 208860 460652
rect 208912 460640 208918 460692
rect 259454 460640 259460 460692
rect 259512 460680 259518 460692
rect 370958 460680 370964 460692
rect 259512 460652 370964 460680
rect 259512 460640 259518 460652
rect 370958 460640 370964 460652
rect 371016 460640 371022 460692
rect 55950 460572 55956 460624
rect 56008 460612 56014 460624
rect 77294 460612 77300 460624
rect 56008 460584 77300 460612
rect 56008 460572 56014 460584
rect 77294 460572 77300 460584
rect 77352 460572 77358 460624
rect 189074 460572 189080 460624
rect 189132 460612 189138 460624
rect 210326 460612 210332 460624
rect 189132 460584 210332 460612
rect 189132 460572 189138 460584
rect 210326 460572 210332 460584
rect 210384 460572 210390 460624
rect 249886 460572 249892 460624
rect 249944 460612 249950 460624
rect 362402 460612 362408 460624
rect 249944 460584 362408 460612
rect 249944 460572 249950 460584
rect 362402 460572 362408 460584
rect 362460 460572 362466 460624
rect 51534 460504 51540 460556
rect 51592 460544 51598 460556
rect 66346 460544 66352 460556
rect 51592 460516 66352 460544
rect 51592 460504 51598 460516
rect 66346 460504 66352 460516
rect 66404 460504 66410 460556
rect 169018 460504 169024 460556
rect 169076 460544 169082 460556
rect 197722 460544 197728 460556
rect 169076 460516 197728 460544
rect 169076 460504 169082 460516
rect 197722 460504 197728 460516
rect 197780 460504 197786 460556
rect 251174 460504 251180 460556
rect 251232 460544 251238 460556
rect 363966 460544 363972 460556
rect 251232 460516 363972 460544
rect 251232 460504 251238 460516
rect 363966 460504 363972 460516
rect 364024 460504 364030 460556
rect 47394 460436 47400 460488
rect 47452 460476 47458 460488
rect 63494 460476 63500 460488
rect 47452 460448 63500 460476
rect 47452 460436 47458 460448
rect 63494 460436 63500 460448
rect 63552 460436 63558 460488
rect 184934 460436 184940 460488
rect 184992 460476 184998 460488
rect 216214 460476 216220 460488
rect 184992 460448 216220 460476
rect 184992 460436 184998 460448
rect 216214 460436 216220 460448
rect 216272 460436 216278 460488
rect 249794 460436 249800 460488
rect 249852 460476 249858 460488
rect 368106 460476 368112 460488
rect 249852 460448 368112 460476
rect 249852 460436 249858 460448
rect 368106 460436 368112 460448
rect 368164 460436 368170 460488
rect 49602 460368 49608 460420
rect 49660 460408 49666 460420
rect 70394 460408 70400 460420
rect 49660 460380 70400 460408
rect 49660 460368 49666 460380
rect 70394 460368 70400 460380
rect 70452 460368 70458 460420
rect 179414 460368 179420 460420
rect 179472 460408 179478 460420
rect 214742 460408 214748 460420
rect 179472 460380 214748 460408
rect 179472 460368 179478 460380
rect 214742 460368 214748 460380
rect 214800 460368 214806 460420
rect 248414 460368 248420 460420
rect 248472 460408 248478 460420
rect 369394 460408 369400 460420
rect 248472 460380 369400 460408
rect 248472 460368 248478 460380
rect 369394 460368 369400 460380
rect 369452 460368 369458 460420
rect 41138 460300 41144 460352
rect 41196 460340 41202 460352
rect 71866 460340 71872 460352
rect 41196 460312 71872 460340
rect 41196 460300 41202 460312
rect 71866 460300 71872 460312
rect 71924 460300 71930 460352
rect 178126 460300 178132 460352
rect 178184 460340 178190 460352
rect 213546 460340 213552 460352
rect 178184 460312 213552 460340
rect 178184 460300 178190 460312
rect 213546 460300 213552 460312
rect 213604 460300 213610 460352
rect 244366 460300 244372 460352
rect 244424 460340 244430 460352
rect 366726 460340 366732 460352
rect 244424 460312 366732 460340
rect 244424 460300 244430 460312
rect 366726 460300 366732 460312
rect 366784 460300 366790 460352
rect 41230 460232 41236 460284
rect 41288 460272 41294 460284
rect 74534 460272 74540 460284
rect 41288 460244 74540 460272
rect 41288 460232 41294 460244
rect 74534 460232 74540 460244
rect 74592 460232 74598 460284
rect 164326 460232 164332 460284
rect 164384 460272 164390 460284
rect 218974 460272 218980 460284
rect 164384 460244 218980 460272
rect 164384 460232 164390 460244
rect 218974 460232 218980 460244
rect 219032 460232 219038 460284
rect 248506 460232 248512 460284
rect 248564 460272 248570 460284
rect 373350 460272 373356 460284
rect 248564 460244 373356 460272
rect 248564 460232 248570 460244
rect 373350 460232 373356 460244
rect 373408 460232 373414 460284
rect 43346 460164 43352 460216
rect 43404 460204 43410 460216
rect 68278 460204 68284 460216
rect 43404 460176 68284 460204
rect 43404 460164 43410 460176
rect 68278 460164 68284 460176
rect 68336 460164 68342 460216
rect 69658 460164 69664 460216
rect 69716 460204 69722 460216
rect 199010 460204 199016 460216
rect 69716 460176 199016 460204
rect 69716 460164 69722 460176
rect 199010 460164 199016 460176
rect 199068 460164 199074 460216
rect 247034 460164 247040 460216
rect 247092 460204 247098 460216
rect 378870 460204 378876 460216
rect 247092 460176 378876 460204
rect 247092 460164 247098 460176
rect 378870 460164 378876 460176
rect 378928 460164 378934 460216
rect 54478 460096 54484 460148
rect 54536 460136 54542 460148
rect 63586 460136 63592 460148
rect 54536 460108 63592 460136
rect 54536 460096 54542 460108
rect 63586 460096 63592 460108
rect 63644 460096 63650 460148
rect 278774 460096 278780 460148
rect 278832 460136 278838 460148
rect 362126 460136 362132 460148
rect 278832 460108 362132 460136
rect 278832 460096 278838 460108
rect 362126 460096 362132 460108
rect 362184 460096 362190 460148
rect 291194 460028 291200 460080
rect 291252 460068 291258 460080
rect 374454 460068 374460 460080
rect 291252 460040 374460 460068
rect 291252 460028 291258 460040
rect 374454 460028 374460 460040
rect 374512 460028 374518 460080
rect 288434 459960 288440 460012
rect 288492 460000 288498 460012
rect 357158 460000 357164 460012
rect 288492 459972 357164 460000
rect 288492 459960 288498 459972
rect 357158 459960 357164 459972
rect 357216 459960 357222 460012
rect 215202 459620 215208 459672
rect 215260 459660 215266 459672
rect 220998 459660 221004 459672
rect 215260 459632 221004 459660
rect 215260 459620 215266 459632
rect 220998 459620 221004 459632
rect 221056 459620 221062 459672
rect 216582 459552 216588 459604
rect 216640 459592 216646 459604
rect 220906 459592 220912 459604
rect 216640 459564 220912 459592
rect 216640 459552 216646 459564
rect 220906 459552 220912 459564
rect 220964 459552 220970 459604
rect 187694 459484 187700 459536
rect 187752 459524 187758 459536
rect 200942 459524 200948 459536
rect 187752 459496 200948 459524
rect 187752 459484 187758 459496
rect 200942 459484 200948 459496
rect 201000 459484 201006 459536
rect 295334 459484 295340 459536
rect 295392 459524 295398 459536
rect 370222 459524 370228 459536
rect 295392 459496 370228 459524
rect 295392 459484 295398 459496
rect 370222 459484 370228 459496
rect 370280 459484 370286 459536
rect 193214 459416 193220 459468
rect 193272 459456 193278 459468
rect 211614 459456 211620 459468
rect 193272 459428 211620 459456
rect 193272 459416 193278 459428
rect 211614 459416 211620 459428
rect 211672 459416 211678 459468
rect 281534 459416 281540 459468
rect 281592 459456 281598 459468
rect 359642 459456 359648 459468
rect 281592 459428 359648 459456
rect 281592 459416 281598 459428
rect 359642 459416 359648 459428
rect 359700 459416 359706 459468
rect 178034 459348 178040 459400
rect 178092 459388 178098 459400
rect 203702 459388 203708 459400
rect 178092 459360 203708 459388
rect 178092 459348 178098 459360
rect 203702 459348 203708 459360
rect 203760 459348 203766 459400
rect 276014 459348 276020 459400
rect 276072 459388 276078 459400
rect 358630 459388 358636 459400
rect 276072 459360 358636 459388
rect 276072 459348 276078 459360
rect 358630 459348 358636 459360
rect 358688 459348 358694 459400
rect 58894 459280 58900 459332
rect 58952 459320 58958 459332
rect 92474 459320 92480 459332
rect 58952 459292 92480 459320
rect 58952 459280 58958 459292
rect 92474 459280 92480 459292
rect 92532 459280 92538 459332
rect 180794 459280 180800 459332
rect 180852 459320 180858 459332
rect 209314 459320 209320 459332
rect 180852 459292 209320 459320
rect 180852 459280 180858 459292
rect 209314 459280 209320 459292
rect 209372 459280 209378 459332
rect 271874 459280 271880 459332
rect 271932 459320 271938 459332
rect 358722 459320 358728 459332
rect 271932 459292 358728 459320
rect 271932 459280 271938 459292
rect 358722 459280 358728 459292
rect 358780 459280 358786 459332
rect 55766 459212 55772 459264
rect 55824 459252 55830 459264
rect 103698 459252 103704 459264
rect 55824 459224 103704 459252
rect 55824 459212 55830 459224
rect 103698 459212 103704 459224
rect 103756 459212 103762 459264
rect 173894 459212 173900 459264
rect 173952 459252 173958 459264
rect 205266 459252 205272 459264
rect 173952 459224 205272 459252
rect 173952 459212 173958 459224
rect 205266 459212 205272 459224
rect 205324 459212 205330 459264
rect 256786 459212 256792 459264
rect 256844 459252 256850 459264
rect 361206 459252 361212 459264
rect 256844 459224 361212 459252
rect 256844 459212 256850 459224
rect 361206 459212 361212 459224
rect 361264 459212 361270 459264
rect 51626 459144 51632 459196
rect 51684 459184 51690 459196
rect 99466 459184 99472 459196
rect 51684 459156 99472 459184
rect 51684 459144 51690 459156
rect 99466 459144 99472 459156
rect 99524 459144 99530 459196
rect 173986 459144 173992 459196
rect 174044 459184 174050 459196
rect 219066 459184 219072 459196
rect 174044 459156 219072 459184
rect 174044 459144 174050 459156
rect 219066 459144 219072 459156
rect 219124 459144 219130 459196
rect 262214 459144 262220 459196
rect 262272 459184 262278 459196
rect 378962 459184 378968 459196
rect 262272 459156 378968 459184
rect 262272 459144 262278 459156
rect 378962 459144 378968 459156
rect 379020 459144 379026 459196
rect 53006 459076 53012 459128
rect 53064 459116 53070 459128
rect 100754 459116 100760 459128
rect 53064 459088 100760 459116
rect 53064 459076 53070 459088
rect 100754 459076 100760 459088
rect 100812 459076 100818 459128
rect 142246 459076 142252 459128
rect 142304 459116 142310 459128
rect 197906 459116 197912 459128
rect 142304 459088 197912 459116
rect 142304 459076 142310 459088
rect 197906 459076 197912 459088
rect 197964 459076 197970 459128
rect 256694 459076 256700 459128
rect 256752 459116 256758 459128
rect 373626 459116 373632 459128
rect 256752 459088 373632 459116
rect 256752 459076 256758 459088
rect 373626 459076 373632 459088
rect 373684 459076 373690 459128
rect 57790 459008 57796 459060
rect 57848 459048 57854 459060
rect 118878 459048 118884 459060
rect 57848 459020 118884 459048
rect 57848 459008 57854 459020
rect 118878 459008 118884 459020
rect 118936 459008 118942 459060
rect 142154 459008 142160 459060
rect 142212 459048 142218 459060
rect 199562 459048 199568 459060
rect 142212 459020 199568 459048
rect 142212 459008 142218 459020
rect 199562 459008 199568 459020
rect 199620 459008 199626 459060
rect 244274 459008 244280 459060
rect 244332 459048 244338 459060
rect 363874 459048 363880 459060
rect 244332 459020 363880 459048
rect 244332 459008 244338 459020
rect 363874 459008 363880 459020
rect 363932 459008 363938 459060
rect 54386 458940 54392 458992
rect 54444 458980 54450 458992
rect 121454 458980 121460 458992
rect 54444 458952 121460 458980
rect 54444 458940 54450 458952
rect 121454 458940 121460 458952
rect 121512 458940 121518 458992
rect 135438 458940 135444 458992
rect 135496 458980 135502 458992
rect 197814 458980 197820 458992
rect 135496 458952 197820 458980
rect 135496 458940 135502 458952
rect 197814 458940 197820 458952
rect 197872 458940 197878 458992
rect 245654 458940 245660 458992
rect 245712 458980 245718 458992
rect 379054 458980 379060 458992
rect 245712 458952 379060 458980
rect 245712 458940 245718 458952
rect 379054 458940 379060 458952
rect 379112 458940 379118 458992
rect 55950 458872 55956 458924
rect 56008 458912 56014 458924
rect 130010 458912 130016 458924
rect 56008 458884 130016 458912
rect 56008 458872 56014 458884
rect 130010 458872 130016 458884
rect 130068 458872 130074 458924
rect 136634 458872 136640 458924
rect 136692 458912 136698 458924
rect 199286 458912 199292 458924
rect 136692 458884 199292 458912
rect 136692 458872 136698 458884
rect 199286 458872 199292 458884
rect 199344 458872 199350 458924
rect 235994 458872 236000 458924
rect 236052 458912 236058 458924
rect 372154 458912 372160 458924
rect 236052 458884 372160 458912
rect 236052 458872 236058 458884
rect 372154 458872 372160 458884
rect 372212 458872 372218 458924
rect 54294 458804 54300 458856
rect 54352 458844 54358 458856
rect 134058 458844 134064 458856
rect 54352 458816 134064 458844
rect 54352 458804 54358 458816
rect 134058 458804 134064 458816
rect 134116 458804 134122 458856
rect 138014 458804 138020 458856
rect 138072 458844 138078 458856
rect 200666 458844 200672 458856
rect 138072 458816 200672 458844
rect 138072 458804 138078 458816
rect 200666 458804 200672 458816
rect 200724 458804 200730 458856
rect 223574 458804 223580 458856
rect 223632 458844 223638 458856
rect 365070 458844 365076 458856
rect 223632 458816 365076 458844
rect 223632 458804 223638 458816
rect 365070 458804 365076 458816
rect 365128 458804 365134 458856
rect 194594 458736 194600 458788
rect 194652 458776 194658 458788
rect 206186 458776 206192 458788
rect 194652 458748 206192 458776
rect 194652 458736 194658 458748
rect 206186 458736 206192 458748
rect 206244 458736 206250 458788
rect 292574 458736 292580 458788
rect 292632 458776 292638 458788
rect 366266 458776 366272 458788
rect 292632 458748 366272 458776
rect 292632 458736 292638 458748
rect 366266 458736 366272 458748
rect 366324 458736 366330 458788
rect 59262 458600 59268 458652
rect 59320 458640 59326 458652
rect 66254 458640 66260 458652
rect 59320 458612 66260 458640
rect 59320 458600 59326 458612
rect 66254 458600 66260 458612
rect 66312 458600 66318 458652
rect 199010 458328 199016 458380
rect 199068 458368 199074 458380
rect 199068 458340 354674 458368
rect 199068 458328 199074 458340
rect 48774 458260 48780 458312
rect 48832 458300 48838 458312
rect 354646 458300 354674 458340
rect 358906 458300 358912 458312
rect 48832 458272 200114 458300
rect 354646 458272 358912 458300
rect 48832 458260 48838 458272
rect 200086 458232 200114 458272
rect 358906 458260 358912 458272
rect 358964 458300 358970 458312
rect 516594 458300 516600 458312
rect 358964 458272 516600 458300
rect 358964 458260 358970 458272
rect 516594 458260 516600 458272
rect 516652 458260 516658 458312
rect 207382 458232 207388 458244
rect 200086 458204 207388 458232
rect 207382 458192 207388 458204
rect 207440 458232 207446 458244
rect 208118 458232 208124 458244
rect 207440 458204 208124 458232
rect 207440 458192 207446 458204
rect 208118 458192 208124 458204
rect 208176 458192 208182 458244
rect 205818 457444 205824 457496
rect 205876 457484 205882 457496
rect 217870 457484 217876 457496
rect 205876 457456 217876 457484
rect 205876 457444 205882 457456
rect 217870 457444 217876 457456
rect 217928 457444 217934 457496
rect 55858 457240 55864 457292
rect 55916 457280 55922 457292
rect 56410 457280 56416 457292
rect 55916 457252 56416 457280
rect 55916 457240 55922 457252
rect 56410 457240 56416 457252
rect 56468 457240 56474 457292
rect 48866 456084 48872 456136
rect 48924 456124 48930 456136
rect 49326 456124 49332 456136
rect 48924 456096 49332 456124
rect 48924 456084 48930 456096
rect 49326 456084 49332 456096
rect 49384 456084 49390 456136
rect 52914 456084 52920 456136
rect 52972 456124 52978 456136
rect 53282 456124 53288 456136
rect 52972 456096 53288 456124
rect 52972 456084 52978 456096
rect 53282 456084 53288 456096
rect 53340 456084 53346 456136
rect 519538 454656 519544 454708
rect 519596 454696 519602 454708
rect 580258 454696 580264 454708
rect 519596 454668 580264 454696
rect 519596 454656 519602 454668
rect 580258 454656 580264 454668
rect 580316 454656 580322 454708
rect 208118 417392 208124 417444
rect 208176 417432 208182 417444
rect 217778 417432 217784 417444
rect 208176 417404 217784 417432
rect 208176 417392 208182 417404
rect 217778 417392 217784 417404
rect 217836 417392 217842 417444
rect 203242 413924 203248 413976
rect 203300 413964 203306 413976
rect 206278 413964 206284 413976
rect 203300 413936 206284 413964
rect 203300 413924 203306 413936
rect 206278 413924 206284 413936
rect 206336 413924 206342 413976
rect 48866 412564 48872 412616
rect 48924 412604 48930 412616
rect 56962 412604 56968 412616
rect 48924 412576 56968 412604
rect 48924 412564 48930 412576
rect 56962 412564 56968 412576
rect 57020 412564 57026 412616
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 15838 411244 15844 411256
rect 3016 411216 15844 411244
rect 3016 411204 3022 411216
rect 15838 411204 15844 411216
rect 15896 411204 15902 411256
rect 44634 409844 44640 409896
rect 44692 409884 44698 409896
rect 57054 409884 57060 409896
rect 44692 409856 57060 409884
rect 44692 409844 44698 409856
rect 57054 409844 57060 409856
rect 57112 409844 57118 409896
rect 205726 409096 205732 409148
rect 205784 409136 205790 409148
rect 216766 409136 216772 409148
rect 205784 409108 216772 409136
rect 205784 409096 205790 409108
rect 216766 409096 216772 409108
rect 216824 409096 216830 409148
rect 360562 409096 360568 409148
rect 360620 409136 360626 409148
rect 377030 409136 377036 409148
rect 360620 409108 377036 409136
rect 360620 409096 360626 409108
rect 377030 409096 377036 409108
rect 377088 409096 377094 409148
rect 55674 408552 55680 408604
rect 55732 408592 55738 408604
rect 56962 408592 56968 408604
rect 55732 408564 56968 408592
rect 55732 408552 55738 408564
rect 56962 408552 56968 408564
rect 57020 408552 57026 408604
rect 46014 408484 46020 408536
rect 46072 408524 46078 408536
rect 57054 408524 57060 408536
rect 46072 408496 57060 408524
rect 46072 408484 46078 408496
rect 57054 408484 57060 408496
rect 57112 408484 57118 408536
rect 359918 407736 359924 407788
rect 359976 407776 359982 407788
rect 376754 407776 376760 407788
rect 359976 407748 376760 407776
rect 359976 407736 359982 407748
rect 376754 407736 376760 407748
rect 376812 407776 376818 407788
rect 376938 407776 376944 407788
rect 376812 407748 376944 407776
rect 376812 407736 376818 407748
rect 376938 407736 376944 407748
rect 376996 407736 377002 407788
rect 48866 407124 48872 407176
rect 48924 407164 48930 407176
rect 56962 407164 56968 407176
rect 48924 407136 56968 407164
rect 48924 407124 48930 407136
rect 56962 407124 56968 407136
rect 57020 407124 57026 407176
rect 357986 406376 357992 406428
rect 358044 406416 358050 406428
rect 377214 406416 377220 406428
rect 358044 406388 377220 406416
rect 358044 406376 358050 406388
rect 377214 406376 377220 406388
rect 377272 406376 377278 406428
rect 48774 405696 48780 405748
rect 48832 405736 48838 405748
rect 57054 405736 57060 405748
rect 48832 405708 57060 405736
rect 48832 405696 48838 405708
rect 57054 405696 57060 405708
rect 57112 405696 57118 405748
rect 377766 405628 377772 405680
rect 377824 405668 377830 405680
rect 378134 405668 378140 405680
rect 377824 405640 378140 405668
rect 377824 405628 377830 405640
rect 378134 405628 378140 405640
rect 378192 405628 378198 405680
rect 51626 404948 51632 405000
rect 51684 404988 51690 405000
rect 55858 404988 55864 405000
rect 51684 404960 55864 404988
rect 51684 404948 51690 404960
rect 55858 404948 55864 404960
rect 55916 404948 55922 405000
rect 204346 404948 204352 405000
rect 204404 404988 204410 405000
rect 216858 404988 216864 405000
rect 204404 404960 216864 404988
rect 204404 404948 204410 404960
rect 216858 404948 216864 404960
rect 216916 404948 216922 405000
rect 359826 404948 359832 405000
rect 359884 404988 359890 405000
rect 377306 404988 377312 405000
rect 359884 404960 377312 404988
rect 359884 404948 359890 404960
rect 377306 404948 377312 404960
rect 377364 404948 377370 405000
rect 51626 404336 51632 404388
rect 51684 404376 51690 404388
rect 57054 404376 57060 404388
rect 51684 404348 57060 404376
rect 51684 404336 51690 404348
rect 57054 404336 57060 404348
rect 57112 404336 57118 404388
rect 359734 403588 359740 403640
rect 359792 403628 359798 403640
rect 377766 403628 377772 403640
rect 359792 403600 377772 403628
rect 359792 403588 359798 403600
rect 377766 403588 377772 403600
rect 377824 403588 377830 403640
rect 52362 402976 52368 403028
rect 52420 403016 52426 403028
rect 57054 403016 57060 403028
rect 52420 402988 57060 403016
rect 52420 402976 52426 402988
rect 57054 402976 57060 402988
rect 57112 402976 57118 403028
rect 199654 393320 199660 393372
rect 199712 393360 199718 393372
rect 203242 393360 203248 393372
rect 199712 393332 203248 393360
rect 199712 393320 199718 393332
rect 203242 393320 203248 393332
rect 203300 393320 203306 393372
rect 199194 390872 199200 390924
rect 199252 390912 199258 390924
rect 199838 390912 199844 390924
rect 199252 390884 199844 390912
rect 199252 390872 199258 390884
rect 199838 390872 199844 390884
rect 199896 390872 199902 390924
rect 198090 390532 198096 390584
rect 198148 390572 198154 390584
rect 199102 390572 199108 390584
rect 198148 390544 199108 390572
rect 198148 390532 198154 390544
rect 199102 390532 199108 390544
rect 199160 390532 199166 390584
rect 198182 389172 198188 389224
rect 198240 389212 198246 389224
rect 199470 389212 199476 389224
rect 198240 389184 199476 389212
rect 198240 389172 198246 389184
rect 199470 389172 199476 389184
rect 199528 389172 199534 389224
rect 520918 388424 520924 388476
rect 520976 388464 520982 388476
rect 580350 388464 580356 388476
rect 520976 388436 580356 388464
rect 520976 388424 520982 388436
rect 580350 388424 580356 388436
rect 580408 388424 580414 388476
rect 44726 384956 44732 385008
rect 44784 384996 44790 385008
rect 56594 384996 56600 385008
rect 44784 384968 56600 384996
rect 44784 384956 44790 384968
rect 56594 384956 56600 384968
rect 56652 384956 56658 385008
rect 206278 384956 206284 385008
rect 206336 384996 206342 385008
rect 216950 384996 216956 385008
rect 206336 384968 216956 384996
rect 206336 384956 206342 384968
rect 216950 384956 216956 384968
rect 217008 384956 217014 385008
rect 359642 384956 359648 385008
rect 359700 384996 359706 385008
rect 376938 384996 376944 385008
rect 359700 384968 376944 384996
rect 359700 384956 359706 384968
rect 376938 384956 376944 384968
rect 376996 384956 377002 385008
rect 208210 384276 208216 384328
rect 208268 384316 208274 384328
rect 216674 384316 216680 384328
rect 208268 384288 216680 384316
rect 208268 384276 208274 384288
rect 216674 384276 216680 384288
rect 216732 384276 216738 384328
rect 57422 384208 57428 384260
rect 57480 384208 57486 384260
rect 57440 384056 57468 384208
rect 57422 384004 57428 384056
rect 57480 384004 57486 384056
rect 46106 383596 46112 383648
rect 46164 383636 46170 383648
rect 56594 383636 56600 383648
rect 46164 383608 56600 383636
rect 46164 383596 46170 383608
rect 56594 383596 56600 383608
rect 56652 383596 56658 383648
rect 57054 383596 57060 383648
rect 57112 383636 57118 383648
rect 57974 383636 57980 383648
rect 57112 383608 57980 383636
rect 57112 383596 57118 383608
rect 57974 383596 57980 383608
rect 58032 383596 58038 383648
rect 207014 383596 207020 383648
rect 207072 383636 207078 383648
rect 216674 383636 216680 383648
rect 207072 383608 216680 383636
rect 207072 383596 207078 383608
rect 216674 383596 216680 383608
rect 216732 383596 216738 383648
rect 359550 383596 359556 383648
rect 359608 383636 359614 383648
rect 376938 383636 376944 383648
rect 359608 383608 376944 383636
rect 359608 383596 359614 383608
rect 376938 383596 376944 383608
rect 376996 383596 377002 383648
rect 51718 383528 51724 383580
rect 51776 383568 51782 383580
rect 52914 383568 52920 383580
rect 51776 383540 52920 383568
rect 51776 383528 51782 383540
rect 52914 383528 52920 383540
rect 52972 383528 52978 383580
rect 202598 383528 202604 383580
rect 202656 383568 202662 383580
rect 217042 383568 217048 383580
rect 202656 383540 217048 383568
rect 202656 383528 202662 383540
rect 217042 383528 217048 383540
rect 217100 383528 217106 383580
rect 206278 382236 206284 382288
rect 206336 382276 206342 382288
rect 207014 382276 207020 382288
rect 206336 382248 207020 382276
rect 206336 382236 206342 382248
rect 207014 382236 207020 382248
rect 207072 382236 207078 382288
rect 41322 382168 41328 382220
rect 41380 382208 41386 382220
rect 57238 382208 57244 382220
rect 41380 382180 57244 382208
rect 41380 382168 41386 382180
rect 57238 382168 57244 382180
rect 57296 382168 57302 382220
rect 367738 382168 367744 382220
rect 367796 382208 367802 382220
rect 375374 382208 375380 382220
rect 367796 382180 375380 382208
rect 367796 382168 367802 382180
rect 375374 382168 375380 382180
rect 375432 382208 375438 382220
rect 376662 382208 376668 382220
rect 375432 382180 376668 382208
rect 375432 382168 375438 382180
rect 376662 382168 376668 382180
rect 376720 382168 376726 382220
rect 56042 380808 56048 380860
rect 56100 380848 56106 380860
rect 57054 380848 57060 380860
rect 56100 380820 57060 380848
rect 56100 380808 56106 380820
rect 57054 380808 57060 380820
rect 57112 380808 57118 380860
rect 57330 378768 57336 378820
rect 57388 378808 57394 378820
rect 57514 378808 57520 378820
rect 57388 378780 57520 378808
rect 57388 378768 57394 378780
rect 57514 378768 57520 378780
rect 57572 378768 57578 378820
rect 373994 378768 374000 378820
rect 374052 378808 374058 378820
rect 374362 378808 374368 378820
rect 374052 378780 374368 378808
rect 374052 378768 374058 378780
rect 374362 378768 374368 378780
rect 374420 378768 374426 378820
rect 57146 378632 57152 378684
rect 57204 378672 57210 378684
rect 57330 378672 57336 378684
rect 57204 378644 57336 378672
rect 57204 378632 57210 378644
rect 57330 378632 57336 378644
rect 57388 378632 57394 378684
rect 55766 375300 55772 375352
rect 55824 375340 55830 375352
rect 59354 375340 59360 375352
rect 55824 375312 59360 375340
rect 55824 375300 55830 375312
rect 59354 375300 59360 375312
rect 59412 375300 59418 375352
rect 217226 375300 217232 375352
rect 217284 375340 217290 375352
rect 217870 375340 217876 375352
rect 217284 375312 217876 375340
rect 217284 375300 217290 375312
rect 217870 375300 217876 375312
rect 217928 375300 217934 375352
rect 377858 375300 377864 375352
rect 377916 375340 377922 375352
rect 379238 375340 379244 375352
rect 377916 375312 379244 375340
rect 377916 375300 377922 375312
rect 379238 375300 379244 375312
rect 379296 375300 379302 375352
rect 48866 375028 48872 375080
rect 48924 375068 48930 375080
rect 217226 375068 217232 375080
rect 48924 375040 217232 375068
rect 48924 375028 48930 375040
rect 217226 375028 217232 375040
rect 217284 375028 217290 375080
rect 51626 374960 51632 375012
rect 51684 375000 51690 375012
rect 216950 375000 216956 375012
rect 51684 374972 216956 375000
rect 51684 374960 51690 374972
rect 216950 374960 216956 374972
rect 217008 374960 217014 375012
rect 379422 374960 379428 375012
rect 379480 375000 379486 375012
rect 380894 375000 380900 375012
rect 379480 374972 380900 375000
rect 379480 374960 379486 374972
rect 380894 374960 380900 374972
rect 380952 374960 380958 375012
rect 54386 374824 54392 374876
rect 54444 374864 54450 374876
rect 56594 374864 56600 374876
rect 54444 374836 56600 374864
rect 54444 374824 54450 374836
rect 56594 374824 56600 374836
rect 56652 374824 56658 374876
rect 201494 374824 201500 374876
rect 201552 374864 201558 374876
rect 275278 374864 275284 374876
rect 201552 374836 275284 374864
rect 201552 374824 201558 374836
rect 275278 374824 275284 374836
rect 275336 374824 275342 374876
rect 200206 374756 200212 374808
rect 200264 374796 200270 374808
rect 295334 374796 295340 374808
rect 200264 374768 295340 374796
rect 200264 374756 200270 374768
rect 295334 374756 295340 374768
rect 295392 374756 295398 374808
rect 201034 374688 201040 374740
rect 201092 374728 201098 374740
rect 304994 374728 305000 374740
rect 201092 374700 305000 374728
rect 201092 374688 201098 374700
rect 304994 374688 305000 374700
rect 305052 374688 305058 374740
rect 356882 374688 356888 374740
rect 356940 374728 356946 374740
rect 452838 374728 452844 374740
rect 356940 374700 452844 374728
rect 356940 374688 356946 374700
rect 452838 374688 452844 374700
rect 452896 374688 452902 374740
rect 53650 374620 53656 374672
rect 53708 374660 53714 374672
rect 59630 374660 59636 374672
rect 53708 374632 59636 374660
rect 53708 374620 53714 374632
rect 59630 374620 59636 374632
rect 59688 374620 59694 374672
rect 203058 374620 203064 374672
rect 203116 374660 203122 374672
rect 312814 374660 312820 374672
rect 203116 374632 312820 374660
rect 203116 374620 203122 374632
rect 312814 374620 312820 374632
rect 312872 374620 312878 374672
rect 165982 374552 165988 374604
rect 166040 374592 166046 374604
rect 199562 374592 199568 374604
rect 166040 374564 199568 374592
rect 166040 374552 166046 374564
rect 199562 374552 199568 374564
rect 199620 374552 199626 374604
rect 379238 374552 379244 374604
rect 379296 374592 379302 374604
rect 425054 374592 425060 374604
rect 379296 374564 425060 374592
rect 379296 374552 379302 374564
rect 425054 374552 425060 374564
rect 425112 374552 425118 374604
rect 163406 374484 163412 374536
rect 163464 374524 163470 374536
rect 197906 374524 197912 374536
rect 163464 374496 197912 374524
rect 163464 374484 163470 374496
rect 197906 374484 197912 374496
rect 197964 374484 197970 374536
rect 203150 374484 203156 374536
rect 203208 374524 203214 374536
rect 213914 374524 213920 374536
rect 203208 374496 213920 374524
rect 203208 374484 203214 374496
rect 213914 374484 213920 374496
rect 213972 374484 213978 374536
rect 362862 374484 362868 374536
rect 362920 374524 362926 374536
rect 410702 374524 410708 374536
rect 362920 374496 410708 374524
rect 362920 374484 362926 374496
rect 410702 374484 410708 374496
rect 410760 374484 410766 374536
rect 158530 374416 158536 374468
rect 158588 374456 158594 374468
rect 201770 374456 201776 374468
rect 158588 374428 201776 374456
rect 158588 374416 158594 374428
rect 201770 374416 201776 374428
rect 201828 374416 201834 374468
rect 209498 374416 209504 374468
rect 209556 374456 209562 374468
rect 320910 374456 320916 374468
rect 209556 374428 320916 374456
rect 209556 374416 209562 374428
rect 320910 374416 320916 374428
rect 320968 374416 320974 374468
rect 359458 374416 359464 374468
rect 359516 374456 359522 374468
rect 407758 374456 407764 374468
rect 359516 374428 407764 374456
rect 359516 374416 359522 374428
rect 407758 374416 407764 374428
rect 407816 374416 407822 374468
rect 153470 374348 153476 374400
rect 153528 374388 153534 374400
rect 200574 374388 200580 374400
rect 153528 374360 200580 374388
rect 153528 374348 153534 374360
rect 200574 374348 200580 374360
rect 200632 374348 200638 374400
rect 210234 374348 210240 374400
rect 210292 374388 210298 374400
rect 210786 374388 210792 374400
rect 210292 374360 210792 374388
rect 210292 374348 210298 374360
rect 210786 374348 210792 374360
rect 210844 374388 210850 374400
rect 244274 374388 244280 374400
rect 210844 374360 244280 374388
rect 210844 374348 210850 374360
rect 244274 374348 244280 374360
rect 244332 374348 244338 374400
rect 372430 374348 372436 374400
rect 372488 374388 372494 374400
rect 438486 374388 438492 374400
rect 372488 374360 438492 374388
rect 372488 374348 372494 374360
rect 438486 374348 438492 374360
rect 438544 374348 438550 374400
rect 160922 374280 160928 374332
rect 160980 374320 160986 374332
rect 208486 374320 208492 374332
rect 160980 374292 208492 374320
rect 160980 374280 160986 374292
rect 208486 374280 208492 374292
rect 208544 374280 208550 374332
rect 369762 374280 369768 374332
rect 369820 374320 369826 374332
rect 440326 374320 440332 374332
rect 369820 374292 440332 374320
rect 369820 374280 369826 374292
rect 440326 374280 440332 374292
rect 440384 374280 440390 374332
rect 156506 374212 156512 374264
rect 156564 374252 156570 374264
rect 204530 374252 204536 374264
rect 156564 374224 204536 374252
rect 156564 374212 156570 374224
rect 204530 374212 204536 374224
rect 204588 374212 204594 374264
rect 217502 374212 217508 374264
rect 217560 374252 217566 374264
rect 256050 374252 256056 374264
rect 217560 374224 256056 374252
rect 217560 374212 217566 374224
rect 256050 374212 256056 374224
rect 256108 374212 256114 374264
rect 360746 374212 360752 374264
rect 360804 374252 360810 374264
rect 436002 374252 436008 374264
rect 360804 374224 436008 374252
rect 360804 374212 360810 374224
rect 436002 374212 436008 374224
rect 436060 374212 436066 374264
rect 58618 374144 58624 374196
rect 58676 374184 58682 374196
rect 93578 374184 93584 374196
rect 58676 374156 93584 374184
rect 58676 374144 58682 374156
rect 93578 374144 93584 374156
rect 93636 374144 93642 374196
rect 148962 374144 148968 374196
rect 149020 374184 149026 374196
rect 197078 374184 197084 374196
rect 149020 374156 197084 374184
rect 149020 374144 149026 374156
rect 197078 374144 197084 374156
rect 197136 374144 197142 374196
rect 199378 374144 199384 374196
rect 199436 374184 199442 374196
rect 250714 374184 250720 374196
rect 199436 374156 250720 374184
rect 199436 374144 199442 374156
rect 250714 374144 250720 374156
rect 250772 374144 250778 374196
rect 358722 374144 358728 374196
rect 358780 374184 358786 374196
rect 433610 374184 433616 374196
rect 358780 374156 433616 374184
rect 358780 374144 358786 374156
rect 433610 374144 433616 374156
rect 433668 374144 433674 374196
rect 56962 374076 56968 374128
rect 57020 374116 57026 374128
rect 103514 374116 103520 374128
rect 57020 374088 103520 374116
rect 57020 374076 57026 374088
rect 103514 374076 103520 374088
rect 103572 374076 103578 374128
rect 146202 374076 146208 374128
rect 146260 374116 146266 374128
rect 207474 374116 207480 374128
rect 146260 374088 207480 374116
rect 146260 374076 146266 374088
rect 207474 374076 207480 374088
rect 207532 374076 207538 374128
rect 241054 374076 241060 374128
rect 241112 374116 241118 374128
rect 250070 374116 250076 374128
rect 241112 374088 250076 374116
rect 241112 374076 241118 374088
rect 250070 374076 250076 374088
rect 250128 374076 250134 374128
rect 366174 374076 366180 374128
rect 366232 374116 366238 374128
rect 443086 374116 443092 374128
rect 366232 374088 443092 374116
rect 366232 374076 366238 374088
rect 443086 374076 443092 374088
rect 443144 374076 443150 374128
rect 54294 374008 54300 374060
rect 54352 374048 54358 374060
rect 116026 374048 116032 374060
rect 54352 374020 116032 374048
rect 54352 374008 54358 374020
rect 116026 374008 116032 374020
rect 116084 374008 116090 374060
rect 143534 374008 143540 374060
rect 143592 374048 143598 374060
rect 205910 374048 205916 374060
rect 143592 374020 205916 374048
rect 143592 374008 143598 374020
rect 205910 374008 205916 374020
rect 205968 374008 205974 374060
rect 213914 374008 213920 374060
rect 213972 374048 213978 374060
rect 215110 374048 215116 374060
rect 213972 374020 215116 374048
rect 213972 374008 213978 374020
rect 215110 374008 215116 374020
rect 215168 374048 215174 374060
rect 235994 374048 236000 374060
rect 215168 374020 236000 374048
rect 215168 374008 215174 374020
rect 235994 374008 236000 374020
rect 236052 374008 236058 374060
rect 380894 374008 380900 374060
rect 380952 374048 380958 374060
rect 405918 374048 405924 374060
rect 380952 374020 405924 374048
rect 380952 374008 380958 374020
rect 405918 374008 405924 374020
rect 405976 374008 405982 374060
rect 44634 373940 44640 373992
rect 44692 373980 44698 373992
rect 217686 373980 217692 373992
rect 44692 373952 217692 373980
rect 44692 373940 44698 373952
rect 217686 373940 217692 373952
rect 217744 373940 217750 373992
rect 48774 373872 48780 373924
rect 48832 373912 48838 373924
rect 217502 373912 217508 373924
rect 48832 373884 217508 373912
rect 48832 373872 48838 373884
rect 217502 373872 217508 373884
rect 217560 373872 217566 373924
rect 40770 373804 40776 373856
rect 40828 373844 40834 373856
rect 199102 373844 199108 373856
rect 40828 373816 199108 373844
rect 40828 373804 40834 373816
rect 199102 373804 199108 373816
rect 199160 373804 199166 373856
rect 375282 373804 375288 373856
rect 375340 373844 375346 373856
rect 416038 373844 416044 373856
rect 375340 373816 416044 373844
rect 375340 373804 375346 373816
rect 416038 373804 416044 373816
rect 416096 373804 416102 373856
rect 59722 373736 59728 373788
rect 59780 373776 59786 373788
rect 107838 373776 107844 373788
rect 59780 373748 107844 373776
rect 59780 373736 59786 373748
rect 107838 373736 107844 373748
rect 107896 373736 107902 373788
rect 136450 373736 136456 373788
rect 136508 373776 136514 373788
rect 200482 373776 200488 373788
rect 136508 373748 200488 373776
rect 136508 373736 136514 373748
rect 200482 373736 200488 373748
rect 200540 373736 200546 373788
rect 215294 373736 215300 373788
rect 215352 373776 215358 373788
rect 217870 373776 217876 373788
rect 215352 373748 217876 373776
rect 215352 373736 215358 373748
rect 217870 373736 217876 373748
rect 217928 373736 217934 373788
rect 375926 373736 375932 373788
rect 375984 373776 375990 373788
rect 418246 373776 418252 373788
rect 375984 373748 418252 373776
rect 375984 373736 375990 373748
rect 418246 373736 418252 373748
rect 418304 373736 418310 373788
rect 42334 373668 42340 373720
rect 42392 373708 42398 373720
rect 100846 373708 100852 373720
rect 42392 373680 100852 373708
rect 42392 373668 42398 373680
rect 100846 373668 100852 373680
rect 100904 373668 100910 373720
rect 131022 373668 131028 373720
rect 131080 373708 131086 373720
rect 199286 373708 199292 373720
rect 131080 373680 199292 373708
rect 131080 373668 131086 373680
rect 199286 373668 199292 373680
rect 199344 373668 199350 373720
rect 371786 373668 371792 373720
rect 371844 373708 371850 373720
rect 423030 373708 423036 373720
rect 371844 373680 423036 373708
rect 371844 373668 371850 373680
rect 423030 373668 423036 373680
rect 423088 373668 423094 373720
rect 57054 373600 57060 373652
rect 57112 373640 57118 373652
rect 118326 373640 118332 373652
rect 57112 373612 118332 373640
rect 57112 373600 57118 373612
rect 118326 373600 118332 373612
rect 118384 373600 118390 373652
rect 128906 373600 128912 373652
rect 128964 373640 128970 373652
rect 198182 373640 198188 373652
rect 128964 373612 198188 373640
rect 128964 373600 128970 373612
rect 198182 373600 198188 373612
rect 198240 373600 198246 373652
rect 204254 373600 204260 373652
rect 204312 373640 204318 373652
rect 215294 373640 215300 373652
rect 204312 373612 215300 373640
rect 204312 373600 204318 373612
rect 215294 373600 215300 373612
rect 215352 373600 215358 373652
rect 369762 373600 369768 373652
rect 369820 373640 369826 373652
rect 375466 373640 375472 373652
rect 369820 373612 375472 373640
rect 369820 373600 369826 373612
rect 375466 373600 375472 373612
rect 375524 373640 375530 373652
rect 426894 373640 426900 373652
rect 375524 373612 426900 373640
rect 375524 373600 375530 373612
rect 426894 373600 426900 373612
rect 426952 373600 426958 373652
rect 52270 373532 52276 373584
rect 52328 373572 52334 373584
rect 113542 373572 113548 373584
rect 52328 373544 113548 373572
rect 52328 373532 52334 373544
rect 113542 373532 113548 373544
rect 113600 373532 113606 373584
rect 133690 373532 133696 373584
rect 133748 373572 133754 373584
rect 204438 373572 204444 373584
rect 133748 373544 204444 373572
rect 133748 373532 133754 373544
rect 204438 373532 204444 373544
rect 204496 373532 204502 373584
rect 368382 373532 368388 373584
rect 368440 373572 368446 373584
rect 445846 373572 445852 373584
rect 368440 373544 445852 373572
rect 368440 373532 368446 373544
rect 445846 373532 445852 373544
rect 445904 373532 445910 373584
rect 48958 373464 48964 373516
rect 49016 373504 49022 373516
rect 110414 373504 110420 373516
rect 49016 373476 110420 373504
rect 49016 373464 49022 373476
rect 110414 373464 110420 373476
rect 110472 373464 110478 373516
rect 125778 373464 125784 373516
rect 125836 373504 125842 373516
rect 201678 373504 201684 373516
rect 125836 373476 201684 373504
rect 125836 373464 125842 373476
rect 201678 373464 201684 373476
rect 201736 373464 201742 373516
rect 214374 373464 214380 373516
rect 214432 373504 214438 373516
rect 224218 373504 224224 373516
rect 214432 373476 224224 373504
rect 214432 373464 214438 373476
rect 224218 373464 224224 373476
rect 224276 373464 224282 373516
rect 370406 373464 370412 373516
rect 370464 373504 370470 373516
rect 450262 373504 450268 373516
rect 370464 373476 450268 373504
rect 370464 373464 370470 373476
rect 450262 373464 450268 373476
rect 450320 373464 450326 373516
rect 43254 373396 43260 373448
rect 43312 373436 43318 373448
rect 105446 373436 105452 373448
rect 43312 373408 105452 373436
rect 43312 373396 43318 373408
rect 105446 373396 105452 373408
rect 105504 373396 105510 373448
rect 121362 373396 121368 373448
rect 121420 373436 121426 373448
rect 197814 373436 197820 373448
rect 121420 373408 197820 373436
rect 121420 373396 121426 373408
rect 197814 373396 197820 373408
rect 197872 373396 197878 373448
rect 210142 373396 210148 373448
rect 210200 373436 210206 373448
rect 212534 373436 212540 373448
rect 210200 373408 212540 373436
rect 210200 373396 210206 373408
rect 212534 373396 212540 373408
rect 212592 373436 212598 373448
rect 256694 373436 256700 373448
rect 212592 373408 256700 373436
rect 212592 373396 212598 373408
rect 256694 373396 256700 373408
rect 256752 373396 256758 373448
rect 373718 373396 373724 373448
rect 373776 373436 373782 373448
rect 455414 373436 455420 373448
rect 373776 373408 455420 373436
rect 373776 373396 373782 373408
rect 455414 373396 455420 373408
rect 455472 373396 455478 373448
rect 50154 373328 50160 373380
rect 50212 373368 50218 373380
rect 98270 373368 98276 373380
rect 50212 373340 98276 373368
rect 50212 373328 50218 373340
rect 98270 373328 98276 373340
rect 98328 373328 98334 373380
rect 99374 373328 99380 373380
rect 99432 373368 99438 373380
rect 204254 373368 204260 373380
rect 99432 373340 204260 373368
rect 99432 373328 99438 373340
rect 204254 373328 204260 373340
rect 204312 373328 204318 373380
rect 213086 373328 213092 373380
rect 213144 373368 213150 373380
rect 214098 373368 214104 373380
rect 213144 373340 214104 373368
rect 213144 373328 213150 373340
rect 214098 373328 214104 373340
rect 214156 373368 214162 373380
rect 260006 373368 260012 373380
rect 214156 373340 260012 373368
rect 214156 373328 214162 373340
rect 260006 373328 260012 373340
rect 260064 373328 260070 373380
rect 363414 373328 363420 373380
rect 363472 373368 363478 373380
rect 447686 373368 447692 373380
rect 363472 373340 447692 373368
rect 363472 373328 363478 373340
rect 447686 373328 447692 373340
rect 447744 373328 447750 373380
rect 57330 373260 57336 373312
rect 57388 373300 57394 373312
rect 122926 373300 122932 373312
rect 57388 373272 122932 373300
rect 57388 373260 57394 373272
rect 122926 373260 122932 373272
rect 122984 373260 122990 373312
rect 191742 373260 191748 373312
rect 191800 373300 191806 373312
rect 206278 373300 206284 373312
rect 191800 373272 206284 373300
rect 191800 373260 191806 373272
rect 206278 373260 206284 373272
rect 206336 373260 206342 373312
rect 262858 373260 262864 373312
rect 262916 373300 262922 373312
rect 269206 373300 269212 373312
rect 262916 373272 269212 373300
rect 262916 373260 262922 373272
rect 269206 373260 269212 373272
rect 269264 373260 269270 373312
rect 358630 373260 358636 373312
rect 358688 373300 358694 373312
rect 462774 373300 462780 373312
rect 358688 373272 462780 373300
rect 358688 373260 358694 373272
rect 462774 373260 462780 373272
rect 462832 373260 462838 373312
rect 49050 373192 49056 373244
rect 49108 373232 49114 373244
rect 96062 373232 96068 373244
rect 49108 373204 96068 373232
rect 49108 373192 49114 373204
rect 96062 373192 96068 373204
rect 96120 373192 96126 373244
rect 139210 373192 139216 373244
rect 139268 373232 139274 373244
rect 200666 373232 200672 373244
rect 139268 373204 200672 373232
rect 139268 373192 139274 373204
rect 200666 373192 200672 373204
rect 200724 373192 200730 373244
rect 215294 373192 215300 373244
rect 215352 373232 215358 373244
rect 216490 373232 216496 373244
rect 215352 373204 216496 373232
rect 215352 373192 215358 373204
rect 216490 373192 216496 373204
rect 216548 373232 216554 373244
rect 236454 373232 236460 373244
rect 216548 373204 236460 373232
rect 216548 373192 216554 373204
rect 236454 373192 236460 373204
rect 236512 373192 236518 373244
rect 47578 373124 47584 373176
rect 47636 373164 47642 373176
rect 88334 373164 88340 373176
rect 47636 373136 88340 373164
rect 47636 373124 47642 373136
rect 88334 373124 88340 373136
rect 88392 373124 88398 373176
rect 141602 373124 141608 373176
rect 141660 373164 141666 373176
rect 203334 373164 203340 373176
rect 141660 373136 203340 373164
rect 141660 373124 141666 373136
rect 203334 373124 203340 373136
rect 203392 373124 203398 373176
rect 207198 373124 207204 373176
rect 207256 373164 207262 373176
rect 213730 373164 213736 373176
rect 207256 373136 213736 373164
rect 207256 373124 207262 373136
rect 213730 373124 213736 373136
rect 213788 373164 213794 373176
rect 242894 373164 242900 373176
rect 213788 373136 242900 373164
rect 213788 373124 213794 373136
rect 242894 373124 242900 373136
rect 242952 373124 242958 373176
rect 55950 373056 55956 373108
rect 56008 373096 56014 373108
rect 90174 373096 90180 373108
rect 56008 373068 90180 373096
rect 56008 373056 56014 373068
rect 90174 373056 90180 373068
rect 90232 373056 90238 373108
rect 151722 373056 151728 373108
rect 151780 373096 151786 373108
rect 198090 373096 198096 373108
rect 151780 373068 198096 373096
rect 151780 373056 151786 373068
rect 198090 373056 198096 373068
rect 198148 373056 198154 373108
rect 220722 373056 220728 373108
rect 220780 373096 220786 373108
rect 253934 373096 253940 373108
rect 220780 373068 253940 373096
rect 220780 373056 220786 373068
rect 253934 373056 253940 373068
rect 253992 373056 253998 373108
rect 42242 372988 42248 373040
rect 42300 373028 42306 373040
rect 59722 373028 59728 373040
rect 42300 373000 59728 373028
rect 42300 372988 42306 373000
rect 59722 372988 59728 373000
rect 59780 372988 59786 373040
rect 212626 372988 212632 373040
rect 212684 373028 212690 373040
rect 217962 373028 217968 373040
rect 212684 373000 217968 373028
rect 212684 372988 212690 373000
rect 217962 372988 217968 373000
rect 218020 373028 218026 373040
rect 255406 373028 255412 373040
rect 218020 373000 255412 373028
rect 218020 372988 218026 373000
rect 255406 372988 255412 373000
rect 255464 372988 255470 373040
rect 213914 372920 213920 372972
rect 213972 372960 213978 372972
rect 219342 372960 219348 372972
rect 213972 372932 219348 372960
rect 213972 372920 213978 372932
rect 219342 372920 219348 372932
rect 219400 372960 219406 372972
rect 261294 372960 261300 372972
rect 219400 372932 261300 372960
rect 219400 372920 219406 372932
rect 261294 372920 261300 372932
rect 261352 372920 261358 372972
rect 212810 372852 212816 372904
rect 212868 372892 212874 372904
rect 217134 372892 217140 372904
rect 212868 372864 217140 372892
rect 212868 372852 212874 372864
rect 217134 372852 217140 372864
rect 217192 372892 217198 372904
rect 258074 372892 258080 372904
rect 217192 372864 258080 372892
rect 217192 372852 217198 372864
rect 258074 372852 258080 372864
rect 258132 372852 258138 372904
rect 214006 372784 214012 372836
rect 214064 372824 214070 372836
rect 259454 372824 259460 372836
rect 214064 372796 259460 372824
rect 214064 372784 214070 372796
rect 259454 372784 259460 372796
rect 259512 372784 259518 372836
rect 215386 372716 215392 372768
rect 215444 372756 215450 372768
rect 262214 372756 262220 372768
rect 215444 372728 262220 372756
rect 215444 372716 215450 372728
rect 262214 372716 262220 372728
rect 262272 372716 262278 372768
rect 379146 372716 379152 372768
rect 379204 372756 379210 372768
rect 379790 372756 379796 372768
rect 379204 372728 379796 372756
rect 379204 372716 379210 372728
rect 379790 372716 379796 372728
rect 379848 372716 379854 372768
rect 217870 372648 217876 372700
rect 217928 372688 217934 372700
rect 264974 372688 264980 372700
rect 217928 372660 264980 372688
rect 217928 372648 217934 372660
rect 264974 372648 264980 372660
rect 265032 372648 265038 372700
rect 211154 372580 211160 372632
rect 211212 372580 211218 372632
rect 217042 372580 217048 372632
rect 217100 372620 217106 372632
rect 217686 372620 217692 372632
rect 217100 372592 217692 372620
rect 217100 372580 217106 372592
rect 217686 372580 217692 372592
rect 217744 372580 217750 372632
rect 219250 372580 219256 372632
rect 219308 372620 219314 372632
rect 266354 372620 266360 372632
rect 219308 372592 266360 372620
rect 219308 372580 219314 372592
rect 266354 372580 266360 372592
rect 266412 372580 266418 372632
rect 362862 372580 362868 372632
rect 362920 372620 362926 372632
rect 371234 372620 371240 372632
rect 362920 372592 371240 372620
rect 362920 372580 362926 372592
rect 371234 372580 371240 372592
rect 371292 372580 371298 372632
rect 379790 372580 379796 372632
rect 379848 372620 379854 372632
rect 402882 372620 402888 372632
rect 379848 372592 402888 372620
rect 379848 372580 379854 372592
rect 402882 372580 402888 372592
rect 402940 372580 402946 372632
rect 84746 372512 84752 372564
rect 84804 372552 84810 372564
rect 208394 372552 208400 372564
rect 84804 372524 208400 372552
rect 84804 372512 84810 372524
rect 208394 372512 208400 372524
rect 208452 372512 208458 372564
rect 210970 372512 210976 372564
rect 211028 372552 211034 372564
rect 211172 372552 211200 372580
rect 211028 372524 211200 372552
rect 211028 372512 211034 372524
rect 212350 372512 212356 372564
rect 212408 372552 212414 372564
rect 218054 372552 218060 372564
rect 212408 372524 218060 372552
rect 212408 372512 212414 372524
rect 218054 372512 218060 372524
rect 218112 372552 218118 372564
rect 271874 372552 271880 372564
rect 218112 372524 271880 372552
rect 218112 372512 218118 372524
rect 271874 372512 271880 372524
rect 271932 372512 271938 372564
rect 275278 372512 275284 372564
rect 275336 372552 275342 372564
rect 314654 372552 314660 372564
rect 275336 372524 314660 372552
rect 275336 372512 275342 372524
rect 314654 372512 314660 372524
rect 314712 372512 314718 372564
rect 373166 372512 373172 372564
rect 373224 372552 373230 372564
rect 377398 372552 377404 372564
rect 373224 372524 377404 372552
rect 373224 372512 373230 372524
rect 377398 372512 377404 372524
rect 377456 372512 377462 372564
rect 86770 372444 86776 372496
rect 86828 372484 86834 372496
rect 208210 372484 208216 372496
rect 86828 372456 208216 372484
rect 86828 372444 86834 372456
rect 208210 372444 208216 372456
rect 208268 372444 208274 372496
rect 208412 372484 208440 372512
rect 215018 372484 215024 372496
rect 208412 372456 215024 372484
rect 215018 372444 215024 372456
rect 215076 372484 215082 372496
rect 215076 372456 219434 372484
rect 215076 372444 215082 372456
rect 89346 372376 89352 372428
rect 89404 372416 89410 372428
rect 209774 372416 209780 372428
rect 89404 372388 209780 372416
rect 89404 372376 89410 372388
rect 209774 372376 209780 372388
rect 209832 372416 209838 372428
rect 210050 372416 210056 372428
rect 209832 372388 210056 372416
rect 209832 372376 209838 372388
rect 210050 372376 210056 372388
rect 210108 372376 210114 372428
rect 219406 372416 219434 372456
rect 295334 372444 295340 372496
rect 295392 372484 295398 372496
rect 310514 372484 310520 372496
rect 295392 372456 310520 372484
rect 295392 372444 295398 372456
rect 310514 372444 310520 372456
rect 310572 372444 310578 372496
rect 312814 372444 312820 372496
rect 312872 372484 312878 372496
rect 322934 372484 322940 372496
rect 312872 372456 322940 372484
rect 312872 372444 312878 372456
rect 322934 372444 322940 372456
rect 322992 372444 322998 372496
rect 244274 372416 244280 372428
rect 219406 372388 244280 372416
rect 244274 372376 244280 372388
rect 244332 372376 244338 372428
rect 304994 372376 305000 372428
rect 305052 372416 305058 372428
rect 313274 372416 313280 372428
rect 305052 372388 313280 372416
rect 305052 372376 305058 372388
rect 313274 372376 313280 372388
rect 313332 372376 313338 372428
rect 92382 372308 92388 372360
rect 92440 372348 92446 372360
rect 211246 372348 211252 372360
rect 92440 372320 211252 372348
rect 92440 372308 92446 372320
rect 211246 372308 211252 372320
rect 211304 372308 211310 372360
rect 372890 372308 372896 372360
rect 372948 372348 372954 372360
rect 400214 372348 400220 372360
rect 372948 372320 400220 372348
rect 372948 372308 372954 372320
rect 400214 372308 400220 372320
rect 400272 372308 400278 372360
rect 77202 372240 77208 372292
rect 77260 372280 77266 372292
rect 99374 372280 99380 372292
rect 77260 372252 99380 372280
rect 77260 372240 77266 372252
rect 99374 372240 99380 372252
rect 99432 372240 99438 372292
rect 114462 372240 114468 372292
rect 114520 372280 114526 372292
rect 219434 372280 219440 372292
rect 114520 372252 219440 372280
rect 114520 372240 114526 372252
rect 219434 372240 219440 372252
rect 219492 372280 219498 372292
rect 220722 372280 220728 372292
rect 219492 372252 220728 372280
rect 219492 372240 219498 372252
rect 220722 372240 220728 372252
rect 220780 372240 220786 372292
rect 93578 372172 93584 372224
rect 93636 372212 93642 372224
rect 210970 372212 210976 372224
rect 93636 372184 210976 372212
rect 93636 372172 93642 372184
rect 210970 372172 210976 372184
rect 211028 372172 211034 372224
rect 214558 372212 214564 372224
rect 211172 372184 214564 372212
rect 211172 372076 211200 372184
rect 214558 372172 214564 372184
rect 214616 372212 214622 372224
rect 219710 372212 219716 372224
rect 214616 372184 219716 372212
rect 214616 372172 214622 372184
rect 219710 372172 219716 372184
rect 219768 372212 219774 372224
rect 220538 372212 220544 372224
rect 219768 372184 220544 372212
rect 219768 372172 219774 372184
rect 220538 372172 220544 372184
rect 220596 372172 220602 372224
rect 375190 372172 375196 372224
rect 375248 372212 375254 372224
rect 379514 372212 379520 372224
rect 375248 372184 379520 372212
rect 375248 372172 375254 372184
rect 379514 372172 379520 372184
rect 379572 372172 379578 372224
rect 211246 372104 211252 372156
rect 211304 372144 211310 372156
rect 221090 372144 221096 372156
rect 211304 372116 221096 372144
rect 211304 372104 211310 372116
rect 221090 372104 221096 372116
rect 221148 372144 221154 372156
rect 222102 372144 222108 372156
rect 221148 372116 222108 372144
rect 221148 372104 221154 372116
rect 222102 372104 222108 372116
rect 222160 372104 222166 372156
rect 371050 372104 371056 372156
rect 371108 372144 371114 372156
rect 377950 372144 377956 372156
rect 371108 372116 377956 372144
rect 371108 372104 371114 372116
rect 377950 372104 377956 372116
rect 378008 372104 378014 372156
rect 379974 372104 379980 372156
rect 380032 372144 380038 372156
rect 396074 372144 396080 372156
rect 380032 372116 396080 372144
rect 380032 372104 380038 372116
rect 396074 372104 396080 372116
rect 396132 372104 396138 372156
rect 219618 372076 219624 372088
rect 205606 372048 211200 372076
rect 219406 372048 219624 372076
rect 47394 371968 47400 372020
rect 47452 372008 47458 372020
rect 78490 372008 78496 372020
rect 47452 371980 78496 372008
rect 47452 371968 47458 371980
rect 78490 371968 78496 371980
rect 78548 371968 78554 372020
rect 92198 371968 92204 372020
rect 92256 372008 92262 372020
rect 205606 372008 205634 372048
rect 92256 371980 205634 372008
rect 92256 371968 92262 371980
rect 208210 371968 208216 372020
rect 208268 372008 208274 372020
rect 213638 372008 213644 372020
rect 208268 371980 213644 372008
rect 208268 371968 208274 371980
rect 213638 371968 213644 371980
rect 213696 371968 213702 372020
rect 46198 371900 46204 371952
rect 46256 371940 46262 371952
rect 79962 371940 79968 371952
rect 46256 371912 79968 371940
rect 46256 371900 46262 371912
rect 79962 371900 79968 371912
rect 80020 371900 80026 371952
rect 212350 371940 212356 371952
rect 200086 371912 212356 371940
rect 47486 371832 47492 371884
rect 47544 371872 47550 371884
rect 80146 371872 80152 371884
rect 47544 371844 80152 371872
rect 47544 371832 47550 371844
rect 80146 371832 80152 371844
rect 80204 371832 80210 371884
rect 85482 371764 85488 371816
rect 85540 371804 85546 371816
rect 105170 371804 105176 371816
rect 85540 371776 105176 371804
rect 85540 371764 85546 371776
rect 105170 371764 105176 371776
rect 105228 371764 105234 371816
rect 112898 371764 112904 371816
rect 112956 371804 112962 371816
rect 200086 371804 200114 371912
rect 212350 371900 212356 371912
rect 212408 371900 212414 371952
rect 208762 371832 208768 371884
rect 208820 371872 208826 371884
rect 209958 371872 209964 371884
rect 208820 371844 209964 371872
rect 208820 371832 208826 371844
rect 209958 371832 209964 371844
rect 210016 371872 210022 371884
rect 219406 371872 219434 372048
rect 219618 372036 219624 372048
rect 219676 372076 219682 372088
rect 241054 372076 241060 372088
rect 219676 372048 241060 372076
rect 219676 372036 219682 372048
rect 241054 372036 241060 372048
rect 241112 372036 241118 372088
rect 357158 372036 357164 372088
rect 357216 372076 357222 372088
rect 380986 372076 380992 372088
rect 357216 372048 380992 372076
rect 357216 372036 357222 372048
rect 380986 372036 380992 372048
rect 381044 372036 381050 372088
rect 220538 371968 220544 372020
rect 220596 372008 220602 372020
rect 251266 372008 251272 372020
rect 220596 371980 251272 372008
rect 220596 371968 220602 371980
rect 251266 371968 251272 371980
rect 251324 371968 251330 372020
rect 369854 371968 369860 372020
rect 369912 372008 369918 372020
rect 370406 372008 370412 372020
rect 369912 371980 370412 372008
rect 369912 371968 369918 371980
rect 370406 371968 370412 371980
rect 370464 372008 370470 372020
rect 397454 372008 397460 372020
rect 370464 371980 397460 372008
rect 370464 371968 370470 371980
rect 397454 371968 397460 371980
rect 397512 371968 397518 372020
rect 220906 371900 220912 371952
rect 220964 371940 220970 371952
rect 221826 371940 221832 371952
rect 220964 371912 221832 371940
rect 220964 371900 220970 371912
rect 221826 371900 221832 371912
rect 221884 371940 221890 371952
rect 252554 371940 252560 371952
rect 221884 371912 252560 371940
rect 221884 371900 221890 371912
rect 252554 371900 252560 371912
rect 252612 371900 252618 371952
rect 377858 371900 377864 371952
rect 377916 371940 377922 371952
rect 404354 371940 404360 371952
rect 377916 371912 404360 371940
rect 377916 371900 377922 371912
rect 404354 371900 404360 371912
rect 404412 371900 404418 371952
rect 210016 371844 219434 371872
rect 210016 371832 210022 371844
rect 224218 371832 224224 371884
rect 224276 371872 224282 371884
rect 247126 371872 247132 371884
rect 224276 371844 247132 371872
rect 224276 371832 224282 371844
rect 247126 371832 247132 371844
rect 247184 371832 247190 371884
rect 362770 371832 362776 371884
rect 362828 371872 362834 371884
rect 362828 371844 373994 371872
rect 362828 371832 362834 371844
rect 112956 371776 200114 371804
rect 112956 371764 112962 371776
rect 210050 371764 210056 371816
rect 210108 371804 210114 371816
rect 219526 371804 219532 371816
rect 210108 371776 219532 371804
rect 210108 371764 210114 371776
rect 219526 371764 219532 371776
rect 219584 371804 219590 371816
rect 248414 371804 248420 371816
rect 219584 371776 248420 371804
rect 219584 371764 219590 371776
rect 248414 371764 248420 371776
rect 248472 371764 248478 371816
rect 278682 371764 278688 371816
rect 278740 371804 278746 371816
rect 356606 371804 356612 371816
rect 278740 371776 356612 371804
rect 278740 371764 278746 371776
rect 356606 371764 356612 371776
rect 356664 371764 356670 371816
rect 373966 371804 373994 371844
rect 379330 371832 379336 371884
rect 379388 371872 379394 371884
rect 422294 371872 422300 371884
rect 379388 371844 422300 371872
rect 379388 371832 379394 371844
rect 422294 371832 422300 371844
rect 422352 371832 422358 371884
rect 518434 371832 518440 371884
rect 518492 371872 518498 371884
rect 580442 371872 580448 371884
rect 518492 371844 580448 371872
rect 518492 371832 518498 371844
rect 580442 371832 580448 371844
rect 580500 371832 580506 371884
rect 379146 371804 379152 371816
rect 373966 371776 379152 371804
rect 379146 371764 379152 371776
rect 379204 371804 379210 371816
rect 407114 371804 407120 371816
rect 379204 371776 407120 371804
rect 379204 371764 379210 371776
rect 407114 371764 407120 371776
rect 407172 371764 407178 371816
rect 208946 371736 208952 371748
rect 84166 371708 208952 371736
rect 46290 371424 46296 371476
rect 46348 371464 46354 371476
rect 49050 371464 49056 371476
rect 46348 371436 49056 371464
rect 46348 371424 46354 371436
rect 49050 371424 49056 371436
rect 49108 371464 49114 371476
rect 81986 371464 81992 371476
rect 49108 371436 81992 371464
rect 49108 371424 49114 371436
rect 81986 371424 81992 371436
rect 82044 371464 82050 371476
rect 84166 371464 84194 371708
rect 208946 371696 208952 371708
rect 209004 371696 209010 371748
rect 214374 371736 214380 371748
rect 210068 371708 214380 371736
rect 88058 371628 88064 371680
rect 88116 371668 88122 371680
rect 209866 371668 209872 371680
rect 88116 371640 209872 371668
rect 88116 371628 88122 371640
rect 209866 371628 209872 371640
rect 209924 371668 209930 371680
rect 210068 371668 210096 371708
rect 214374 371696 214380 371708
rect 214432 371696 214438 371748
rect 241698 371736 241704 371748
rect 219406 371708 241704 371736
rect 219406 371668 219434 371708
rect 241698 371696 241704 371708
rect 241756 371736 241762 371748
rect 242802 371736 242808 371748
rect 241756 371708 242808 371736
rect 241756 371696 241762 371708
rect 242802 371696 242808 371708
rect 242860 371696 242866 371748
rect 276014 371696 276020 371748
rect 276072 371736 276078 371748
rect 276934 371736 276940 371748
rect 276072 371708 276940 371736
rect 276072 371696 276078 371708
rect 276934 371696 276940 371708
rect 276992 371736 276998 371748
rect 356882 371736 356888 371748
rect 276992 371708 356888 371736
rect 276992 371696 276998 371708
rect 356882 371696 356888 371708
rect 356940 371696 356946 371748
rect 371234 371696 371240 371748
rect 371292 371736 371298 371748
rect 371602 371736 371608 371748
rect 371292 371708 371608 371736
rect 371292 371696 371298 371708
rect 371602 371696 371608 371708
rect 371660 371736 371666 371748
rect 401594 371736 401600 371748
rect 371660 371708 401600 371736
rect 371660 371696 371666 371708
rect 401594 371696 401600 371708
rect 401652 371696 401658 371748
rect 209924 371640 210096 371668
rect 210252 371640 219434 371668
rect 209924 371628 209930 371640
rect 82044 371436 84194 371464
rect 82044 371424 82050 371436
rect 90726 371424 90732 371476
rect 90784 371464 90790 371476
rect 208762 371464 208768 371476
rect 90784 371436 208768 371464
rect 90784 371424 90790 371436
rect 208762 371424 208768 371436
rect 208820 371424 208826 371476
rect 208946 371424 208952 371476
rect 209004 371464 209010 371476
rect 210252 371464 210280 371640
rect 222102 371628 222108 371680
rect 222160 371668 222166 371680
rect 251174 371668 251180 371680
rect 222160 371640 251180 371668
rect 222160 371628 222166 371640
rect 251174 371628 251180 371640
rect 251232 371628 251238 371680
rect 273346 371628 273352 371680
rect 273404 371668 273410 371680
rect 304994 371668 305000 371680
rect 273404 371640 305000 371668
rect 273404 371628 273410 371640
rect 304994 371628 305000 371640
rect 305052 371628 305058 371680
rect 368382 371628 368388 371680
rect 368440 371668 368446 371680
rect 378134 371668 378140 371680
rect 368440 371640 378140 371668
rect 368440 371628 368446 371640
rect 378134 371628 378140 371640
rect 378192 371628 378198 371680
rect 379514 371628 379520 371680
rect 379572 371668 379578 371680
rect 379698 371668 379704 371680
rect 379572 371640 379704 371668
rect 379572 371628 379578 371640
rect 379698 371628 379704 371640
rect 379756 371668 379762 371680
rect 409874 371668 409880 371680
rect 379756 371640 409880 371668
rect 379756 371628 379762 371640
rect 409874 371628 409880 371640
rect 409932 371628 409938 371680
rect 210970 371560 210976 371612
rect 211028 371600 211034 371612
rect 239306 371600 239312 371612
rect 211028 371572 239312 371600
rect 211028 371560 211034 371572
rect 239306 371560 239312 371572
rect 239364 371600 239370 371612
rect 367738 371600 367744 371612
rect 239364 371572 367744 371600
rect 239364 371560 239370 371572
rect 367738 371560 367744 371572
rect 367796 371600 367802 371612
rect 398834 371600 398840 371612
rect 367796 371572 398840 371600
rect 367796 371560 367802 371572
rect 398834 371560 398840 371572
rect 398892 371560 398898 371612
rect 240410 371532 240416 371544
rect 215266 371504 240416 371532
rect 212442 371464 212448 371476
rect 209004 371436 210280 371464
rect 210344 371436 212448 371464
rect 209004 371424 209010 371436
rect 79962 371356 79968 371408
rect 80020 371396 80026 371408
rect 210050 371396 210056 371408
rect 80020 371368 210056 371396
rect 80020 371356 80026 371368
rect 210050 371356 210056 371368
rect 210108 371356 210114 371408
rect 80146 371288 80152 371340
rect 80204 371328 80210 371340
rect 210344 371328 210372 371436
rect 212442 371424 212448 371436
rect 212500 371464 212506 371476
rect 215266 371464 215294 371504
rect 240410 371492 240416 371504
rect 240468 371532 240474 371544
rect 241422 371532 241428 371544
rect 240468 371504 241428 371532
rect 240468 371492 240474 371504
rect 241422 371492 241428 371504
rect 241480 371492 241486 371544
rect 242802 371492 242808 371544
rect 242860 371532 242866 371544
rect 371234 371532 371240 371544
rect 242860 371504 371240 371532
rect 242860 371492 242866 371504
rect 371234 371492 371240 371504
rect 371292 371492 371298 371544
rect 377950 371492 377956 371544
rect 378008 371532 378014 371544
rect 378008 371504 380572 371532
rect 378008 371492 378014 371504
rect 369854 371464 369860 371476
rect 212500 371436 215294 371464
rect 238726 371436 369860 371464
rect 212500 371424 212506 371436
rect 216398 371396 216404 371408
rect 80204 371300 210372 371328
rect 210436 371368 216404 371396
rect 80204 371288 80210 371300
rect 47394 371220 47400 371272
rect 47452 371260 47458 371272
rect 47578 371260 47584 371272
rect 47452 371232 47584 371260
rect 47452 371220 47458 371232
rect 47578 371220 47584 371232
rect 47636 371220 47642 371272
rect 78490 371220 78496 371272
rect 78548 371260 78554 371272
rect 210436 371260 210464 371368
rect 216398 371356 216404 371368
rect 216456 371396 216462 371408
rect 238110 371396 238116 371408
rect 216456 371368 238116 371396
rect 216456 371356 216462 371368
rect 238110 371356 238116 371368
rect 238168 371396 238174 371408
rect 238726 371396 238754 371436
rect 369854 371424 369860 371436
rect 369912 371424 369918 371476
rect 376570 371424 376576 371476
rect 376628 371464 376634 371476
rect 380544 371464 380572 371504
rect 380986 371492 380992 371544
rect 381044 371532 381050 371544
rect 411254 371532 411260 371544
rect 381044 371504 411260 371532
rect 381044 371492 381050 371504
rect 411254 371492 411260 371504
rect 411312 371492 411318 371544
rect 411346 371464 411352 371476
rect 376628 371436 380480 371464
rect 380544 371436 411352 371464
rect 376628 371424 376634 371436
rect 238168 371368 238754 371396
rect 238168 371356 238174 371368
rect 241422 371356 241428 371408
rect 241480 371396 241486 371408
rect 372890 371396 372896 371408
rect 241480 371368 372896 371396
rect 241480 371356 241486 371368
rect 372890 371356 372896 371368
rect 372948 371396 372954 371408
rect 373718 371396 373724 371408
rect 372948 371368 373724 371396
rect 372948 371356 372954 371368
rect 373718 371356 373724 371368
rect 373776 371356 373782 371408
rect 377030 371356 377036 371408
rect 377088 371396 377094 371408
rect 377858 371396 377864 371408
rect 377088 371368 377864 371396
rect 377088 371356 377094 371368
rect 377858 371356 377864 371368
rect 377916 371356 377922 371408
rect 380452 371396 380480 371436
rect 411346 371424 411352 371436
rect 411404 371424 411410 371476
rect 380986 371396 380992 371408
rect 380452 371368 380992 371396
rect 380986 371356 380992 371368
rect 381044 371396 381050 371408
rect 426434 371396 426440 371408
rect 381044 371368 426440 371396
rect 381044 371356 381050 371368
rect 426434 371356 426440 371368
rect 426492 371356 426498 371408
rect 213638 371288 213644 371340
rect 213696 371328 213702 371340
rect 245654 371328 245660 371340
rect 213696 371300 245660 371328
rect 213696 371288 213702 371300
rect 245654 371288 245660 371300
rect 245712 371288 245718 371340
rect 342254 371288 342260 371340
rect 342312 371328 342318 371340
rect 343358 371328 343364 371340
rect 342312 371300 343364 371328
rect 342312 371288 342318 371300
rect 343358 371288 343364 371300
rect 343416 371328 343422 371340
rect 360194 371328 360200 371340
rect 343416 371300 360200 371328
rect 343416 371288 343422 371300
rect 360194 371288 360200 371300
rect 360252 371328 360258 371340
rect 503530 371328 503536 371340
rect 360252 371300 503536 371328
rect 360252 371288 360258 371300
rect 503530 371288 503536 371300
rect 503588 371328 503594 371340
rect 517882 371328 517888 371340
rect 503588 371300 517888 371328
rect 503588 371288 503594 371300
rect 517882 371288 517888 371300
rect 517940 371328 517946 371340
rect 518434 371328 518440 371340
rect 517940 371300 518440 371328
rect 517940 371288 517946 371300
rect 518434 371288 518440 371300
rect 518492 371288 518498 371340
rect 78548 371232 210464 371260
rect 78548 371220 78554 371232
rect 220722 371220 220728 371272
rect 220780 371260 220786 371272
rect 220998 371260 221004 371272
rect 220780 371232 221004 371260
rect 220780 371220 220786 371232
rect 220998 371220 221004 371232
rect 221056 371260 221062 371272
rect 273254 371260 273260 371272
rect 221056 371232 273260 371260
rect 221056 371220 221062 371232
rect 273254 371220 273260 371232
rect 273312 371220 273318 371272
rect 342898 371220 342904 371272
rect 342956 371260 342962 371272
rect 357250 371260 357256 371272
rect 342956 371232 357256 371260
rect 342956 371220 342962 371232
rect 357250 371220 357256 371232
rect 357308 371260 357314 371272
rect 503162 371260 503168 371272
rect 357308 371232 503168 371260
rect 357308 371220 357314 371232
rect 503162 371220 503168 371232
rect 503220 371260 503226 371272
rect 517974 371260 517980 371272
rect 503220 371232 517980 371260
rect 503220 371220 503226 371232
rect 517974 371220 517980 371232
rect 518032 371260 518038 371272
rect 580258 371260 580264 371272
rect 518032 371232 580264 371260
rect 518032 371220 518038 371232
rect 580258 371220 580264 371232
rect 580316 371220 580322 371272
rect 40954 371152 40960 371204
rect 41012 371192 41018 371204
rect 182818 371192 182824 371204
rect 41012 371164 182824 371192
rect 41012 371152 41018 371164
rect 182818 371152 182824 371164
rect 182876 371152 182882 371204
rect 198734 371152 198740 371204
rect 198792 371192 198798 371204
rect 302234 371192 302240 371204
rect 198792 371164 302240 371192
rect 198792 371152 198798 371164
rect 302234 371152 302240 371164
rect 302292 371152 302298 371204
rect 356974 371152 356980 371204
rect 357032 371192 357038 371204
rect 477494 371192 477500 371204
rect 357032 371164 477500 371192
rect 357032 371152 357038 371164
rect 477494 371152 477500 371164
rect 477552 371152 477558 371204
rect 54478 371084 54484 371136
rect 54536 371124 54542 371136
rect 183462 371124 183468 371136
rect 54536 371096 183468 371124
rect 54536 371084 54542 371096
rect 183462 371084 183468 371096
rect 183520 371084 183526 371136
rect 198918 371084 198924 371136
rect 198976 371124 198982 371136
rect 300854 371124 300860 371136
rect 198976 371096 300860 371124
rect 198976 371084 198982 371096
rect 300854 371084 300860 371096
rect 300912 371084 300918 371136
rect 362126 371084 362132 371136
rect 362184 371124 362190 371136
rect 474734 371124 474740 371136
rect 362184 371096 474740 371124
rect 362184 371084 362190 371096
rect 474734 371084 474740 371096
rect 474792 371084 474798 371136
rect 102042 371016 102048 371068
rect 102100 371056 102106 371068
rect 213914 371056 213920 371068
rect 102100 371028 213920 371056
rect 102100 371016 102106 371028
rect 213914 371016 213920 371028
rect 213972 371016 213978 371068
rect 217410 371016 217416 371068
rect 217468 371056 217474 371068
rect 317414 371056 317420 371068
rect 217468 371028 317420 371056
rect 217468 371016 217474 371028
rect 317414 371016 317420 371028
rect 317472 371016 317478 371068
rect 364886 371016 364892 371068
rect 364944 371056 364950 371068
rect 473354 371056 473360 371068
rect 364944 371028 473360 371056
rect 364944 371016 364950 371028
rect 473354 371016 473360 371028
rect 473412 371016 473418 371068
rect 197538 370948 197544 371000
rect 197596 370988 197602 371000
rect 298094 370988 298100 371000
rect 197596 370960 298100 370988
rect 197596 370948 197602 370960
rect 298094 370948 298100 370960
rect 298152 370948 298158 371000
rect 360654 370948 360660 371000
rect 360712 370988 360718 371000
rect 465074 370988 465080 371000
rect 360712 370960 465080 370988
rect 360712 370948 360718 370960
rect 465074 370948 465080 370960
rect 465132 370948 465138 371000
rect 197446 370880 197452 370932
rect 197504 370920 197510 370932
rect 295334 370920 295340 370932
rect 197504 370892 295340 370920
rect 197504 370880 197510 370892
rect 295334 370880 295340 370892
rect 295392 370880 295398 370932
rect 367554 370880 367560 370932
rect 367612 370920 367618 370932
rect 470594 370920 470600 370932
rect 367612 370892 470600 370920
rect 367612 370880 367618 370892
rect 470594 370880 470600 370892
rect 470652 370880 470658 370932
rect 210050 370812 210056 370864
rect 210108 370852 210114 370864
rect 210970 370852 210976 370864
rect 210108 370824 210976 370852
rect 210108 370812 210114 370824
rect 210970 370812 210976 370824
rect 211028 370812 211034 370864
rect 212258 370812 212264 370864
rect 212316 370852 212322 370864
rect 307754 370852 307760 370864
rect 212316 370824 307760 370852
rect 212316 370812 212322 370824
rect 307754 370812 307760 370824
rect 307812 370812 307818 370864
rect 364794 370812 364800 370864
rect 364852 370852 364858 370864
rect 458174 370852 458180 370864
rect 364852 370824 458180 370852
rect 364852 370812 364858 370824
rect 458174 370812 458180 370824
rect 458232 370812 458238 370864
rect 198274 370744 198280 370796
rect 198332 370784 198338 370796
rect 292574 370784 292580 370796
rect 198332 370756 292580 370784
rect 198332 370744 198338 370756
rect 292574 370744 292580 370756
rect 292632 370744 292638 370796
rect 365622 370744 365628 370796
rect 365680 370784 365686 370796
rect 374546 370784 374552 370796
rect 365680 370756 374552 370784
rect 365680 370744 365686 370756
rect 374546 370744 374552 370756
rect 374604 370784 374610 370796
rect 375190 370784 375196 370796
rect 374604 370756 375196 370784
rect 374604 370744 374610 370756
rect 375190 370744 375196 370756
rect 375248 370744 375254 370796
rect 378134 370744 378140 370796
rect 378192 370784 378198 370796
rect 427814 370784 427820 370796
rect 378192 370756 427820 370784
rect 378192 370744 378198 370756
rect 427814 370744 427820 370756
rect 427872 370744 427878 370796
rect 196802 370676 196808 370728
rect 196860 370716 196866 370728
rect 289814 370716 289820 370728
rect 196860 370688 289820 370716
rect 196860 370676 196866 370688
rect 289814 370676 289820 370688
rect 289872 370676 289878 370728
rect 367002 370676 367008 370728
rect 367060 370716 367066 370728
rect 413186 370716 413192 370728
rect 367060 370688 413192 370716
rect 367060 370676 367066 370688
rect 413186 370676 413192 370688
rect 413244 370676 413250 370728
rect 196710 370608 196716 370660
rect 196768 370648 196774 370660
rect 287330 370648 287336 370660
rect 196768 370620 287336 370648
rect 196768 370608 196774 370620
rect 287330 370608 287336 370620
rect 287388 370608 287394 370660
rect 363506 370608 363512 370660
rect 363564 370648 363570 370660
rect 374914 370648 374920 370660
rect 363564 370620 374920 370648
rect 363564 370608 363570 370620
rect 374914 370608 374920 370620
rect 374972 370648 374978 370660
rect 375282 370648 375288 370660
rect 374972 370620 375288 370648
rect 374972 370608 374978 370620
rect 375282 370608 375288 370620
rect 375340 370608 375346 370660
rect 378042 370608 378048 370660
rect 378100 370648 378106 370660
rect 416774 370648 416780 370660
rect 378100 370620 416780 370648
rect 378100 370608 378106 370620
rect 416774 370608 416780 370620
rect 416832 370608 416838 370660
rect 196618 370540 196624 370592
rect 196676 370580 196682 370592
rect 285674 370580 285680 370592
rect 196676 370552 285680 370580
rect 196676 370540 196682 370552
rect 285674 370540 285680 370552
rect 285732 370540 285738 370592
rect 362678 370540 362684 370592
rect 362736 370580 362742 370592
rect 379882 370580 379888 370592
rect 362736 370552 379888 370580
rect 362736 370540 362742 370552
rect 379882 370540 379888 370552
rect 379940 370580 379946 370592
rect 414014 370580 414020 370592
rect 379940 370552 414020 370580
rect 379940 370540 379946 370552
rect 414014 370540 414020 370552
rect 414072 370540 414078 370592
rect 183462 370472 183468 370524
rect 183520 370512 183526 370524
rect 195974 370512 195980 370524
rect 183520 370484 195980 370512
rect 183520 370472 183526 370484
rect 195974 370472 195980 370484
rect 196032 370472 196038 370524
rect 196894 370472 196900 370524
rect 196952 370512 196958 370524
rect 282914 370512 282920 370524
rect 196952 370484 282920 370512
rect 196952 370472 196958 370484
rect 282914 370472 282920 370484
rect 282972 370472 282978 370524
rect 357066 370472 357072 370524
rect 357124 370512 357130 370524
rect 373074 370512 373080 370524
rect 357124 370484 373080 370512
rect 357124 370472 357130 370484
rect 373074 370472 373080 370484
rect 373132 370512 373138 370524
rect 373132 370484 373994 370512
rect 373132 370472 373138 370484
rect 196986 370404 196992 370456
rect 197044 370444 197050 370456
rect 277670 370444 277676 370456
rect 197044 370416 277676 370444
rect 197044 370404 197050 370416
rect 277670 370404 277676 370416
rect 277728 370404 277734 370456
rect 373966 370444 373994 370484
rect 375190 370472 375196 370524
rect 375248 370512 375254 370524
rect 415394 370512 415400 370524
rect 375248 370484 415400 370512
rect 375248 370472 375254 370484
rect 415394 370472 415400 370484
rect 415452 370472 415458 370524
rect 402974 370444 402980 370456
rect 373966 370416 402980 370444
rect 402974 370404 402980 370416
rect 403032 370404 403038 370456
rect 198826 370336 198832 370388
rect 198884 370376 198890 370388
rect 273346 370376 273352 370388
rect 198884 370348 273352 370376
rect 198884 370336 198890 370348
rect 273346 370336 273352 370348
rect 273404 370336 273410 370388
rect 375282 370336 375288 370388
rect 375340 370376 375346 370388
rect 396074 370376 396080 370388
rect 375340 370348 396080 370376
rect 375340 370336 375346 370348
rect 396074 370336 396080 370348
rect 396132 370336 396138 370388
rect 202874 369792 202880 369844
rect 202932 369832 202938 369844
rect 326154 369832 326160 369844
rect 202932 369804 326160 369832
rect 202932 369792 202938 369804
rect 326154 369792 326160 369804
rect 326212 369792 326218 369844
rect 363322 369792 363328 369844
rect 363380 369832 363386 369844
rect 480254 369832 480260 369844
rect 363380 369804 480260 369832
rect 363380 369792 363386 369804
rect 480254 369792 480260 369804
rect 480312 369792 480318 369844
rect 202506 369724 202512 369776
rect 202564 369764 202570 369776
rect 270494 369764 270500 369776
rect 202564 369736 270500 369764
rect 202564 369724 202570 369736
rect 270494 369724 270500 369736
rect 270552 369724 270558 369776
rect 369670 369724 369676 369776
rect 369728 369764 369734 369776
rect 483014 369764 483020 369776
rect 369728 369736 483020 369764
rect 369728 369724 369734 369736
rect 483014 369724 483020 369736
rect 483072 369724 483078 369776
rect 77018 369656 77024 369708
rect 77076 369696 77082 369708
rect 203150 369696 203156 369708
rect 77076 369668 203156 369696
rect 77076 369656 77082 369668
rect 203150 369656 203156 369668
rect 203208 369656 203214 369708
rect 206186 369656 206192 369708
rect 206244 369696 206250 369708
rect 280154 369696 280160 369708
rect 206244 369668 280160 369696
rect 206244 369656 206250 369668
rect 280154 369656 280160 369668
rect 280212 369656 280218 369708
rect 361298 369656 361304 369708
rect 361356 369696 361362 369708
rect 430574 369696 430580 369708
rect 361356 369668 430580 369696
rect 361356 369656 361362 369668
rect 430574 369656 430580 369668
rect 430632 369656 430638 369708
rect 211614 369588 211620 369640
rect 211672 369628 211678 369640
rect 276014 369628 276020 369640
rect 211672 369600 276020 369628
rect 211672 369588 211678 369600
rect 276014 369588 276020 369600
rect 276072 369588 276078 369640
rect 358446 369588 358452 369640
rect 358504 369628 358510 369640
rect 425054 369628 425060 369640
rect 358504 369600 425060 369628
rect 358504 369588 358510 369600
rect 425054 369588 425060 369600
rect 425112 369588 425118 369640
rect 208026 369520 208032 369572
rect 208084 369560 208090 369572
rect 264974 369560 264980 369572
rect 208084 369532 264980 369560
rect 208084 369520 208090 369532
rect 264974 369520 264980 369532
rect 265032 369520 265038 369572
rect 372430 369520 372436 369572
rect 372488 369560 372494 369572
rect 374362 369560 374368 369572
rect 372488 369532 374368 369560
rect 372488 369520 372494 369532
rect 374362 369520 374368 369532
rect 374420 369520 374426 369572
rect 378686 369520 378692 369572
rect 378744 369560 378750 369572
rect 430666 369560 430672 369572
rect 378744 369532 430672 369560
rect 378744 369520 378750 369532
rect 430666 369520 430672 369532
rect 430724 369520 430730 369572
rect 208854 369452 208860 369504
rect 208912 369492 208918 369504
rect 273438 369492 273444 369504
rect 208912 369464 273444 369492
rect 208912 369452 208918 369464
rect 273438 369452 273444 369464
rect 273496 369452 273502 369504
rect 373810 369452 373816 369504
rect 373868 369492 373874 369504
rect 429194 369492 429200 369504
rect 373868 369464 429200 369492
rect 373868 369452 373874 369464
rect 429194 369452 429200 369464
rect 429252 369452 429258 369504
rect 205358 369384 205364 369436
rect 205416 369424 205422 369436
rect 267734 369424 267740 369436
rect 205416 369396 267740 369424
rect 205416 369384 205422 369396
rect 267734 369384 267740 369396
rect 267792 369384 267798 369436
rect 370314 369384 370320 369436
rect 370372 369424 370378 369436
rect 420914 369424 420920 369436
rect 370372 369396 420920 369424
rect 370372 369384 370378 369396
rect 420914 369384 420920 369396
rect 420972 369384 420978 369436
rect 203794 369316 203800 369368
rect 203852 369356 203858 369368
rect 252554 369356 252560 369368
rect 203852 369328 252560 369356
rect 203852 369316 203858 369328
rect 252554 369316 252560 369328
rect 252612 369316 252618 369368
rect 358538 369316 358544 369368
rect 358596 369356 358602 369368
rect 376938 369356 376944 369368
rect 358596 369328 376944 369356
rect 358596 369316 358602 369328
rect 376938 369316 376944 369328
rect 376996 369356 377002 369368
rect 423674 369356 423680 369368
rect 376996 369328 423680 369356
rect 376996 369316 377002 369328
rect 423674 369316 423680 369328
rect 423732 369316 423738 369368
rect 99282 369248 99288 369300
rect 99340 369288 99346 369300
rect 212718 369288 212724 369300
rect 99340 369260 212724 369288
rect 99340 369248 99346 369260
rect 212718 369248 212724 369260
rect 212776 369248 212782 369300
rect 216306 369248 216312 369300
rect 216364 369288 216370 369300
rect 260834 369288 260840 369300
rect 216364 369260 260840 369288
rect 216364 369248 216370 369260
rect 260834 369248 260840 369260
rect 260892 369248 260898 369300
rect 373902 369248 373908 369300
rect 373960 369288 373966 369300
rect 375190 369288 375196 369300
rect 373960 369260 375196 369288
rect 373960 369248 373966 369260
rect 375190 369248 375196 369260
rect 375248 369288 375254 369300
rect 418154 369288 418160 369300
rect 375248 369260 418160 369288
rect 375248 369248 375254 369260
rect 418154 369248 418160 369260
rect 418212 369248 418218 369300
rect 106090 369180 106096 369232
rect 106148 369220 106154 369232
rect 217870 369220 217876 369232
rect 106148 369192 217876 369220
rect 106148 369180 106154 369192
rect 217870 369180 217876 369192
rect 217928 369180 217934 369232
rect 219158 369180 219164 369232
rect 219216 369220 219222 369232
rect 263594 369220 263600 369232
rect 219216 369192 263600 369220
rect 219216 369180 219222 369192
rect 263594 369180 263600 369192
rect 263652 369180 263658 369232
rect 366266 369180 366272 369232
rect 366324 369220 366330 369232
rect 375834 369220 375840 369232
rect 366324 369192 375840 369220
rect 366324 369180 366330 369192
rect 375834 369180 375840 369192
rect 375892 369220 375898 369232
rect 419534 369220 419540 369232
rect 375892 369192 419540 369220
rect 375892 369180 375898 369192
rect 419534 369180 419540 369192
rect 419592 369180 419598 369232
rect 100478 369112 100484 369164
rect 100536 369152 100542 369164
rect 212258 369152 212264 369164
rect 100536 369124 212264 369152
rect 100536 369112 100542 369124
rect 212258 369112 212264 369124
rect 212316 369152 212322 369164
rect 214006 369152 214012 369164
rect 212316 369124 214012 369152
rect 212316 369112 212322 369124
rect 214006 369112 214012 369124
rect 214064 369112 214070 369164
rect 214834 369112 214840 369164
rect 214892 369152 214898 369164
rect 258166 369152 258172 369164
rect 214892 369124 258172 369152
rect 214892 369112 214898 369124
rect 258166 369112 258172 369124
rect 258224 369112 258230 369164
rect 421006 369152 421012 369164
rect 373966 369124 421012 369152
rect 210326 369044 210332 369096
rect 210384 369084 210390 369096
rect 247034 369084 247040 369096
rect 210384 369056 247040 369084
rect 210384 369044 210390 369056
rect 247034 369044 247040 369056
rect 247092 369044 247098 369096
rect 367646 369044 367652 369096
rect 367704 369084 367710 369096
rect 371786 369084 371792 369096
rect 367704 369056 371792 369084
rect 367704 369044 367710 369056
rect 371786 369044 371792 369056
rect 371844 369084 371850 369096
rect 373966 369084 373994 369124
rect 421006 369112 421012 369124
rect 421064 369112 421070 369164
rect 371844 369056 373994 369084
rect 371844 369044 371850 369056
rect 374454 369044 374460 369096
rect 374512 369084 374518 369096
rect 375926 369084 375932 369096
rect 374512 369056 375932 369084
rect 374512 369044 374518 369056
rect 375926 369044 375932 369056
rect 375984 369084 375990 369096
rect 418246 369084 418252 369096
rect 375984 369056 418252 369084
rect 375984 369044 375990 369056
rect 418246 369044 418252 369056
rect 418304 369044 418310 369096
rect 97718 368976 97724 369028
rect 97776 369016 97782 369028
rect 210142 369016 210148 369028
rect 97776 368988 210148 369016
rect 97776 368976 97782 368988
rect 210142 368976 210148 368988
rect 210200 369016 210206 369028
rect 210878 369016 210884 369028
rect 210200 368988 210884 369016
rect 210200 368976 210206 368988
rect 210878 368976 210884 368988
rect 210936 368976 210942 369028
rect 370222 368976 370228 369028
rect 370280 369016 370286 369028
rect 371050 369016 371056 369028
rect 370280 368988 371056 369016
rect 370280 368976 370286 368988
rect 371050 368976 371056 368988
rect 371108 369016 371114 369028
rect 378686 369016 378692 369028
rect 371108 368988 378692 369016
rect 371108 368976 371114 368988
rect 378686 368976 378692 368988
rect 378744 368976 378750 369028
rect 105170 368908 105176 368960
rect 105228 368948 105234 368960
rect 210234 368948 210240 368960
rect 105228 368920 210240 368948
rect 105228 368908 105234 368920
rect 210234 368908 210240 368920
rect 210292 368948 210298 368960
rect 210786 368948 210792 368960
rect 210292 368920 210792 368948
rect 210292 368908 210298 368920
rect 210786 368908 210792 368920
rect 210844 368908 210850 368960
rect 101122 368840 101128 368892
rect 101180 368880 101186 368892
rect 213086 368880 213092 368892
rect 101180 368852 213092 368880
rect 101180 368840 101186 368852
rect 213086 368840 213092 368852
rect 213144 368840 213150 368892
rect 195974 368432 195980 368484
rect 196032 368472 196038 368484
rect 196710 368472 196716 368484
rect 196032 368444 196716 368472
rect 196032 368432 196038 368444
rect 196710 368432 196716 368444
rect 196768 368472 196774 368484
rect 342254 368472 342260 368484
rect 196768 368444 342260 368472
rect 196768 368432 196774 368444
rect 342254 368432 342260 368444
rect 342312 368432 342318 368484
rect 372522 368432 372528 368484
rect 372580 368472 372586 368484
rect 374454 368472 374460 368484
rect 372580 368444 374460 368472
rect 372580 368432 372586 368444
rect 374454 368432 374460 368444
rect 374512 368472 374518 368484
rect 375282 368472 375288 368484
rect 374512 368444 375288 368472
rect 374512 368432 374518 368444
rect 375282 368432 375288 368444
rect 375340 368432 375346 368484
rect 375742 368432 375748 368484
rect 375800 368472 375806 368484
rect 376570 368472 376576 368484
rect 375800 368444 376576 368472
rect 375800 368432 375806 368444
rect 376570 368432 376576 368444
rect 376628 368472 376634 368484
rect 436094 368472 436100 368484
rect 376628 368444 436100 368472
rect 376628 368432 376634 368444
rect 436094 368432 436100 368444
rect 436152 368432 436158 368484
rect 374362 368364 374368 368416
rect 374420 368404 374426 368416
rect 434714 368404 434720 368416
rect 374420 368376 434720 368404
rect 374420 368364 374426 368376
rect 434714 368364 434720 368376
rect 434772 368364 434778 368416
rect 361390 367888 361396 367940
rect 361448 367928 361454 367940
rect 379330 367928 379336 367940
rect 361448 367900 379336 367928
rect 361448 367888 361454 367900
rect 379330 367888 379336 367900
rect 379388 367928 379394 367940
rect 412634 367928 412640 367940
rect 379388 367900 412640 367928
rect 379388 367888 379394 367900
rect 412634 367888 412640 367900
rect 412692 367888 412698 367940
rect 375282 367820 375288 367872
rect 375340 367860 375346 367872
rect 431954 367860 431960 367872
rect 375340 367832 431960 367860
rect 375340 367820 375346 367832
rect 431954 367820 431960 367832
rect 432012 367820 432018 367872
rect 107562 367752 107568 367804
rect 107620 367792 107626 367804
rect 214834 367792 214840 367804
rect 107620 367764 214840 367792
rect 107620 367752 107626 367764
rect 214834 367752 214840 367764
rect 214892 367752 214898 367804
rect 369026 367752 369032 367804
rect 369084 367792 369090 367804
rect 373166 367792 373172 367804
rect 369084 367764 373172 367792
rect 369084 367752 369090 367764
rect 373166 367752 373172 367764
rect 373224 367792 373230 367804
rect 433334 367792 433340 367804
rect 373224 367764 433340 367792
rect 373224 367752 373230 367764
rect 433334 367752 433340 367764
rect 433392 367752 433398 367804
rect 374914 367548 374920 367600
rect 374972 367588 374978 367600
rect 375190 367588 375196 367600
rect 374972 367560 375196 367588
rect 374972 367548 374978 367560
rect 375190 367548 375196 367560
rect 375248 367548 375254 367600
rect 199378 365644 199384 365696
rect 199436 365684 199442 365696
rect 199562 365684 199568 365696
rect 199436 365656 199568 365684
rect 199436 365644 199442 365656
rect 199562 365644 199568 365656
rect 199620 365644 199626 365696
rect 199378 364964 199384 365016
rect 199436 365004 199442 365016
rect 359182 365004 359188 365016
rect 199436 364976 359188 365004
rect 199436 364964 199442 364976
rect 359182 364964 359188 364976
rect 359240 364964 359246 365016
rect 359734 364964 359740 365016
rect 359792 365004 359798 365016
rect 519170 365004 519176 365016
rect 359792 364976 519176 365004
rect 359792 364964 359798 364976
rect 519170 364964 519176 364976
rect 519228 365004 519234 365016
rect 519446 365004 519452 365016
rect 519228 364976 519452 365004
rect 519228 364964 519234 364976
rect 519446 364964 519452 364976
rect 519504 364964 519510 365016
rect 359826 363604 359832 363656
rect 359884 363644 359890 363656
rect 519170 363644 519176 363656
rect 359884 363616 519176 363644
rect 359884 363604 359890 363616
rect 519170 363604 519176 363616
rect 519228 363604 519234 363656
rect 199654 362176 199660 362228
rect 199712 362216 199718 362228
rect 200022 362216 200028 362228
rect 199712 362188 200028 362216
rect 199712 362176 199718 362188
rect 200022 362176 200028 362188
rect 200080 362216 200086 362228
rect 358998 362216 359004 362228
rect 200080 362188 359004 362216
rect 200080 362176 200086 362188
rect 358998 362176 359004 362188
rect 359056 362216 359062 362228
rect 359182 362216 359188 362228
rect 359056 362188 359188 362216
rect 359056 362176 359062 362188
rect 359182 362176 359188 362188
rect 359240 362216 359246 362228
rect 518986 362216 518992 362228
rect 359240 362188 518992 362216
rect 359240 362176 359246 362188
rect 518986 362176 518992 362188
rect 519044 362216 519050 362228
rect 519262 362216 519268 362228
rect 519044 362188 519268 362216
rect 519044 362176 519050 362188
rect 519262 362176 519268 362188
rect 519320 362176 519326 362228
rect 182818 360816 182824 360868
rect 182876 360856 182882 360868
rect 197446 360856 197452 360868
rect 182876 360828 197452 360856
rect 182876 360816 182882 360828
rect 197446 360816 197452 360828
rect 197504 360856 197510 360868
rect 342898 360856 342904 360868
rect 197504 360828 342904 360856
rect 197504 360816 197510 360828
rect 342898 360816 342904 360828
rect 342956 360816 342962 360868
rect 359458 359524 359464 359576
rect 359516 359564 359522 359576
rect 519078 359564 519084 359576
rect 359516 359536 519084 359564
rect 359516 359524 359522 359536
rect 519078 359524 519084 359536
rect 519136 359524 519142 359576
rect 199470 359456 199476 359508
rect 199528 359496 199534 359508
rect 358998 359496 359004 359508
rect 199528 359468 359004 359496
rect 199528 359456 199534 359468
rect 358998 359456 359004 359468
rect 359056 359496 359062 359508
rect 359734 359496 359740 359508
rect 359056 359468 359740 359496
rect 359056 359456 359062 359468
rect 359734 359456 359740 359468
rect 359792 359456 359798 359508
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 18598 358748 18604 358760
rect 3384 358720 18604 358748
rect 3384 358708 3390 358720
rect 18598 358708 18604 358720
rect 18656 358708 18662 358760
rect 359090 357348 359096 357400
rect 359148 357388 359154 357400
rect 359826 357388 359832 357400
rect 359148 357360 359832 357388
rect 359148 357348 359154 357360
rect 359826 357348 359832 357360
rect 359884 357348 359890 357400
rect 199562 356668 199568 356720
rect 199620 356708 199626 356720
rect 199838 356708 199844 356720
rect 199620 356680 199844 356708
rect 199620 356668 199626 356680
rect 199838 356668 199844 356680
rect 199896 356708 199902 356720
rect 359090 356708 359096 356720
rect 199896 356680 359096 356708
rect 199896 356668 199902 356680
rect 359090 356668 359096 356680
rect 359148 356668 359154 356720
rect 179138 355988 179144 356040
rect 179196 356028 179202 356040
rect 197262 356028 197268 356040
rect 179196 356000 197268 356028
rect 179196 355988 179202 356000
rect 197262 355988 197268 356000
rect 197320 355988 197326 356040
rect 357342 355988 357348 356040
rect 357400 356028 357406 356040
rect 358814 356028 358820 356040
rect 357400 356000 358820 356028
rect 357400 355988 357406 356000
rect 358814 355988 358820 356000
rect 358872 355988 358878 356040
rect 500862 355444 500868 355496
rect 500920 355484 500926 355496
rect 517606 355484 517612 355496
rect 500920 355456 517612 355484
rect 500920 355444 500926 355456
rect 517606 355444 517612 355456
rect 517664 355444 517670 355496
rect 338482 355376 338488 355428
rect 338540 355416 338546 355428
rect 357434 355416 357440 355428
rect 338540 355388 357440 355416
rect 338540 355376 338546 355388
rect 357434 355376 357440 355388
rect 357492 355376 357498 355428
rect 498838 355376 498844 355428
rect 498896 355416 498902 355428
rect 517698 355416 517704 355428
rect 498896 355388 517704 355416
rect 498896 355376 498902 355388
rect 517698 355376 517704 355388
rect 517756 355376 517762 355428
rect 191466 355308 191472 355360
rect 191524 355348 191530 355360
rect 191742 355348 191748 355360
rect 191524 355320 191748 355348
rect 191524 355308 191530 355320
rect 191742 355308 191748 355320
rect 191800 355348 191806 355360
rect 214558 355348 214564 355360
rect 191800 355320 214564 355348
rect 191800 355308 191806 355320
rect 214558 355308 214564 355320
rect 214616 355308 214622 355360
rect 351730 355308 351736 355360
rect 351788 355348 351794 355360
rect 375374 355348 375380 355360
rect 351788 355320 375380 355348
rect 351788 355308 351794 355320
rect 375374 355308 375380 355320
rect 375432 355308 375438 355360
rect 375374 355104 375380 355156
rect 375432 355144 375438 355156
rect 376018 355144 376024 355156
rect 375432 355116 376024 355144
rect 375432 355104 375438 355116
rect 376018 355104 376024 355116
rect 376076 355104 376082 355156
rect 179690 354696 179696 354748
rect 179748 354736 179754 354748
rect 197538 354736 197544 354748
rect 179748 354708 197544 354736
rect 179748 354696 179754 354708
rect 197538 354696 197544 354708
rect 197596 354736 197602 354748
rect 201586 354736 201592 354748
rect 197596 354708 201592 354736
rect 197596 354696 197602 354708
rect 201586 354696 201592 354708
rect 201644 354696 201650 354748
rect 339770 354696 339776 354748
rect 339828 354736 339834 354748
rect 357342 354736 357348 354748
rect 339828 354708 357348 354736
rect 339828 354696 339834 354708
rect 357342 354696 357348 354708
rect 357400 354696 357406 354748
rect 510890 354696 510896 354748
rect 510948 354736 510954 354748
rect 517514 354736 517520 354748
rect 510948 354708 517520 354736
rect 510948 354696 510954 354708
rect 517514 354696 517520 354708
rect 517572 354696 517578 354748
rect 371694 353948 371700 354000
rect 371752 353988 371758 354000
rect 380894 353988 380900 354000
rect 371752 353960 380900 353988
rect 371752 353948 371758 353960
rect 380894 353948 380900 353960
rect 380952 353948 380958 354000
rect 218422 353404 218428 353456
rect 218480 353444 218486 353456
rect 221090 353444 221096 353456
rect 218480 353416 221096 353444
rect 218480 353404 218486 353416
rect 221090 353404 221096 353416
rect 221148 353404 221154 353456
rect 56042 353336 56048 353388
rect 56100 353376 56106 353388
rect 59814 353376 59820 353388
rect 56100 353348 59820 353376
rect 56100 353336 56106 353348
rect 59814 353336 59820 353348
rect 59872 353336 59878 353388
rect 218606 353336 218612 353388
rect 218664 353376 218670 353388
rect 220906 353376 220912 353388
rect 218664 353348 220912 353376
rect 218664 353336 218670 353348
rect 220906 353336 220912 353348
rect 220964 353336 220970 353388
rect 378686 353336 378692 353388
rect 378744 353376 378750 353388
rect 381078 353376 381084 353388
rect 378744 353348 381084 353376
rect 378744 353336 378750 353348
rect 381078 353336 381084 353348
rect 381136 353336 381142 353388
rect 58526 353268 58532 353320
rect 58584 353308 58590 353320
rect 60734 353308 60740 353320
rect 58584 353280 60740 353308
rect 58584 353268 58590 353280
rect 60734 353268 60740 353280
rect 60792 353268 60798 353320
rect 218514 353268 218520 353320
rect 218572 353308 218578 353320
rect 220814 353308 220820 353320
rect 218572 353280 220820 353308
rect 218572 353268 218578 353280
rect 220814 353268 220820 353280
rect 220872 353268 220878 353320
rect 378594 353268 378600 353320
rect 378652 353308 378658 353320
rect 380986 353308 380992 353320
rect 378652 353280 380992 353308
rect 378652 353268 378658 353280
rect 380986 353268 380992 353280
rect 381044 353268 381050 353320
rect 57054 351976 57060 352028
rect 57112 352016 57118 352028
rect 59354 352016 59360 352028
rect 57112 351988 59360 352016
rect 57112 351976 57118 351988
rect 59354 351976 59360 351988
rect 59412 351976 59418 352028
rect 55950 351908 55956 351960
rect 56008 351948 56014 351960
rect 57974 351948 57980 351960
rect 56008 351920 57980 351948
rect 56008 351908 56014 351920
rect 57974 351908 57980 351920
rect 58032 351908 58038 351960
rect 54478 303764 54484 303816
rect 54536 303804 54542 303816
rect 56594 303804 56600 303816
rect 54536 303776 56600 303804
rect 54536 303764 54542 303776
rect 56594 303764 56600 303776
rect 56652 303764 56658 303816
rect 46382 299412 46388 299464
rect 46440 299452 46446 299464
rect 56962 299452 56968 299464
rect 46440 299424 56968 299452
rect 46440 299412 46446 299424
rect 56962 299412 56968 299424
rect 57020 299452 57026 299464
rect 57422 299452 57428 299464
rect 57020 299424 57428 299452
rect 57020 299412 57026 299424
rect 57422 299412 57428 299424
rect 57480 299412 57486 299464
rect 46474 298052 46480 298104
rect 46532 298092 46538 298104
rect 57422 298092 57428 298104
rect 46532 298064 57428 298092
rect 46532 298052 46538 298064
rect 57422 298052 57428 298064
rect 57480 298052 57486 298104
rect 519906 284316 519912 284368
rect 519964 284356 519970 284368
rect 580258 284356 580264 284368
rect 519964 284328 580264 284356
rect 519964 284316 519970 284328
rect 580258 284316 580264 284328
rect 580316 284316 580322 284368
rect 519170 282888 519176 282940
rect 519228 282928 519234 282940
rect 580350 282928 580356 282940
rect 519228 282900 580356 282928
rect 519228 282888 519234 282900
rect 580350 282888 580356 282900
rect 580408 282888 580414 282940
rect 377766 282208 377772 282260
rect 377824 282248 377830 282260
rect 377950 282248 377956 282260
rect 377824 282220 377956 282248
rect 377824 282208 377830 282220
rect 377950 282208 377956 282220
rect 378008 282208 378014 282260
rect 200942 280100 200948 280152
rect 201000 280140 201006 280152
rect 216674 280140 216680 280152
rect 201000 280112 216680 280140
rect 201000 280100 201006 280112
rect 216674 280100 216680 280112
rect 216732 280100 216738 280152
rect 368290 280100 368296 280152
rect 368348 280140 368354 280152
rect 377030 280140 377036 280152
rect 368348 280112 377036 280140
rect 368348 280100 368354 280112
rect 377030 280100 377036 280112
rect 377088 280100 377094 280152
rect 205266 278672 205272 278724
rect 205324 278712 205330 278724
rect 216858 278712 216864 278724
rect 205324 278684 216864 278712
rect 205324 278672 205330 278684
rect 216858 278672 216864 278684
rect 216916 278672 216922 278724
rect 366910 278672 366916 278724
rect 366968 278712 366974 278724
rect 377030 278712 377036 278724
rect 366968 278684 377036 278712
rect 366968 278672 366974 278684
rect 377030 278672 377036 278684
rect 377088 278672 377094 278724
rect 214558 278264 214564 278316
rect 214616 278304 214622 278316
rect 216674 278304 216680 278316
rect 214616 278276 216680 278304
rect 214616 278264 214622 278276
rect 216674 278264 216680 278276
rect 216732 278264 216738 278316
rect 376018 278264 376024 278316
rect 376076 278304 376082 278316
rect 377398 278304 377404 278316
rect 376076 278276 377404 278304
rect 376076 278264 376082 278276
rect 377398 278264 377404 278276
rect 377456 278264 377462 278316
rect 214558 276564 214564 276616
rect 214616 276604 214622 276616
rect 215294 276604 215300 276616
rect 214616 276576 215300 276604
rect 214616 276564 214622 276576
rect 215294 276564 215300 276576
rect 215352 276564 215358 276616
rect 377766 274116 377772 274168
rect 377824 274156 377830 274168
rect 377950 274156 377956 274168
rect 377824 274128 377956 274156
rect 377824 274116 377830 274128
rect 377950 274116 377956 274128
rect 378008 274116 378014 274168
rect 213086 272552 213092 272604
rect 213144 272592 213150 272604
rect 213638 272592 213644 272604
rect 213144 272564 213644 272592
rect 213144 272552 213150 272564
rect 213638 272552 213644 272564
rect 213696 272552 213702 272604
rect 211706 270444 211712 270496
rect 211764 270484 211770 270496
rect 212902 270484 212908 270496
rect 211764 270456 212908 270484
rect 211764 270444 211770 270456
rect 212902 270444 212908 270456
rect 212960 270444 212966 270496
rect 378594 270444 378600 270496
rect 378652 270484 378658 270496
rect 379514 270484 379520 270496
rect 378652 270456 379520 270484
rect 378652 270444 378658 270456
rect 379514 270444 379520 270456
rect 379572 270444 379578 270496
rect 219250 270036 219256 270088
rect 219308 270076 219314 270088
rect 219802 270076 219808 270088
rect 219308 270048 219808 270076
rect 219308 270036 219314 270048
rect 219802 270036 219808 270048
rect 219860 270036 219866 270088
rect 60826 269628 60832 269680
rect 60884 269668 60890 269680
rect 107562 269668 107568 269680
rect 60884 269640 107568 269668
rect 60884 269628 60890 269640
rect 107562 269628 107568 269640
rect 107620 269628 107626 269680
rect 55858 269560 55864 269612
rect 55916 269600 55922 269612
rect 110966 269600 110972 269612
rect 55916 269572 110972 269600
rect 55916 269560 55922 269572
rect 110966 269560 110972 269572
rect 111024 269560 111030 269612
rect 219802 269560 219808 269612
rect 219860 269600 219866 269612
rect 263502 269600 263508 269612
rect 219860 269572 263508 269600
rect 219860 269560 219866 269572
rect 263502 269560 263508 269572
rect 263560 269560 263566 269612
rect 52914 269492 52920 269544
rect 52972 269532 52978 269544
rect 108298 269532 108304 269544
rect 52972 269504 108304 269532
rect 52972 269492 52978 269504
rect 108298 269492 108304 269504
rect 108356 269492 108362 269544
rect 200850 269492 200856 269544
rect 200908 269532 200914 269544
rect 250714 269532 250720 269544
rect 200908 269504 250720 269532
rect 200908 269492 200914 269504
rect 250714 269492 250720 269504
rect 250772 269492 250778 269544
rect 43346 269424 43352 269476
rect 43404 269464 43410 269476
rect 133414 269464 133420 269476
rect 43404 269436 133420 269464
rect 43404 269424 43410 269436
rect 133414 269424 133420 269436
rect 133472 269424 133478 269476
rect 218514 269424 218520 269476
rect 218572 269464 218578 269476
rect 279142 269464 279148 269476
rect 218572 269436 279148 269464
rect 218572 269424 218578 269436
rect 279142 269424 279148 269436
rect 279200 269424 279206 269476
rect 379238 269424 379244 269476
rect 379296 269464 379302 269476
rect 425238 269464 425244 269476
rect 379296 269436 425244 269464
rect 379296 269424 379302 269436
rect 425238 269424 425244 269436
rect 425296 269424 425302 269476
rect 45370 269356 45376 269408
rect 45428 269396 45434 269408
rect 135898 269396 135904 269408
rect 45428 269368 135904 269396
rect 45428 269356 45434 269368
rect 135898 269356 135904 269368
rect 135956 269356 135962 269408
rect 212902 269356 212908 269408
rect 212960 269396 212966 269408
rect 275738 269396 275744 269408
rect 212960 269368 275744 269396
rect 212960 269356 212966 269368
rect 275738 269356 275744 269368
rect 275796 269356 275802 269408
rect 379514 269356 379520 269408
rect 379572 269396 379578 269408
rect 426434 269396 426440 269408
rect 379572 269368 426440 269396
rect 379572 269356 379578 269368
rect 426434 269356 426440 269368
rect 426492 269356 426498 269408
rect 44818 269288 44824 269340
rect 44876 269328 44882 269340
rect 138474 269328 138480 269340
rect 44876 269300 138480 269328
rect 44876 269288 44882 269300
rect 138474 269288 138480 269300
rect 138532 269288 138538 269340
rect 214742 269288 214748 269340
rect 214800 269328 214806 269340
rect 280890 269328 280896 269340
rect 214800 269300 280896 269328
rect 214800 269288 214806 269300
rect 280890 269288 280896 269300
rect 280948 269288 280954 269340
rect 364150 269288 364156 269340
rect 364208 269328 364214 269340
rect 418430 269328 418436 269340
rect 364208 269300 418436 269328
rect 364208 269288 364214 269300
rect 418430 269288 418436 269300
rect 418488 269288 418494 269340
rect 45002 269220 45008 269272
rect 45060 269260 45066 269272
rect 140866 269260 140872 269272
rect 45060 269232 140872 269260
rect 45060 269220 45066 269232
rect 140866 269220 140872 269232
rect 140924 269220 140930 269272
rect 210694 269220 210700 269272
rect 210752 269260 210758 269272
rect 283466 269260 283472 269272
rect 210752 269232 283472 269260
rect 210752 269220 210758 269232
rect 283466 269220 283472 269232
rect 283524 269220 283530 269272
rect 373626 269220 373632 269272
rect 373684 269260 373690 269272
rect 433610 269260 433616 269272
rect 373684 269232 433616 269260
rect 373684 269220 373690 269232
rect 433610 269220 433616 269232
rect 433668 269220 433674 269272
rect 45094 269152 45100 269204
rect 45152 269192 45158 269204
rect 143534 269192 143540 269204
rect 45152 269164 143540 269192
rect 45152 269152 45158 269164
rect 143534 269152 143540 269164
rect 143592 269152 143598 269204
rect 212166 269152 212172 269204
rect 212224 269192 212230 269204
rect 288250 269192 288256 269204
rect 212224 269164 288256 269192
rect 212224 269152 212230 269164
rect 288250 269152 288256 269164
rect 288308 269152 288314 269204
rect 370958 269152 370964 269204
rect 371016 269192 371022 269204
rect 453390 269192 453396 269204
rect 371016 269164 453396 269192
rect 371016 269152 371022 269164
rect 453390 269152 453396 269164
rect 453448 269152 453454 269204
rect 44910 269084 44916 269136
rect 44968 269124 44974 269136
rect 145926 269124 145932 269136
rect 44968 269096 145932 269124
rect 44968 269084 44974 269096
rect 145926 269084 145932 269096
rect 145984 269084 145990 269136
rect 209314 269084 209320 269136
rect 209372 269124 209378 269136
rect 285950 269124 285956 269136
rect 209372 269096 285956 269124
rect 209372 269084 209378 269096
rect 285950 269084 285956 269096
rect 286008 269084 286014 269136
rect 368198 269084 368204 269136
rect 368256 269124 368262 269136
rect 468478 269124 468484 269136
rect 368256 269096 468484 269124
rect 368256 269084 368262 269096
rect 468478 269084 468484 269096
rect 468536 269084 468542 269136
rect 42518 269016 42524 269068
rect 42576 269056 42582 269068
rect 42576 269028 45554 269056
rect 42576 269016 42582 269028
rect 45526 268988 45554 269028
rect 59630 269016 59636 269068
rect 59688 269056 59694 269068
rect 60734 269056 60740 269068
rect 59688 269028 60740 269056
rect 59688 269016 59694 269028
rect 60734 269016 60740 269028
rect 60792 269016 60798 269068
rect 196618 269016 196624 269068
rect 196676 269056 196682 269068
rect 197630 269056 197636 269068
rect 196676 269028 197636 269056
rect 196676 269016 196682 269028
rect 197630 269016 197636 269028
rect 197688 269016 197694 269068
rect 213638 269016 213644 269068
rect 213696 269056 213702 269068
rect 214282 269056 214288 269068
rect 213696 269028 214288 269056
rect 213696 269016 213702 269028
rect 214282 269016 214288 269028
rect 214340 269016 214346 269068
rect 217134 269016 217140 269068
rect 217192 269056 217198 269068
rect 217778 269056 217784 269068
rect 217192 269028 217784 269056
rect 217192 269016 217198 269028
rect 217778 269016 217784 269028
rect 217836 269016 217842 269068
rect 374454 269016 374460 269068
rect 374512 269056 374518 269068
rect 374914 269056 374920 269068
rect 374512 269028 374920 269056
rect 374512 269016 374518 269028
rect 374914 269016 374920 269028
rect 374972 269016 374978 269068
rect 60826 268988 60832 269000
rect 45526 268960 60832 268988
rect 60826 268948 60832 268960
rect 60884 268948 60890 269000
rect 374546 268880 374552 268932
rect 374604 268920 374610 268932
rect 396074 268920 396080 268932
rect 374604 268892 396080 268920
rect 374604 268880 374610 268892
rect 396074 268880 396080 268892
rect 396132 268880 396138 268932
rect 206554 268812 206560 268864
rect 206612 268852 206618 268864
rect 290918 268852 290924 268864
rect 206612 268824 290924 268852
rect 206612 268812 206618 268824
rect 290918 268812 290924 268824
rect 290976 268812 290982 268864
rect 369118 268812 369124 268864
rect 369176 268852 369182 268864
rect 423490 268852 423496 268864
rect 369176 268824 423496 268852
rect 369176 268812 369182 268824
rect 423490 268812 423496 268824
rect 423548 268812 423554 268864
rect 49234 268744 49240 268796
rect 49292 268784 49298 268796
rect 83090 268784 83096 268796
rect 49292 268756 83096 268784
rect 49292 268744 49298 268756
rect 83090 268744 83096 268756
rect 83148 268744 83154 268796
rect 207934 268744 207940 268796
rect 207992 268784 207998 268796
rect 295886 268784 295892 268796
rect 207992 268756 295892 268784
rect 207992 268744 207998 268756
rect 295886 268744 295892 268756
rect 295944 268744 295950 268796
rect 366818 268744 366824 268796
rect 366876 268784 366882 268796
rect 421006 268784 421012 268796
rect 366876 268756 421012 268784
rect 366876 268744 366882 268756
rect 421006 268744 421012 268756
rect 421064 268744 421070 268796
rect 42610 268676 42616 268728
rect 42668 268716 42674 268728
rect 57790 268716 57796 268728
rect 42668 268688 57796 268716
rect 42668 268676 42674 268688
rect 57790 268676 57796 268688
rect 57848 268676 57854 268728
rect 203610 268676 203616 268728
rect 203668 268716 203674 268728
rect 293402 268716 293408 268728
rect 203668 268688 293408 268716
rect 203668 268676 203674 268688
rect 293402 268676 293408 268688
rect 293460 268676 293466 268728
rect 376386 268676 376392 268728
rect 376444 268716 376450 268728
rect 430942 268716 430948 268728
rect 376444 268688 430948 268716
rect 376444 268676 376450 268688
rect 430942 268676 430948 268688
rect 431000 268676 431006 268728
rect 47762 268608 47768 268660
rect 47820 268648 47826 268660
rect 77110 268648 77116 268660
rect 47820 268620 77116 268648
rect 47820 268608 47826 268620
rect 77110 268608 77116 268620
rect 77168 268608 77174 268660
rect 216214 268608 216220 268660
rect 216272 268648 216278 268660
rect 308490 268648 308496 268660
rect 216272 268620 308496 268648
rect 216272 268608 216278 268620
rect 308490 268608 308496 268620
rect 308548 268608 308554 268660
rect 375098 268608 375104 268660
rect 375156 268648 375162 268660
rect 478414 268648 478420 268660
rect 375156 268620 478420 268648
rect 375156 268608 375162 268620
rect 478414 268608 478420 268620
rect 478472 268608 478478 268660
rect 45186 268540 45192 268592
rect 45244 268580 45250 268592
rect 47394 268580 47400 268592
rect 45244 268552 47400 268580
rect 45244 268540 45250 268552
rect 47394 268540 47400 268552
rect 47452 268540 47458 268592
rect 47946 268540 47952 268592
rect 48004 268580 48010 268592
rect 90726 268580 90732 268592
rect 48004 268552 90732 268580
rect 48004 268540 48010 268552
rect 90726 268540 90732 268552
rect 90784 268540 90790 268592
rect 202414 268540 202420 268592
rect 202472 268580 202478 268592
rect 298462 268580 298468 268592
rect 202472 268552 298468 268580
rect 202472 268540 202478 268552
rect 298462 268540 298468 268552
rect 298520 268540 298526 268592
rect 372338 268540 372344 268592
rect 372396 268580 372402 268592
rect 475838 268580 475844 268592
rect 372396 268552 475844 268580
rect 372396 268540 372402 268552
rect 475838 268540 475844 268552
rect 475896 268540 475902 268592
rect 48038 268472 48044 268524
rect 48096 268512 48102 268524
rect 93578 268512 93584 268524
rect 48096 268484 93584 268512
rect 48096 268472 48102 268484
rect 93578 268472 93584 268484
rect 93636 268472 93642 268524
rect 205174 268472 205180 268524
rect 205232 268512 205238 268524
rect 300854 268512 300860 268524
rect 205232 268484 300860 268512
rect 205232 268472 205238 268484
rect 300854 268472 300860 268484
rect 300912 268472 300918 268524
rect 362586 268472 362592 268524
rect 362644 268512 362650 268524
rect 473354 268512 473360 268524
rect 362644 268484 473360 268512
rect 362644 268472 362650 268484
rect 473354 268472 473360 268484
rect 473412 268472 473418 268524
rect 43438 268404 43444 268456
rect 43496 268444 43502 268456
rect 47302 268444 47308 268456
rect 43496 268416 47308 268444
rect 43496 268404 43502 268416
rect 47302 268404 47308 268416
rect 47360 268404 47366 268456
rect 49142 268404 49148 268456
rect 49200 268444 49206 268456
rect 96062 268444 96068 268456
rect 49200 268416 96068 268444
rect 49200 268404 49206 268416
rect 96062 268404 96068 268416
rect 96120 268404 96126 268456
rect 213454 268404 213460 268456
rect 213512 268444 213518 268456
rect 318426 268444 318432 268456
rect 213512 268416 318432 268444
rect 213512 268404 213518 268416
rect 318426 268404 318432 268416
rect 318484 268404 318490 268456
rect 365530 268404 365536 268456
rect 365588 268444 365594 268456
rect 480898 268444 480904 268456
rect 365588 268416 480904 268444
rect 365588 268404 365594 268416
rect 480898 268404 480904 268416
rect 480956 268404 480962 268456
rect 51810 268336 51816 268388
rect 51868 268376 51874 268388
rect 98454 268376 98460 268388
rect 51868 268348 98460 268376
rect 51868 268336 51874 268348
rect 98454 268336 98460 268348
rect 98512 268336 98518 268388
rect 197998 268336 198004 268388
rect 198056 268376 198062 268388
rect 315850 268376 315856 268388
rect 198056 268348 315856 268376
rect 198056 268336 198062 268348
rect 315850 268336 315856 268348
rect 315908 268336 315914 268388
rect 361022 268336 361028 268388
rect 361080 268376 361086 268388
rect 483382 268376 483388 268388
rect 361080 268348 483388 268376
rect 361080 268336 361086 268348
rect 483382 268336 483388 268348
rect 483440 268336 483446 268388
rect 46658 268268 46664 268320
rect 46716 268308 46722 268320
rect 76006 268308 76012 268320
rect 46716 268280 76012 268308
rect 46716 268268 46722 268280
rect 76006 268268 76012 268280
rect 76064 268268 76070 268320
rect 47210 268200 47216 268252
rect 47268 268240 47274 268252
rect 47762 268240 47768 268252
rect 47268 268212 47768 268240
rect 47268 268200 47274 268212
rect 47762 268200 47768 268212
rect 47820 268200 47826 268252
rect 64874 268200 64880 268252
rect 64932 268240 64938 268252
rect 95878 268240 95884 268252
rect 64932 268212 95884 268240
rect 64932 268200 64938 268212
rect 95878 268200 95884 268212
rect 95936 268200 95942 268252
rect 62114 268132 62120 268184
rect 62172 268172 62178 268184
rect 94498 268172 94504 268184
rect 62172 268144 94504 268172
rect 62172 268132 62178 268144
rect 94498 268132 94504 268144
rect 94556 268132 94562 268184
rect 53834 268064 53840 268116
rect 53892 268104 53898 268116
rect 86954 268104 86960 268116
rect 53892 268076 86960 268104
rect 53892 268064 53898 268076
rect 86954 268064 86960 268076
rect 87012 268064 87018 268116
rect 373166 268064 373172 268116
rect 373224 268104 373230 268116
rect 374270 268104 374276 268116
rect 373224 268076 374276 268104
rect 373224 268064 373230 268076
rect 374270 268064 374276 268076
rect 374328 268104 374334 268116
rect 433334 268104 433340 268116
rect 374328 268076 433340 268104
rect 374328 268064 374334 268076
rect 433334 268064 433340 268076
rect 433392 268064 433398 268116
rect 58618 267996 58624 268048
rect 58676 268036 58682 268048
rect 58676 268008 64874 268036
rect 58676 267996 58682 268008
rect 64846 267968 64874 268008
rect 82078 267996 82084 268048
rect 82136 268036 82142 268048
rect 108666 268036 108672 268048
rect 82136 268008 108672 268036
rect 82136 267996 82142 268008
rect 108666 267996 108672 268008
rect 108724 267996 108730 268048
rect 396074 267996 396080 268048
rect 396132 268036 396138 268048
rect 415854 268036 415860 268048
rect 396132 268008 415860 268036
rect 396132 267996 396138 268008
rect 415854 267996 415860 268008
rect 415912 267996 415918 268048
rect 99374 267968 99380 267980
rect 64846 267940 99380 267968
rect 99374 267928 99380 267940
rect 99432 267928 99438 267980
rect 236638 267928 236644 267980
rect 236696 267968 236702 267980
rect 255774 267968 255780 267980
rect 236696 267940 255780 267968
rect 236696 267928 236702 267940
rect 255774 267928 255780 267940
rect 255832 267928 255838 267980
rect 356514 267928 356520 267980
rect 356572 267968 356578 267980
rect 360194 267968 360200 267980
rect 356572 267940 360200 267968
rect 356572 267928 356578 267940
rect 360194 267928 360200 267940
rect 360252 267928 360258 267980
rect 373074 267928 373080 267980
rect 373132 267968 373138 267980
rect 375650 267968 375656 267980
rect 373132 267940 375656 267968
rect 373132 267928 373138 267940
rect 375650 267928 375656 267940
rect 375708 267968 375714 267980
rect 402974 267968 402980 267980
rect 375708 267940 402980 267968
rect 375708 267928 375714 267940
rect 402974 267928 402980 267940
rect 403032 267928 403038 267980
rect 57790 267860 57796 267912
rect 57848 267900 57854 267912
rect 105262 267900 105268 267912
rect 57848 267872 105268 267900
rect 57848 267860 57854 267872
rect 105262 267860 105268 267872
rect 105320 267860 105326 267912
rect 214282 267860 214288 267912
rect 214340 267900 214346 267912
rect 243078 267900 243084 267912
rect 214340 267872 243084 267900
rect 214340 267860 214346 267872
rect 243078 267860 243084 267872
rect 243136 267860 243142 267912
rect 379882 267860 379888 267912
rect 379940 267900 379946 267912
rect 414382 267900 414388 267912
rect 379940 267872 414388 267900
rect 379940 267860 379946 267872
rect 414382 267860 414388 267872
rect 414440 267860 414446 267912
rect 421558 267860 421564 267912
rect 421616 267900 421622 267912
rect 435726 267900 435732 267912
rect 421616 267872 435732 267900
rect 421616 267860 421622 267872
rect 435726 267860 435732 267872
rect 435784 267860 435790 267912
rect 59722 267792 59728 267844
rect 59780 267832 59786 267844
rect 106366 267832 106372 267844
rect 59780 267804 106372 267832
rect 59780 267792 59786 267804
rect 106366 267792 106372 267804
rect 106424 267792 106430 267844
rect 217778 267792 217784 267844
rect 217836 267832 217842 267844
rect 258074 267832 258080 267844
rect 217836 267804 258080 267832
rect 217836 267792 217842 267804
rect 258074 267792 258080 267804
rect 258132 267792 258138 267844
rect 374914 267792 374920 267844
rect 374972 267832 374978 267844
rect 432138 267832 432144 267844
rect 374972 267804 432144 267832
rect 374972 267792 374978 267804
rect 432138 267792 432144 267804
rect 432196 267792 432202 267844
rect 54478 267724 54484 267776
rect 54536 267764 54542 267776
rect 102686 267764 102692 267776
rect 54536 267736 102692 267764
rect 54536 267724 54542 267736
rect 102686 267724 102692 267736
rect 102744 267724 102750 267776
rect 117130 267724 117136 267776
rect 117188 267764 117194 267776
rect 196618 267764 196624 267776
rect 117188 267736 196624 267764
rect 117188 267724 117194 267736
rect 196618 267724 196624 267736
rect 196676 267724 196682 267776
rect 219342 267724 219348 267776
rect 219400 267764 219406 267776
rect 261662 267764 261668 267776
rect 219400 267736 261668 267764
rect 219400 267724 219406 267736
rect 261662 267724 261668 267736
rect 261720 267724 261726 267776
rect 42426 267656 42432 267708
rect 42484 267696 42490 267708
rect 122834 267696 122840 267708
rect 42484 267668 122840 267696
rect 42484 267656 42490 267668
rect 122834 267656 122840 267668
rect 122892 267656 122898 267708
rect 158530 267656 158536 267708
rect 158588 267696 158594 267708
rect 206002 267696 206008 267708
rect 158588 267668 206008 267696
rect 158588 267656 158594 267668
rect 206002 267656 206008 267668
rect 206060 267656 206066 267708
rect 357250 267656 357256 267708
rect 357308 267696 357314 267708
rect 357526 267696 357532 267708
rect 357308 267668 357532 267696
rect 357308 267656 357314 267668
rect 357526 267656 357532 267668
rect 357584 267656 357590 267708
rect 361114 267656 361120 267708
rect 361172 267696 361178 267708
rect 458174 267696 458180 267708
rect 361172 267668 458180 267696
rect 361172 267656 361178 267668
rect 458174 267656 458180 267668
rect 458232 267656 458238 267708
rect 47670 267588 47676 267640
rect 47728 267628 47734 267640
rect 53834 267628 53840 267640
rect 47728 267600 53840 267628
rect 47728 267588 47734 267600
rect 53834 267588 53840 267600
rect 53892 267588 53898 267640
rect 55950 267588 55956 267640
rect 56008 267628 56014 267640
rect 129734 267628 129740 267640
rect 56008 267600 129740 267628
rect 56008 267588 56014 267600
rect 129734 267588 129740 267600
rect 129792 267588 129798 267640
rect 153562 267588 153568 267640
rect 153620 267628 153626 267640
rect 200298 267628 200304 267640
rect 153620 267600 200304 267628
rect 153620 267588 153626 267600
rect 200298 267588 200304 267600
rect 200356 267588 200362 267640
rect 216122 267588 216128 267640
rect 216180 267628 216186 267640
rect 302234 267628 302240 267640
rect 216180 267600 302240 267628
rect 216180 267588 216186 267600
rect 302234 267588 302240 267600
rect 302292 267588 302298 267640
rect 362494 267588 362500 267640
rect 362552 267628 362558 267640
rect 455782 267628 455788 267640
rect 362552 267600 455788 267628
rect 362552 267588 362558 267600
rect 455782 267588 455788 267600
rect 455840 267588 455846 267640
rect 57054 267520 57060 267572
rect 57112 267560 57118 267572
rect 128354 267560 128360 267572
rect 57112 267532 128360 267560
rect 57112 267520 57118 267532
rect 128354 267520 128360 267532
rect 128412 267520 128418 267572
rect 155954 267520 155960 267572
rect 156012 267560 156018 267572
rect 202966 267560 202972 267572
rect 156012 267532 202972 267560
rect 156012 267520 156018 267532
rect 202966 267520 202972 267532
rect 203024 267520 203030 267572
rect 206738 267520 206744 267572
rect 206796 267560 206802 267572
rect 276014 267560 276020 267572
rect 206796 267532 276020 267560
rect 206796 267520 206802 267532
rect 276014 267520 276020 267532
rect 276072 267520 276078 267572
rect 364058 267520 364064 267572
rect 364116 267560 364122 267572
rect 445754 267560 445760 267572
rect 364116 267532 445760 267560
rect 364116 267520 364122 267532
rect 445754 267520 445760 267532
rect 445812 267520 445818 267572
rect 56042 267452 56048 267504
rect 56100 267492 56106 267504
rect 125594 267492 125600 267504
rect 56100 267464 125600 267492
rect 56100 267452 56106 267464
rect 125594 267452 125600 267464
rect 125652 267452 125658 267504
rect 163498 267452 163504 267504
rect 163556 267492 163562 267504
rect 197722 267492 197728 267504
rect 163556 267464 197728 267492
rect 163556 267452 163562 267464
rect 197722 267452 197728 267464
rect 197780 267452 197786 267504
rect 202322 267452 202328 267504
rect 202380 267492 202386 267504
rect 270862 267492 270868 267504
rect 202380 267464 270868 267492
rect 202380 267452 202386 267464
rect 270862 267452 270868 267464
rect 270920 267452 270926 267504
rect 370866 267452 370872 267504
rect 370924 267492 370930 267504
rect 449894 267492 449900 267504
rect 370924 267464 449900 267492
rect 370924 267452 370930 267464
rect 449894 267452 449900 267464
rect 449952 267452 449958 267504
rect 54754 267384 54760 267436
rect 54812 267424 54818 267436
rect 120074 267424 120080 267436
rect 54812 267396 120080 267424
rect 54812 267384 54818 267396
rect 120074 267384 120080 267396
rect 120132 267384 120138 267436
rect 166166 267384 166172 267436
rect 166224 267424 166230 267436
rect 200390 267424 200396 267436
rect 166224 267396 200396 267424
rect 166224 267384 166230 267396
rect 200390 267384 200396 267396
rect 200448 267384 200454 267436
rect 203702 267384 203708 267436
rect 203760 267424 203766 267436
rect 268194 267424 268200 267436
rect 203760 267396 268200 267424
rect 203760 267384 203766 267396
rect 268194 267384 268200 267396
rect 268252 267384 268258 267436
rect 369486 267384 369492 267436
rect 369544 267424 369550 267436
rect 447134 267424 447140 267436
rect 369544 267396 447140 267424
rect 369544 267384 369550 267396
rect 447134 267384 447140 267396
rect 447192 267384 447198 267436
rect 46750 267316 46756 267368
rect 46808 267356 46814 267368
rect 51350 267356 51356 267368
rect 46808 267328 51356 267356
rect 46808 267316 46814 267328
rect 51350 267316 51356 267328
rect 51408 267316 51414 267368
rect 53006 267316 53012 267368
rect 53064 267356 53070 267368
rect 117314 267356 117320 267368
rect 53064 267328 117320 267356
rect 53064 267316 53070 267328
rect 117314 267316 117320 267328
rect 117372 267316 117378 267368
rect 160922 267316 160928 267368
rect 160980 267356 160986 267368
rect 207106 267356 207112 267368
rect 160980 267328 207112 267356
rect 160980 267316 160986 267328
rect 207106 267316 207112 267328
rect 207164 267316 207170 267368
rect 213546 267316 213552 267368
rect 213604 267356 213610 267368
rect 273254 267356 273260 267368
rect 213604 267328 273260 267356
rect 213604 267316 213610 267328
rect 273254 267316 273260 267328
rect 273312 267316 273318 267368
rect 356514 267356 356520 267368
rect 354646 267328 356520 267356
rect 53190 267248 53196 267300
rect 53248 267288 53254 267300
rect 115934 267288 115940 267300
rect 53248 267260 115940 267288
rect 53248 267248 53254 267260
rect 115934 267248 115940 267260
rect 115992 267248 115998 267300
rect 204990 267248 204996 267300
rect 205048 267288 205054 267300
rect 263594 267288 263600 267300
rect 205048 267260 263600 267288
rect 205048 267248 205054 267260
rect 263594 267248 263600 267260
rect 263652 267248 263658 267300
rect 53098 267180 53104 267232
rect 53156 267220 53162 267232
rect 113174 267220 113180 267232
rect 53156 267192 113180 267220
rect 53156 267180 53162 267192
rect 113174 267180 113180 267192
rect 113232 267180 113238 267232
rect 207842 267180 207848 267232
rect 207900 267220 207906 267232
rect 260834 267220 260840 267232
rect 207900 267192 260840 267220
rect 207900 267180 207906 267192
rect 260834 267180 260840 267192
rect 260892 267180 260898 267232
rect 343450 267180 343456 267232
rect 343508 267220 343514 267232
rect 354646 267220 354674 267328
rect 356514 267316 356520 267328
rect 356572 267356 356578 267368
rect 356974 267356 356980 267368
rect 356572 267328 356980 267356
rect 356572 267316 356578 267328
rect 356974 267316 356980 267328
rect 357032 267316 357038 267368
rect 358354 267316 358360 267368
rect 358412 267356 358418 267368
rect 435910 267356 435916 267368
rect 358412 267328 435916 267356
rect 358412 267316 358418 267328
rect 435910 267316 435916 267328
rect 435968 267316 435974 267368
rect 361206 267248 361212 267300
rect 361264 267288 361270 267300
rect 437474 267288 437480 267300
rect 361264 267260 437480 267288
rect 361264 267248 361270 267260
rect 437474 267248 437480 267260
rect 437532 267248 437538 267300
rect 343508 267192 354674 267220
rect 343508 267180 343514 267192
rect 356514 267180 356520 267232
rect 356572 267220 356578 267232
rect 356882 267220 356888 267232
rect 356572 267192 356888 267220
rect 356572 267180 356578 267192
rect 356882 267180 356888 267192
rect 356940 267180 356946 267232
rect 372246 267180 372252 267232
rect 372304 267220 372310 267232
rect 442994 267220 443000 267232
rect 372304 267192 443000 267220
rect 372304 267180 372310 267192
rect 442994 267180 443000 267192
rect 443052 267180 443058 267232
rect 51902 267112 51908 267164
rect 51960 267152 51966 267164
rect 104894 267152 104900 267164
rect 51960 267124 104900 267152
rect 51960 267112 51966 267124
rect 104894 267112 104900 267124
rect 104952 267112 104958 267164
rect 183462 267112 183468 267164
rect 183520 267152 183526 267164
rect 196710 267152 196716 267164
rect 183520 267124 196716 267152
rect 183520 267112 183526 267124
rect 196710 267112 196716 267124
rect 196768 267112 196774 267164
rect 211982 267112 211988 267164
rect 212040 267152 212046 267164
rect 265802 267152 265808 267164
rect 212040 267124 265808 267152
rect 212040 267112 212046 267124
rect 265802 267112 265808 267124
rect 265860 267112 265866 267164
rect 278130 267112 278136 267164
rect 278188 267152 278194 267164
rect 356606 267152 356612 267164
rect 278188 267124 356612 267152
rect 278188 267112 278194 267124
rect 356606 267112 356612 267124
rect 356664 267112 356670 267164
rect 373442 267112 373448 267164
rect 373500 267152 373506 267164
rect 440234 267152 440240 267164
rect 373500 267124 440240 267152
rect 373500 267112 373506 267124
rect 440234 267112 440240 267124
rect 440292 267112 440298 267164
rect 503530 267112 503536 267164
rect 503588 267152 503594 267164
rect 517882 267152 517888 267164
rect 503588 267124 517888 267152
rect 503588 267112 503594 267124
rect 517882 267112 517888 267124
rect 517940 267112 517946 267164
rect 47486 267044 47492 267096
rect 47544 267084 47550 267096
rect 47762 267084 47768 267096
rect 47544 267056 47768 267084
rect 47544 267044 47550 267056
rect 47762 267044 47768 267056
rect 47820 267044 47826 267096
rect 51994 267044 52000 267096
rect 52052 267084 52058 267096
rect 103514 267084 103520 267096
rect 52052 267056 103520 267084
rect 52052 267044 52058 267056
rect 103514 267044 103520 267056
rect 103572 267044 103578 267096
rect 206646 267044 206652 267096
rect 206704 267084 206710 267096
rect 258258 267084 258264 267096
rect 206704 267056 258264 267084
rect 206704 267044 206710 267056
rect 258258 267044 258264 267056
rect 258316 267044 258322 267096
rect 343542 267044 343548 267096
rect 343600 267084 343606 267096
rect 357526 267084 357532 267096
rect 343600 267056 357532 267084
rect 343600 267044 343606 267056
rect 357526 267044 357532 267056
rect 357584 267044 357590 267096
rect 369578 267044 369584 267096
rect 369636 267084 369642 267096
rect 416038 267084 416044 267096
rect 369636 267056 416044 267084
rect 369636 267044 369642 267056
rect 416038 267044 416044 267056
rect 416096 267044 416102 267096
rect 50338 266976 50344 267028
rect 50396 267016 50402 267028
rect 100754 267016 100760 267028
rect 50396 266988 100760 267016
rect 50396 266976 50402 266988
rect 100754 266976 100760 266988
rect 100812 266976 100818 267028
rect 183278 266976 183284 267028
rect 183336 267016 183342 267028
rect 197446 267016 197452 267028
rect 183336 266988 197452 267016
rect 183336 266976 183342 266988
rect 197446 266976 197452 266988
rect 197504 266976 197510 267028
rect 214926 266976 214932 267028
rect 214984 267016 214990 267028
rect 273254 267016 273260 267028
rect 214984 266988 273260 267016
rect 214984 266976 214990 266988
rect 273254 266976 273260 266988
rect 273312 266976 273318 267028
rect 277118 266976 277124 267028
rect 277176 267016 277182 267028
rect 356514 267016 356520 267028
rect 277176 266988 356520 267016
rect 277176 266976 277182 266988
rect 356514 266976 356520 266988
rect 356572 266976 356578 267028
rect 365438 266976 365444 267028
rect 365496 267016 365502 267028
rect 409874 267016 409880 267028
rect 365496 266988 409880 267016
rect 365496 266976 365502 266988
rect 409874 266976 409880 266988
rect 409932 266976 409938 267028
rect 503438 266976 503444 267028
rect 503496 267016 503502 267028
rect 517974 267016 517980 267028
rect 503496 266988 517980 267016
rect 503496 266976 503502 266988
rect 517974 266976 517980 266988
rect 518032 266976 518038 267028
rect 54662 266908 54668 266960
rect 54720 266948 54726 266960
rect 88334 266948 88340 266960
rect 54720 266920 88340 266948
rect 54720 266908 54726 266920
rect 88334 266908 88340 266920
rect 88392 266908 88398 266960
rect 210602 266908 210608 266960
rect 210660 266948 210666 266960
rect 255314 266948 255320 266960
rect 210660 266920 255320 266948
rect 210660 266908 210666 266920
rect 255314 266908 255320 266920
rect 255372 266908 255378 266960
rect 379422 266908 379428 266960
rect 379480 266948 379486 266960
rect 422570 266948 422576 266960
rect 379480 266920 422576 266948
rect 379480 266908 379486 266920
rect 422570 266908 422576 266920
rect 422628 266908 422634 266960
rect 47762 266840 47768 266892
rect 47820 266880 47826 266892
rect 80054 266880 80060 266892
rect 47820 266852 80060 266880
rect 47820 266840 47826 266852
rect 80054 266840 80060 266852
rect 80112 266840 80118 266892
rect 213178 266840 213184 266892
rect 213236 266880 213242 266892
rect 252554 266880 252560 266892
rect 213236 266852 252560 266880
rect 213236 266840 213242 266852
rect 252554 266840 252560 266852
rect 252612 266840 252618 266892
rect 375006 266840 375012 266892
rect 375064 266880 375070 266892
rect 412910 266880 412916 266892
rect 375064 266852 412916 266880
rect 375064 266840 375070 266852
rect 412910 266840 412916 266852
rect 412968 266840 412974 266892
rect 47578 266772 47584 266824
rect 47636 266812 47642 266824
rect 77294 266812 77300 266824
rect 47636 266784 77300 266812
rect 47636 266772 47642 266784
rect 77294 266772 77300 266784
rect 77352 266772 77358 266824
rect 219066 266772 219072 266824
rect 219124 266812 219130 266824
rect 247034 266812 247040 266824
rect 219124 266784 247040 266812
rect 219124 266772 219130 266784
rect 247034 266772 247040 266784
rect 247092 266772 247098 266824
rect 376478 266772 376484 266824
rect 376536 266812 376542 266824
rect 407114 266812 407120 266824
rect 376536 266784 407120 266812
rect 376536 266772 376542 266784
rect 407114 266772 407120 266784
rect 407172 266772 407178 266824
rect 214650 266704 214656 266756
rect 214708 266744 214714 266756
rect 310514 266744 310520 266756
rect 214708 266716 310520 266744
rect 214708 266704 214714 266716
rect 310514 266704 310520 266716
rect 310572 266704 310578 266756
rect 214558 266432 214564 266484
rect 214616 266472 214622 266484
rect 214926 266472 214932 266484
rect 214616 266444 214932 266472
rect 214616 266432 214622 266444
rect 214926 266432 214932 266444
rect 214984 266432 214990 266484
rect 214650 266364 214656 266416
rect 214708 266404 214714 266416
rect 215386 266404 215392 266416
rect 214708 266376 215392 266404
rect 214708 266364 214714 266376
rect 215386 266364 215392 266376
rect 215444 266364 215450 266416
rect 356606 266364 356612 266416
rect 356664 266404 356670 266416
rect 356790 266404 356796 266416
rect 356664 266376 356796 266404
rect 356664 266364 356670 266376
rect 356790 266364 356796 266376
rect 356848 266364 356854 266416
rect 425698 266364 425704 266416
rect 425756 266404 425762 266416
rect 434254 266404 434260 266416
rect 425756 266376 434260 266404
rect 425756 266364 425762 266376
rect 434254 266364 434260 266376
rect 434312 266364 434318 266416
rect 517698 266364 517704 266416
rect 517756 266404 517762 266416
rect 517882 266404 517888 266416
rect 517756 266376 517888 266404
rect 517756 266364 517762 266376
rect 517882 266364 517888 266376
rect 517940 266364 517946 266416
rect 50338 266296 50344 266348
rect 50396 266336 50402 266348
rect 57698 266336 57704 266348
rect 50396 266308 57704 266336
rect 50396 266296 50402 266308
rect 57698 266296 57704 266308
rect 57756 266336 57762 266348
rect 92382 266336 92388 266348
rect 57756 266308 92388 266336
rect 57756 266296 57762 266308
rect 92382 266296 92388 266308
rect 92440 266296 92446 266348
rect 215404 266336 215432 266364
rect 262214 266336 262220 266348
rect 215404 266308 262220 266336
rect 262214 266296 262220 266308
rect 262272 266296 262278 266348
rect 379790 266296 379796 266348
rect 379848 266336 379854 266348
rect 403158 266336 403164 266348
rect 379848 266308 403164 266336
rect 379848 266296 379854 266308
rect 403158 266296 403164 266308
rect 403216 266296 403222 266348
rect 63494 266228 63500 266280
rect 63552 266268 63558 266280
rect 92474 266268 92480 266280
rect 63552 266240 92480 266268
rect 63552 266228 63558 266240
rect 92474 266228 92480 266240
rect 92532 266228 92538 266280
rect 218606 266228 218612 266280
rect 218664 266268 218670 266280
rect 219158 266268 219164 266280
rect 218664 266240 219164 266268
rect 218664 266228 218670 266240
rect 219158 266228 219164 266240
rect 219216 266268 219222 266280
rect 252554 266268 252560 266280
rect 219216 266240 252560 266268
rect 219216 266228 219222 266240
rect 252554 266228 252560 266240
rect 252612 266228 252618 266280
rect 378686 266228 378692 266280
rect 378744 266268 378750 266280
rect 411254 266268 411260 266280
rect 378744 266240 411260 266268
rect 378744 266228 378750 266240
rect 411254 266228 411260 266240
rect 411312 266228 411318 266280
rect 54110 266160 54116 266212
rect 54168 266200 54174 266212
rect 84194 266200 84200 266212
rect 54168 266172 84200 266200
rect 54168 266160 54174 266172
rect 84194 266160 84200 266172
rect 84252 266160 84258 266212
rect 216766 266160 216772 266212
rect 216824 266200 216830 266212
rect 218422 266200 218428 266212
rect 216824 266172 218428 266200
rect 216824 266160 216830 266172
rect 218422 266160 218428 266172
rect 218480 266200 218486 266212
rect 251266 266200 251272 266212
rect 218480 266172 251272 266200
rect 218480 266160 218486 266172
rect 251266 266160 251272 266172
rect 251324 266160 251330 266212
rect 379698 266160 379704 266212
rect 379756 266200 379762 266212
rect 409874 266200 409880 266212
rect 379756 266172 409880 266200
rect 379756 266160 379762 266172
rect 409874 266160 409880 266172
rect 409932 266160 409938 266212
rect 58710 266092 58716 266144
rect 58768 266132 58774 266144
rect 89714 266132 89720 266144
rect 58768 266104 89720 266132
rect 58768 266092 58774 266104
rect 89714 266092 89720 266104
rect 89772 266092 89778 266144
rect 213638 266092 213644 266144
rect 213696 266132 213702 266144
rect 245654 266132 245660 266144
rect 213696 266104 245660 266132
rect 213696 266092 213702 266104
rect 245654 266092 245660 266104
rect 245712 266092 245718 266144
rect 371602 266092 371608 266144
rect 371660 266132 371666 266144
rect 372338 266132 372344 266144
rect 371660 266104 372344 266132
rect 371660 266092 371666 266104
rect 372338 266092 372344 266104
rect 372396 266132 372402 266144
rect 401686 266132 401692 266144
rect 372396 266104 401692 266132
rect 372396 266092 372402 266104
rect 401686 266092 401692 266104
rect 401744 266092 401750 266144
rect 53926 266024 53932 266076
rect 53984 266064 53990 266076
rect 85574 266064 85580 266076
rect 53984 266036 85580 266064
rect 53984 266024 53990 266036
rect 85574 266024 85580 266036
rect 85632 266024 85638 266076
rect 219066 266024 219072 266076
rect 219124 266064 219130 266076
rect 219710 266064 219716 266076
rect 219124 266036 219716 266064
rect 219124 266024 219130 266036
rect 219710 266024 219716 266036
rect 219768 266064 219774 266076
rect 251174 266064 251180 266076
rect 219768 266036 251180 266064
rect 219768 266024 219774 266036
rect 251174 266024 251180 266036
rect 251232 266024 251238 266076
rect 379146 266024 379152 266076
rect 379204 266064 379210 266076
rect 407114 266064 407120 266076
rect 379204 266036 407120 266064
rect 379204 266024 379210 266036
rect 407114 266024 407120 266036
rect 407172 266024 407178 266076
rect 85390 265996 85396 266008
rect 52012 265968 85396 265996
rect 52012 265872 52040 265968
rect 85390 265956 85396 265968
rect 85448 265956 85454 266008
rect 220722 265956 220728 266008
rect 220780 265996 220786 266008
rect 249794 265996 249800 266008
rect 220780 265968 249800 265996
rect 220780 265956 220786 265968
rect 249794 265956 249800 265968
rect 249852 265956 249858 266008
rect 373626 265956 373632 266008
rect 373684 265996 373690 266008
rect 400214 265996 400220 266008
rect 373684 265968 400220 265996
rect 373684 265956 373690 265968
rect 400214 265956 400220 265968
rect 400272 265956 400278 266008
rect 54570 265888 54576 265940
rect 54628 265928 54634 265940
rect 56042 265928 56048 265940
rect 54628 265900 56048 265928
rect 54628 265888 54634 265900
rect 56042 265888 56048 265900
rect 56100 265928 56106 265940
rect 88334 265928 88340 265940
rect 56100 265900 88340 265928
rect 56100 265888 56106 265900
rect 88334 265888 88340 265900
rect 88392 265888 88398 265940
rect 213086 265888 213092 265940
rect 213144 265928 213150 265940
rect 213638 265928 213644 265940
rect 213144 265900 213644 265928
rect 213144 265888 213150 265900
rect 213638 265888 213644 265900
rect 213696 265888 213702 265940
rect 219250 265888 219256 265940
rect 219308 265928 219314 265940
rect 219526 265928 219532 265940
rect 219308 265900 219532 265928
rect 219308 265888 219314 265900
rect 219526 265888 219532 265900
rect 219584 265928 219590 265940
rect 248506 265928 248512 265940
rect 219584 265900 248512 265928
rect 219584 265888 219590 265900
rect 248506 265888 248512 265900
rect 248564 265888 248570 265940
rect 376570 265888 376576 265940
rect 376628 265928 376634 265940
rect 377858 265928 377864 265940
rect 376628 265900 377864 265928
rect 376628 265888 376634 265900
rect 377858 265888 377864 265900
rect 377916 265928 377922 265940
rect 404354 265928 404360 265940
rect 377916 265900 404360 265928
rect 377916 265888 377922 265900
rect 404354 265888 404360 265900
rect 404412 265888 404418 265940
rect 50246 265820 50252 265872
rect 50304 265860 50310 265872
rect 51994 265860 52000 265872
rect 50304 265832 52000 265860
rect 50304 265820 50310 265832
rect 51994 265820 52000 265832
rect 52052 265820 52058 265872
rect 78582 265820 78588 265872
rect 78640 265860 78646 265872
rect 111794 265860 111800 265872
rect 78640 265832 111800 265860
rect 78640 265820 78646 265832
rect 111794 265820 111800 265832
rect 111852 265820 111858 265872
rect 244274 265860 244280 265872
rect 216324 265832 244280 265860
rect 57698 265752 57704 265804
rect 57756 265792 57762 265804
rect 91094 265792 91100 265804
rect 57756 265764 91100 265792
rect 57756 265752 57762 265764
rect 91094 265752 91100 265764
rect 91152 265752 91158 265804
rect 216324 265736 216352 265832
rect 244274 265820 244280 265832
rect 244332 265820 244338 265872
rect 370406 265820 370412 265872
rect 370464 265860 370470 265872
rect 372522 265860 372528 265872
rect 370464 265832 372528 265860
rect 370464 265820 370470 265832
rect 372522 265820 372528 265832
rect 372580 265860 372586 265872
rect 398190 265860 398196 265872
rect 372580 265832 398196 265860
rect 372580 265820 372586 265832
rect 398190 265820 398196 265832
rect 398248 265820 398254 265872
rect 247034 265792 247040 265804
rect 216692 265764 247040 265792
rect 52546 265684 52552 265736
rect 52604 265724 52610 265736
rect 100754 265724 100760 265736
rect 52604 265696 100760 265724
rect 52604 265684 52610 265696
rect 100754 265684 100760 265696
rect 100812 265684 100818 265736
rect 215018 265684 215024 265736
rect 215076 265724 215082 265736
rect 216306 265724 216312 265736
rect 215076 265696 216312 265724
rect 215076 265684 215082 265696
rect 216306 265684 216312 265696
rect 216364 265684 216370 265736
rect 52730 265616 52736 265668
rect 52788 265656 52794 265668
rect 113266 265656 113272 265668
rect 52788 265628 113272 265656
rect 52788 265616 52794 265628
rect 113266 265616 113272 265628
rect 113324 265616 113330 265668
rect 214374 265616 214380 265668
rect 214432 265656 214438 265668
rect 216214 265656 216220 265668
rect 214432 265628 216220 265656
rect 214432 265616 214438 265628
rect 216214 265616 216220 265628
rect 216272 265656 216278 265668
rect 216692 265656 216720 265764
rect 247034 265752 247040 265764
rect 247092 265752 247098 265804
rect 367738 265752 367744 265804
rect 367796 265792 367802 265804
rect 370958 265792 370964 265804
rect 367796 265764 370964 265792
rect 367796 265752 367802 265764
rect 370958 265752 370964 265764
rect 371016 265792 371022 265804
rect 398834 265792 398840 265804
rect 371016 265764 398840 265792
rect 371016 265752 371022 265764
rect 398834 265752 398840 265764
rect 398892 265752 398898 265804
rect 217870 265684 217876 265736
rect 217928 265724 217934 265736
rect 219710 265724 219716 265736
rect 217928 265696 219716 265724
rect 217928 265684 217934 265696
rect 219710 265684 219716 265696
rect 219768 265724 219774 265736
rect 265158 265724 265164 265736
rect 219768 265696 265164 265724
rect 219768 265684 219774 265696
rect 265158 265684 265164 265696
rect 265216 265684 265222 265736
rect 373718 265684 373724 265736
rect 373776 265724 373782 265736
rect 376570 265724 376576 265736
rect 373776 265696 376576 265724
rect 373776 265684 373782 265696
rect 376570 265684 376576 265696
rect 376628 265684 376634 265736
rect 376662 265684 376668 265736
rect 376720 265724 376726 265736
rect 378594 265724 378600 265736
rect 376720 265696 378600 265724
rect 376720 265684 376726 265696
rect 378594 265684 378600 265696
rect 378652 265724 378658 265736
rect 408494 265724 408500 265736
rect 378652 265696 408500 265724
rect 378652 265684 378658 265696
rect 408494 265684 408500 265696
rect 408552 265684 408558 265736
rect 267090 265656 267096 265668
rect 216272 265628 216720 265656
rect 219406 265628 267096 265656
rect 216272 265616 216278 265628
rect 214834 265548 214840 265600
rect 214892 265588 214898 265600
rect 218514 265588 218520 265600
rect 214892 265560 218520 265588
rect 214892 265548 214898 265560
rect 218514 265548 218520 265560
rect 218572 265588 218578 265600
rect 219406 265588 219434 265628
rect 267090 265616 267096 265628
rect 267148 265616 267154 265668
rect 371694 265616 371700 265668
rect 371752 265656 371758 265668
rect 373166 265656 373172 265668
rect 371752 265628 373172 265656
rect 371752 265616 371758 265628
rect 373166 265616 373172 265628
rect 373224 265656 373230 265668
rect 405734 265656 405740 265668
rect 373224 265628 405740 265656
rect 373224 265616 373230 265628
rect 405734 265616 405740 265628
rect 405792 265616 405798 265668
rect 218572 265560 219434 265588
rect 218572 265548 218578 265560
rect 377950 265480 377956 265532
rect 378008 265520 378014 265532
rect 411346 265520 411352 265532
rect 378008 265492 411352 265520
rect 378008 265480 378014 265492
rect 411346 265480 411352 265492
rect 411404 265480 411410 265532
rect 375282 265344 375288 265396
rect 375340 265384 375346 265396
rect 375340 265356 383654 265384
rect 375340 265344 375346 265356
rect 375098 265276 375104 265328
rect 375156 265316 375162 265328
rect 379790 265316 379796 265328
rect 375156 265288 379796 265316
rect 375156 265276 375162 265288
rect 379790 265276 379796 265288
rect 379848 265276 379854 265328
rect 375190 265208 375196 265260
rect 375248 265248 375254 265260
rect 379974 265248 379980 265260
rect 375248 265220 379980 265248
rect 375248 265208 375254 265220
rect 379974 265208 379980 265220
rect 380032 265208 380038 265260
rect 377030 265140 377036 265192
rect 377088 265180 377094 265192
rect 377950 265180 377956 265192
rect 377088 265152 377956 265180
rect 377088 265140 377094 265152
rect 377950 265140 377956 265152
rect 378008 265140 378014 265192
rect 212994 265072 213000 265124
rect 213052 265112 213058 265124
rect 215754 265112 215760 265124
rect 213052 265084 215760 265112
rect 213052 265072 213058 265084
rect 215754 265072 215760 265084
rect 215812 265112 215818 265124
rect 230382 265112 230388 265124
rect 215812 265084 230388 265112
rect 215812 265072 215818 265084
rect 230382 265072 230388 265084
rect 230440 265072 230446 265124
rect 375742 265072 375748 265124
rect 375800 265112 375806 265124
rect 379146 265112 379152 265124
rect 375800 265084 379152 265112
rect 375800 265072 375806 265084
rect 379146 265072 379152 265084
rect 379204 265072 379210 265124
rect 212258 265004 212264 265056
rect 212316 265044 212322 265056
rect 215662 265044 215668 265056
rect 212316 265016 215668 265044
rect 212316 265004 212322 265016
rect 215662 265004 215668 265016
rect 215720 265044 215726 265056
rect 233142 265044 233148 265056
rect 215720 265016 233148 265044
rect 215720 265004 215726 265016
rect 233142 265004 233148 265016
rect 233200 265004 233206 265056
rect 377950 265004 377956 265056
rect 378008 265044 378014 265056
rect 379698 265044 379704 265056
rect 378008 265016 379704 265044
rect 378008 265004 378014 265016
rect 379698 265004 379704 265016
rect 379756 265004 379762 265056
rect 210878 264936 210884 264988
rect 210936 264976 210942 264988
rect 214742 264976 214748 264988
rect 210936 264948 214748 264976
rect 210936 264936 210942 264948
rect 214742 264936 214748 264948
rect 214800 264976 214806 264988
rect 231762 264976 231768 264988
rect 214800 264948 231768 264976
rect 214800 264936 214806 264948
rect 231762 264936 231768 264948
rect 231820 264936 231826 264988
rect 374546 264936 374552 264988
rect 374604 264976 374610 264988
rect 375282 264976 375288 264988
rect 374604 264948 375288 264976
rect 374604 264936 374610 264948
rect 375282 264936 375288 264948
rect 375340 264936 375346 264988
rect 378686 264936 378692 264988
rect 378744 264976 378750 264988
rect 379238 264976 379244 264988
rect 378744 264948 379244 264976
rect 378744 264936 378750 264948
rect 379238 264936 379244 264948
rect 379296 264936 379302 264988
rect 383626 264976 383654 265356
rect 391934 264976 391940 264988
rect 383626 264948 391940 264976
rect 391934 264936 391940 264948
rect 391992 264936 391998 264988
rect 48130 264868 48136 264920
rect 48188 264908 48194 264920
rect 54110 264908 54116 264920
rect 48188 264880 54116 264908
rect 48188 264868 48194 264880
rect 54110 264868 54116 264880
rect 54168 264908 54174 264920
rect 54478 264908 54484 264920
rect 54168 264880 54484 264908
rect 54168 264868 54174 264880
rect 54478 264868 54484 264880
rect 54536 264868 54542 264920
rect 212350 264868 212356 264920
rect 212408 264908 212414 264920
rect 272150 264908 272156 264920
rect 212408 264880 272156 264908
rect 212408 264868 212414 264880
rect 272150 264868 272156 264880
rect 272208 264868 272214 264920
rect 378042 264868 378048 264920
rect 378100 264908 378106 264920
rect 416774 264908 416780 264920
rect 378100 264880 416780 264908
rect 378100 264868 378106 264880
rect 416774 264868 416780 264880
rect 416832 264868 416838 264920
rect 45462 264800 45468 264852
rect 45520 264840 45526 264852
rect 58710 264840 58716 264852
rect 45520 264812 58716 264840
rect 45520 264800 45526 264812
rect 58710 264800 58716 264812
rect 58768 264800 58774 264852
rect 219894 264800 219900 264852
rect 219952 264840 219958 264852
rect 253934 264840 253940 264852
rect 219952 264812 253940 264840
rect 219952 264800 219958 264812
rect 253934 264800 253940 264812
rect 253992 264800 253998 264852
rect 379330 264800 379336 264852
rect 379388 264840 379394 264852
rect 412910 264840 412916 264852
rect 379388 264812 412916 264840
rect 379388 264800 379394 264812
rect 412910 264800 412916 264812
rect 412968 264800 412974 264852
rect 43990 264732 43996 264784
rect 44048 264772 44054 264784
rect 57238 264772 57244 264784
rect 44048 264744 57244 264772
rect 44048 264732 44054 264744
rect 57238 264732 57244 264744
rect 57296 264772 57302 264784
rect 57698 264772 57704 264784
rect 57296 264744 57704 264772
rect 57296 264732 57302 264744
rect 57698 264732 57704 264744
rect 57756 264732 57762 264784
rect 230382 264732 230388 264784
rect 230440 264772 230446 264784
rect 259546 264772 259552 264784
rect 230440 264744 259552 264772
rect 230440 264732 230446 264744
rect 259546 264732 259552 264744
rect 259604 264732 259610 264784
rect 369762 264732 369768 264784
rect 369820 264772 369826 264784
rect 378962 264772 378968 264784
rect 369820 264744 378968 264772
rect 369820 264732 369826 264744
rect 378962 264732 378968 264744
rect 379020 264732 379026 264784
rect 388162 264732 388168 264784
rect 388220 264772 388226 264784
rect 420914 264772 420920 264784
rect 388220 264744 420920 264772
rect 388220 264732 388226 264744
rect 420914 264732 420920 264744
rect 420972 264732 420978 264784
rect 43806 264664 43812 264716
rect 43864 264704 43870 264716
rect 52546 264704 52552 264716
rect 43864 264676 52552 264704
rect 43864 264664 43870 264676
rect 52546 264664 52552 264676
rect 52604 264704 52610 264716
rect 53098 264704 53104 264716
rect 52604 264676 53104 264704
rect 52604 264664 52610 264676
rect 53098 264664 53104 264676
rect 53156 264664 53162 264716
rect 233142 264664 233148 264716
rect 233200 264704 233206 264716
rect 259454 264704 259460 264716
rect 233200 264676 259460 264704
rect 233200 264664 233206 264676
rect 259454 264664 259460 264676
rect 259512 264664 259518 264716
rect 389174 264664 389180 264716
rect 389232 264704 389238 264716
rect 419534 264704 419540 264716
rect 389232 264676 419540 264704
rect 389232 264664 389238 264676
rect 419534 264664 419540 264676
rect 419592 264664 419598 264716
rect 46842 264596 46848 264648
rect 46900 264636 46906 264648
rect 53926 264636 53932 264648
rect 46900 264608 53932 264636
rect 46900 264596 46906 264608
rect 53926 264596 53932 264608
rect 53984 264636 53990 264648
rect 54570 264636 54576 264648
rect 53984 264608 54576 264636
rect 53984 264596 53990 264608
rect 54570 264596 54576 264608
rect 54628 264596 54634 264648
rect 231762 264596 231768 264648
rect 231820 264636 231826 264648
rect 256694 264636 256700 264648
rect 231820 264608 256700 264636
rect 231820 264596 231826 264608
rect 256694 264596 256700 264608
rect 256752 264596 256758 264648
rect 390554 264596 390560 264648
rect 390612 264636 390618 264648
rect 418246 264636 418252 264648
rect 390612 264608 418252 264636
rect 390612 264596 390618 264608
rect 418246 264596 418252 264608
rect 418304 264596 418310 264648
rect 46566 264528 46572 264580
rect 46624 264568 46630 264580
rect 147674 264568 147680 264580
rect 46624 264540 147680 264568
rect 46624 264528 46630 264540
rect 147674 264528 147680 264540
rect 147732 264528 147738 264580
rect 391934 264528 391940 264580
rect 391992 264568 391998 264580
rect 418154 264568 418160 264580
rect 391992 264540 418160 264568
rect 391992 264528 391998 264540
rect 418154 264528 418160 264540
rect 418212 264528 418218 264580
rect 43898 264392 43904 264444
rect 43956 264432 43962 264444
rect 47946 264432 47952 264444
rect 43956 264404 47952 264432
rect 43956 264392 43962 264404
rect 47946 264392 47952 264404
rect 48004 264432 48010 264444
rect 63494 264432 63500 264444
rect 48004 264404 63500 264432
rect 48004 264392 48010 264404
rect 63494 264392 63500 264404
rect 63552 264392 63558 264444
rect 45278 264324 45284 264376
rect 45336 264364 45342 264376
rect 47486 264364 47492 264376
rect 45336 264336 47492 264364
rect 45336 264324 45342 264336
rect 47486 264324 47492 264336
rect 47544 264364 47550 264376
rect 78582 264364 78588 264376
rect 47544 264336 78588 264364
rect 47544 264324 47550 264336
rect 78582 264324 78588 264336
rect 78640 264324 78646 264376
rect 210786 264324 210792 264376
rect 210844 264364 210850 264376
rect 215018 264364 215024 264376
rect 210844 264336 215024 264364
rect 210844 264324 210850 264336
rect 215018 264324 215024 264336
rect 215076 264364 215082 264376
rect 244366 264364 244372 264376
rect 215076 264336 244372 264364
rect 215076 264324 215082 264336
rect 244366 264324 244372 264336
rect 244424 264324 244430 264376
rect 43714 264256 43720 264308
rect 43772 264296 43778 264308
rect 49142 264296 49148 264308
rect 43772 264268 49148 264296
rect 43772 264256 43778 264268
rect 49142 264256 49148 264268
rect 49200 264296 49206 264308
rect 82078 264296 82084 264308
rect 49200 264268 82084 264296
rect 49200 264256 49206 264268
rect 82078 264256 82084 264268
rect 82136 264256 82142 264308
rect 208118 264256 208124 264308
rect 208176 264296 208182 264308
rect 214926 264296 214932 264308
rect 208176 264268 214932 264296
rect 208176 264256 208182 264268
rect 214926 264256 214932 264268
rect 214984 264296 214990 264308
rect 269758 264296 269764 264308
rect 214984 264268 269764 264296
rect 214984 264256 214990 264268
rect 269758 264256 269764 264268
rect 269816 264256 269822 264308
rect 43622 264188 43628 264240
rect 43680 264228 43686 264240
rect 47854 264228 47860 264240
rect 43680 264200 47860 264228
rect 43680 264188 43686 264200
rect 47854 264188 47860 264200
rect 47912 264228 47918 264240
rect 96614 264228 96620 264240
rect 47912 264200 96620 264228
rect 47912 264188 47918 264200
rect 96614 264188 96620 264200
rect 96672 264188 96678 264240
rect 209498 264188 209504 264240
rect 209556 264228 209562 264240
rect 213454 264228 213460 264240
rect 209556 264200 213460 264228
rect 209556 264188 209562 264200
rect 213454 264188 213460 264200
rect 213512 264228 213518 264240
rect 271230 264228 271236 264240
rect 213512 264200 271236 264228
rect 213512 264188 213518 264200
rect 271230 264188 271236 264200
rect 271288 264188 271294 264240
rect 377122 263576 377128 263628
rect 377180 263616 377186 263628
rect 378042 263616 378048 263628
rect 377180 263588 378048 263616
rect 377180 263576 377186 263588
rect 378042 263576 378048 263588
rect 378100 263576 378106 263628
rect 378686 263576 378692 263628
rect 378744 263616 378750 263628
rect 379330 263616 379336 263628
rect 378744 263588 379336 263616
rect 378744 263576 378750 263588
rect 379330 263576 379336 263588
rect 379388 263576 379394 263628
rect 376386 263508 376392 263560
rect 376444 263548 376450 263560
rect 436094 263548 436100 263560
rect 376444 263520 436100 263548
rect 376444 263508 376450 263520
rect 436094 263508 436100 263520
rect 436152 263508 436158 263560
rect 378042 263440 378048 263492
rect 378100 263480 378106 263492
rect 437474 263480 437480 263492
rect 378100 263452 437480 263480
rect 378100 263440 378106 263452
rect 437474 263440 437480 263452
rect 437532 263440 437538 263492
rect 375834 263100 375840 263152
rect 375892 263140 375898 263152
rect 376386 263140 376392 263152
rect 375892 263112 376392 263140
rect 375892 263100 375898 263112
rect 376386 263100 376392 263112
rect 376444 263100 376450 263152
rect 357434 252560 357440 252612
rect 357492 252560 357498 252612
rect 356882 252492 356888 252544
rect 356940 252532 356946 252544
rect 357452 252532 357480 252560
rect 356940 252504 357480 252532
rect 356940 252492 356946 252504
rect 357434 251240 357440 251252
rect 356440 251212 357440 251240
rect 213178 251132 213184 251184
rect 213236 251172 213242 251184
rect 215294 251172 215300 251184
rect 213236 251144 215300 251172
rect 213236 251132 213242 251144
rect 215294 251132 215300 251144
rect 215352 251132 215358 251184
rect 215846 251132 215852 251184
rect 215904 251172 215910 251184
rect 263594 251172 263600 251184
rect 215904 251144 263600 251172
rect 215904 251132 215910 251144
rect 263594 251132 263600 251144
rect 263652 251132 263658 251184
rect 340230 251132 340236 251184
rect 340288 251172 340294 251184
rect 356440 251172 356468 251212
rect 357434 251200 357440 251212
rect 357492 251200 357498 251252
rect 340288 251144 356468 251172
rect 340288 251132 340294 251144
rect 368382 251132 368388 251184
rect 368440 251172 368446 251184
rect 371786 251172 371792 251184
rect 368440 251144 371792 251172
rect 368440 251132 368446 251144
rect 371786 251132 371792 251144
rect 371844 251132 371850 251184
rect 373442 251132 373448 251184
rect 373500 251172 373506 251184
rect 373810 251172 373816 251184
rect 373500 251144 373816 251172
rect 373500 251132 373506 251144
rect 373810 251132 373816 251144
rect 373868 251172 373874 251184
rect 430574 251172 430580 251184
rect 373868 251144 430580 251172
rect 373868 251132 373874 251144
rect 430574 251132 430580 251144
rect 430632 251132 430638 251184
rect 217134 251064 217140 251116
rect 217192 251104 217198 251116
rect 217962 251104 217968 251116
rect 217192 251076 217968 251104
rect 217192 251064 217198 251076
rect 217962 251064 217968 251076
rect 218020 251104 218026 251116
rect 236638 251104 236644 251116
rect 218020 251076 236644 251104
rect 218020 251064 218026 251076
rect 236638 251064 236644 251076
rect 236696 251064 236702 251116
rect 372246 251064 372252 251116
rect 372304 251104 372310 251116
rect 372430 251104 372436 251116
rect 372304 251076 372436 251104
rect 372304 251064 372310 251076
rect 372430 251064 372436 251076
rect 372488 251104 372494 251116
rect 421558 251104 421564 251116
rect 372488 251076 421564 251104
rect 372488 251064 372494 251076
rect 421558 251064 421564 251076
rect 421616 251064 421622 251116
rect 517606 251064 517612 251116
rect 517664 251104 517670 251116
rect 517882 251104 517888 251116
rect 517664 251076 517888 251104
rect 517664 251064 517670 251076
rect 517882 251064 517888 251076
rect 517940 251064 517946 251116
rect 197354 250928 197360 250980
rect 197412 250968 197418 250980
rect 197538 250968 197544 250980
rect 197412 250940 197544 250968
rect 197412 250928 197418 250940
rect 197538 250928 197544 250940
rect 197596 250928 197602 250980
rect 371142 250724 371148 250776
rect 371200 250764 371206 250776
rect 374454 250764 374460 250776
rect 371200 250736 374460 250764
rect 371200 250724 371206 250736
rect 374454 250724 374460 250736
rect 374512 250764 374518 250776
rect 425698 250764 425704 250776
rect 374512 250736 425704 250764
rect 374512 250724 374518 250736
rect 425698 250724 425704 250736
rect 425756 250724 425762 250776
rect 371050 250656 371056 250708
rect 371108 250696 371114 250708
rect 373534 250696 373540 250708
rect 371108 250668 373540 250696
rect 371108 250656 371114 250668
rect 373534 250656 373540 250668
rect 373592 250696 373598 250708
rect 430666 250696 430672 250708
rect 373592 250668 430672 250696
rect 373592 250656 373598 250668
rect 430666 250656 430672 250668
rect 430724 250656 430730 250708
rect 180242 250588 180248 250640
rect 180300 250628 180306 250640
rect 197630 250628 197636 250640
rect 180300 250600 197636 250628
rect 180300 250588 180306 250600
rect 197630 250588 197636 250600
rect 197688 250588 197694 250640
rect 371786 250588 371792 250640
rect 371844 250628 371850 250640
rect 429194 250628 429200 250640
rect 371844 250600 429200 250628
rect 371844 250588 371850 250600
rect 429194 250588 429200 250600
rect 429252 250588 429258 250640
rect 500402 250588 500408 250640
rect 500460 250628 500466 250640
rect 517882 250628 517888 250640
rect 500460 250600 517888 250628
rect 500460 250588 500466 250600
rect 517882 250588 517888 250600
rect 517940 250588 517946 250640
rect 82814 250520 82820 250572
rect 82872 250560 82878 250572
rect 100846 250560 100852 250572
rect 82872 250532 100852 250560
rect 82872 250520 82878 250532
rect 100846 250520 100852 250532
rect 100904 250520 100910 250572
rect 209590 250520 209596 250572
rect 209648 250560 209654 250572
rect 209648 250532 219434 250560
rect 209648 250520 209654 250532
rect 67542 250452 67548 250504
rect 67600 250492 67606 250504
rect 97994 250492 98000 250504
rect 67600 250464 98000 250492
rect 67600 250452 67606 250464
rect 97994 250452 98000 250464
rect 98052 250452 98058 250504
rect 179322 250452 179328 250504
rect 179380 250492 179386 250504
rect 197538 250492 197544 250504
rect 179380 250464 197544 250492
rect 179380 250452 179386 250464
rect 197538 250452 197544 250464
rect 197596 250452 197602 250504
rect 219406 250492 219434 250532
rect 338482 250520 338488 250572
rect 338540 250560 338546 250572
rect 356882 250560 356888 250572
rect 338540 250532 356888 250560
rect 338540 250520 338546 250532
rect 356882 250520 356888 250532
rect 356940 250520 356946 250572
rect 362862 250520 362868 250572
rect 362920 250560 362926 250572
rect 372430 250560 372436 250572
rect 362920 250532 372436 250560
rect 362920 250520 362926 250532
rect 372430 250520 372436 250532
rect 372488 250560 372494 250572
rect 438854 250560 438860 250572
rect 372488 250532 438860 250560
rect 372488 250520 372494 250532
rect 438854 250520 438860 250532
rect 438912 250520 438918 250572
rect 499022 250520 499028 250572
rect 499080 250560 499086 250572
rect 517790 250560 517796 250572
rect 499080 250532 517796 250560
rect 499080 250520 499086 250532
rect 517790 250520 517796 250532
rect 517848 250520 517854 250572
rect 219618 250492 219624 250504
rect 219406 250464 219624 250492
rect 219618 250452 219624 250464
rect 219676 250492 219682 250504
rect 267734 250492 267740 250504
rect 219676 250464 267740 250492
rect 219676 250452 219682 250464
rect 267734 250452 267740 250464
rect 267792 250452 267798 250504
rect 279970 250452 279976 250504
rect 280028 250492 280034 250504
rect 357618 250492 357624 250504
rect 280028 250464 357624 250492
rect 280028 250452 280034 250464
rect 357618 250452 357624 250464
rect 357676 250452 357682 250504
rect 379698 250452 379704 250504
rect 379756 250492 379762 250504
rect 396074 250492 396080 250504
rect 379756 250464 396080 250492
rect 379756 250452 379762 250464
rect 396074 250452 396080 250464
rect 396132 250452 396138 250504
rect 510890 249840 510896 249892
rect 510948 249880 510954 249892
rect 517514 249880 517520 249892
rect 510948 249852 517520 249880
rect 510948 249840 510954 249852
rect 517514 249840 517520 249852
rect 517572 249840 517578 249892
rect 190914 249772 190920 249824
rect 190972 249812 190978 249824
rect 213178 249812 213184 249824
rect 190972 249784 213184 249812
rect 190972 249772 190978 249784
rect 213178 249772 213184 249784
rect 213236 249772 213242 249824
rect 350994 249772 351000 249824
rect 351052 249812 351058 249824
rect 369118 249812 369124 249824
rect 351052 249784 369124 249812
rect 351052 249772 351058 249784
rect 369118 249772 369124 249784
rect 369176 249812 369182 249824
rect 376018 249812 376024 249824
rect 369176 249784 376024 249812
rect 369176 249772 369182 249784
rect 376018 249772 376024 249784
rect 376076 249772 376082 249824
rect 50430 249704 50436 249756
rect 50488 249744 50494 249756
rect 52730 249744 52736 249756
rect 50488 249716 52736 249744
rect 50488 249704 50494 249716
rect 52730 249704 52736 249716
rect 52788 249704 52794 249756
rect 58434 249704 58440 249756
rect 58492 249744 58498 249756
rect 60918 249744 60924 249756
rect 58492 249716 60924 249744
rect 58492 249704 58498 249716
rect 60918 249704 60924 249716
rect 60976 249704 60982 249756
rect 58526 249636 58532 249688
rect 58584 249676 58590 249688
rect 60826 249676 60832 249688
rect 58584 249648 60832 249676
rect 58584 249636 58590 249648
rect 60826 249636 60832 249648
rect 60884 249636 60890 249688
rect 55950 249364 55956 249416
rect 56008 249404 56014 249416
rect 61010 249404 61016 249416
rect 56008 249376 61016 249404
rect 56008 249364 56014 249376
rect 61010 249364 61016 249376
rect 61068 249364 61074 249416
rect 54662 249160 54668 249212
rect 54720 249200 54726 249212
rect 60734 249200 60740 249212
rect 54720 249172 60740 249200
rect 54720 249160 54726 249172
rect 60734 249160 60740 249172
rect 60792 249160 60798 249212
rect 52730 249092 52736 249144
rect 52788 249132 52794 249144
rect 67542 249132 67548 249144
rect 52788 249104 67548 249132
rect 52788 249092 52794 249104
rect 67542 249092 67548 249104
rect 67600 249092 67606 249144
rect 53006 249024 53012 249076
rect 53064 249064 53070 249076
rect 82814 249064 82820 249076
rect 53064 249036 82820 249064
rect 53064 249024 53070 249036
rect 82814 249024 82820 249036
rect 82872 249024 82878 249076
rect 42702 248344 42708 248396
rect 42760 248384 42766 248396
rect 52914 248384 52920 248396
rect 42760 248356 52920 248384
rect 42760 248344 42766 248356
rect 52914 248344 52920 248356
rect 52972 248344 52978 248396
rect 52730 243652 52736 243704
rect 52788 243692 52794 243704
rect 53006 243692 53012 243704
rect 52788 243664 53012 243692
rect 52788 243652 52794 243664
rect 53006 243652 53012 243664
rect 53064 243652 53070 243704
rect 52822 243584 52828 243636
rect 52880 243584 52886 243636
rect 52840 243432 52868 243584
rect 52822 243380 52828 243432
rect 52880 243380 52886 243432
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 40678 202824 40684 202836
rect 3108 202796 40684 202824
rect 3108 202784 3114 202796
rect 40678 202784 40684 202796
rect 40736 202784 40742 202836
rect 520182 182180 520188 182232
rect 520240 182220 520246 182232
rect 580258 182220 580264 182232
rect 520240 182192 580264 182220
rect 520240 182180 520246 182192
rect 580258 182180 580264 182192
rect 580316 182180 580322 182232
rect 519262 182112 519268 182164
rect 519320 182152 519326 182164
rect 519446 182152 519452 182164
rect 519320 182124 519452 182152
rect 519320 182112 519326 182124
rect 519446 182112 519452 182124
rect 519504 182152 519510 182164
rect 580350 182152 580356 182164
rect 519504 182124 580356 182152
rect 519504 182112 519510 182124
rect 580350 182112 580356 182124
rect 580408 182112 580414 182164
rect 207750 175176 207756 175228
rect 207808 175216 207814 175228
rect 216674 175216 216680 175228
rect 207808 175188 216680 175216
rect 207808 175176 207814 175188
rect 216674 175176 216680 175188
rect 216732 175176 216738 175228
rect 363966 175176 363972 175228
rect 364024 175216 364030 175228
rect 376846 175216 376852 175228
rect 364024 175188 376852 175216
rect 364024 175176 364030 175188
rect 376846 175176 376852 175188
rect 376904 175176 376910 175228
rect 369118 173816 369124 173868
rect 369176 173856 369182 173868
rect 376846 173856 376852 173868
rect 369176 173828 376852 173856
rect 369176 173816 369182 173828
rect 376846 173816 376852 173828
rect 376904 173816 376910 173868
rect 203518 173748 203524 173800
rect 203576 173788 203582 173800
rect 217042 173788 217048 173800
rect 203576 173760 217048 173788
rect 203576 173748 203582 173760
rect 217042 173748 217048 173760
rect 217100 173748 217106 173800
rect 372154 173748 372160 173800
rect 372212 173788 372218 173800
rect 376754 173788 376760 173800
rect 372212 173760 376760 173788
rect 372212 173748 372218 173760
rect 376754 173748 376760 173760
rect 376812 173748 376818 173800
rect 197998 173136 198004 173188
rect 198056 173176 198062 173188
rect 213178 173176 213184 173188
rect 198056 173148 213184 173176
rect 198056 173136 198062 173148
rect 213178 173136 213184 173148
rect 213236 173176 213242 173188
rect 216674 173176 216680 173188
rect 213236 173148 216680 173176
rect 213236 173136 213242 173148
rect 216674 173136 216680 173148
rect 216732 173136 216738 173188
rect 358722 173136 358728 173188
rect 358780 173176 358786 173188
rect 369118 173176 369124 173188
rect 358780 173148 369124 173176
rect 358780 173136 358786 173148
rect 369118 173136 369124 173148
rect 369176 173136 369182 173188
rect 374454 165520 374460 165572
rect 374512 165560 374518 165572
rect 375558 165560 375564 165572
rect 374512 165532 375564 165560
rect 374512 165520 374518 165532
rect 375558 165520 375564 165532
rect 375616 165520 375622 165572
rect 375558 164432 375564 164484
rect 375616 164472 375622 164484
rect 434346 164472 434352 164484
rect 375616 164444 434352 164472
rect 375616 164432 375622 164444
rect 434346 164432 434352 164444
rect 434404 164432 434410 164484
rect 50522 164364 50528 164416
rect 50580 164404 50586 164416
rect 96062 164404 96068 164416
rect 50580 164376 96068 164404
rect 50580 164364 50586 164376
rect 96062 164364 96068 164376
rect 96120 164364 96126 164416
rect 363782 164364 363788 164416
rect 363840 164404 363846 164416
rect 425974 164404 425980 164416
rect 363840 164376 425980 164404
rect 363840 164364 363846 164376
rect 425974 164364 425980 164376
rect 426032 164364 426038 164416
rect 59078 164296 59084 164348
rect 59136 164336 59142 164348
rect 140866 164336 140872 164348
rect 59136 164308 140872 164336
rect 59136 164296 59142 164308
rect 140866 164296 140872 164308
rect 140924 164296 140930 164348
rect 205082 164296 205088 164348
rect 205140 164336 205146 164348
rect 258442 164336 258448 164348
rect 205140 164308 258448 164336
rect 205140 164296 205146 164308
rect 258442 164296 258448 164308
rect 258500 164296 258506 164348
rect 366726 164296 366732 164348
rect 366784 164336 366790 164348
rect 450998 164336 451004 164348
rect 366784 164308 451004 164336
rect 366784 164296 366790 164308
rect 450998 164296 451004 164308
rect 451056 164296 451062 164348
rect 41046 164228 41052 164280
rect 41104 164268 41110 164280
rect 163314 164268 163320 164280
rect 41104 164240 163320 164268
rect 41104 164228 41110 164240
rect 163314 164228 163320 164240
rect 163372 164228 163378 164280
rect 202230 164228 202236 164280
rect 202288 164268 202294 164280
rect 318426 164268 318432 164280
rect 202288 164240 318432 164268
rect 202288 164228 202294 164240
rect 318426 164228 318432 164240
rect 318484 164228 318490 164280
rect 362402 164228 362408 164280
rect 362460 164268 362466 164280
rect 480898 164268 480904 164280
rect 362460 164240 480904 164268
rect 362460 164228 362466 164240
rect 480898 164228 480904 164240
rect 480956 164228 480962 164280
rect 375834 164160 375840 164212
rect 375892 164200 375898 164212
rect 376386 164200 376392 164212
rect 375892 164172 376392 164200
rect 375892 164160 375898 164172
rect 376386 164160 376392 164172
rect 376444 164160 376450 164212
rect 374546 164092 374552 164144
rect 374604 164132 374610 164144
rect 393314 164132 393320 164144
rect 374604 164104 393320 164132
rect 374604 164092 374610 164104
rect 393314 164092 393320 164104
rect 393372 164132 393378 164144
rect 394510 164132 394516 164144
rect 393372 164104 394516 164132
rect 393372 164092 393378 164104
rect 394510 164092 394516 164104
rect 394568 164092 394574 164144
rect 49418 164024 49424 164076
rect 49476 164064 49482 164076
rect 98454 164064 98460 164076
rect 49476 164036 98460 164064
rect 49476 164024 49482 164036
rect 98454 164024 98460 164036
rect 98512 164024 98518 164076
rect 365162 164024 365168 164076
rect 365220 164064 365226 164076
rect 423490 164064 423496 164076
rect 365220 164036 423496 164064
rect 365220 164024 365226 164036
rect 423490 164024 423496 164036
rect 423548 164024 423554 164076
rect 52086 163956 52092 164008
rect 52144 163996 52150 164008
rect 101030 163996 101036 164008
rect 52144 163968 101036 163996
rect 52144 163956 52150 163968
rect 101030 163956 101036 163968
rect 101088 163956 101094 164008
rect 362310 163956 362316 164008
rect 362368 163996 362374 164008
rect 421006 163996 421012 164008
rect 362368 163968 421012 163996
rect 362368 163956 362374 163968
rect 421006 163956 421012 163968
rect 421064 163956 421070 164008
rect 50798 163888 50804 163940
rect 50856 163928 50862 163940
rect 103514 163928 103520 163940
rect 50856 163900 103520 163928
rect 50856 163888 50862 163900
rect 103514 163888 103520 163900
rect 103572 163888 103578 163940
rect 356698 163888 356704 163940
rect 356756 163928 356762 163940
rect 416038 163928 416044 163940
rect 356756 163900 416044 163928
rect 356756 163888 356762 163900
rect 416038 163888 416044 163900
rect 416096 163888 416102 163940
rect 52178 163820 52184 163872
rect 52236 163860 52242 163872
rect 105906 163860 105912 163872
rect 52236 163832 105912 163860
rect 52236 163820 52242 163832
rect 105906 163820 105912 163832
rect 105964 163820 105970 163872
rect 366634 163820 366640 163872
rect 366692 163860 366698 163872
rect 428182 163860 428188 163872
rect 366692 163832 428188 163860
rect 366692 163820 366698 163832
rect 428182 163820 428188 163832
rect 428240 163820 428246 163872
rect 50706 163752 50712 163804
rect 50764 163792 50770 163804
rect 108206 163792 108212 163804
rect 50764 163764 108212 163792
rect 50764 163752 50770 163764
rect 108206 163752 108212 163764
rect 108264 163752 108270 163804
rect 116210 163752 116216 163804
rect 116268 163792 116274 163804
rect 117038 163792 117044 163804
rect 116268 163764 117044 163792
rect 116268 163752 116274 163764
rect 117038 163752 117044 163764
rect 117096 163792 117102 163804
rect 196618 163792 196624 163804
rect 117096 163764 196624 163792
rect 117096 163752 117102 163764
rect 196618 163752 196624 163764
rect 196676 163752 196682 163804
rect 369302 163752 369308 163804
rect 369360 163792 369366 163804
rect 430942 163792 430948 163804
rect 369360 163764 430948 163792
rect 369360 163752 369366 163764
rect 430942 163752 430948 163764
rect 431000 163752 431006 163804
rect 59998 163684 60004 163736
rect 60056 163724 60062 163736
rect 145926 163724 145932 163736
rect 60056 163696 145932 163724
rect 60056 163684 60062 163696
rect 145926 163684 145932 163696
rect 145984 163684 145990 163736
rect 213362 163684 213368 163736
rect 213420 163724 213426 163736
rect 261018 163724 261024 163736
rect 213420 163696 261024 163724
rect 213420 163684 213426 163696
rect 261018 163684 261024 163696
rect 261076 163684 261082 163736
rect 369394 163684 369400 163736
rect 369452 163724 369458 163736
rect 470594 163724 470600 163736
rect 369452 163696 470600 163724
rect 369452 163684 369458 163696
rect 470594 163684 470600 163696
rect 470652 163684 470658 163736
rect 59170 163616 59176 163668
rect 59228 163656 59234 163668
rect 148502 163656 148508 163668
rect 59228 163628 148508 163656
rect 59228 163616 59234 163628
rect 148502 163616 148508 163628
rect 148560 163616 148566 163668
rect 209130 163616 209136 163668
rect 209188 163656 209194 163668
rect 298462 163656 298468 163668
rect 209188 163628 298468 163656
rect 209188 163616 209194 163628
rect 298462 163616 298468 163628
rect 298520 163616 298526 163668
rect 372062 163616 372068 163668
rect 372120 163656 372126 163668
rect 473446 163656 473452 163668
rect 372120 163628 473452 163656
rect 372120 163616 372126 163628
rect 473446 163616 473452 163628
rect 473504 163616 473510 163668
rect 510522 163616 510528 163668
rect 510580 163656 510586 163668
rect 517514 163656 517520 163668
rect 510580 163628 517520 163656
rect 510580 163616 510586 163628
rect 517514 163616 517520 163628
rect 517572 163616 517578 163668
rect 59906 163548 59912 163600
rect 59964 163588 59970 163600
rect 150894 163588 150900 163600
rect 59964 163560 150900 163588
rect 59964 163548 59970 163560
rect 150894 163548 150900 163560
rect 150952 163548 150958 163600
rect 211890 163548 211896 163600
rect 211948 163588 211954 163600
rect 305914 163588 305920 163600
rect 211948 163560 305920 163588
rect 211948 163548 211954 163560
rect 305914 163548 305920 163560
rect 305972 163548 305978 163600
rect 373350 163548 373356 163600
rect 373408 163588 373414 163600
rect 475838 163588 475844 163600
rect 373408 163560 475844 163588
rect 373408 163548 373414 163560
rect 475838 163548 475844 163560
rect 475896 163548 475902 163600
rect 58894 163480 58900 163532
rect 58952 163520 58958 163532
rect 153378 163520 153384 163532
rect 58952 163492 153384 163520
rect 58952 163480 58958 163492
rect 153378 163480 153384 163492
rect 153436 163480 153442 163532
rect 206370 163480 206376 163532
rect 206428 163520 206434 163532
rect 300854 163520 300860 163532
rect 206428 163492 300860 163520
rect 206428 163480 206434 163492
rect 300854 163480 300860 163492
rect 300912 163480 300918 163532
rect 368106 163480 368112 163532
rect 368164 163520 368170 163532
rect 478414 163520 478420 163532
rect 368164 163492 478420 163520
rect 368164 163480 368170 163492
rect 478414 163480 478420 163492
rect 478472 163480 478478 163532
rect 196710 163412 196716 163464
rect 196768 163452 196774 163464
rect 197354 163452 197360 163464
rect 196768 163424 197360 163452
rect 196768 163412 196774 163424
rect 197354 163412 197360 163424
rect 197412 163412 197418 163464
rect 377122 163140 377128 163192
rect 377180 163180 377186 163192
rect 396718 163180 396724 163192
rect 377180 163152 396724 163180
rect 377180 163140 377186 163152
rect 396718 163140 396724 163152
rect 396776 163140 396782 163192
rect 394510 163072 394516 163124
rect 394568 163112 394574 163124
rect 415302 163112 415308 163124
rect 394568 163084 415308 163112
rect 394568 163072 394574 163084
rect 415302 163072 415308 163084
rect 415360 163072 415366 163124
rect 374914 163004 374920 163056
rect 374972 163044 374978 163056
rect 431954 163044 431960 163056
rect 374972 163016 431960 163044
rect 374972 163004 374978 163016
rect 431954 163004 431960 163016
rect 432012 163004 432018 163056
rect 378410 162936 378416 162988
rect 378468 162976 378474 162988
rect 438026 162976 438032 162988
rect 378468 162948 438032 162976
rect 378468 162936 378474 162948
rect 438026 162936 438032 162948
rect 438084 162936 438090 162988
rect 52914 162868 52920 162920
rect 52972 162908 52978 162920
rect 54386 162908 54392 162920
rect 52972 162880 54392 162908
rect 52972 162868 52978 162880
rect 54386 162868 54392 162880
rect 54444 162908 54450 162920
rect 73798 162908 73804 162920
rect 54444 162880 73804 162908
rect 54444 162868 54450 162880
rect 73798 162868 73804 162880
rect 73856 162868 73862 162920
rect 218238 162868 218244 162920
rect 218296 162908 218302 162920
rect 218514 162908 218520 162920
rect 218296 162880 218520 162908
rect 218296 162868 218302 162880
rect 218514 162868 218520 162880
rect 218572 162908 218578 162920
rect 267550 162908 267556 162920
rect 218572 162880 267556 162908
rect 218572 162868 218578 162880
rect 267550 162868 267556 162880
rect 267608 162868 267614 162920
rect 376386 162868 376392 162920
rect 376444 162908 376450 162920
rect 436922 162908 436928 162920
rect 376444 162880 436928 162908
rect 376444 162868 376450 162880
rect 436922 162868 436928 162880
rect 436980 162868 436986 162920
rect 55122 162800 55128 162852
rect 55180 162840 55186 162852
rect 133414 162840 133420 162852
rect 55180 162812 133420 162840
rect 55180 162800 55186 162812
rect 133414 162800 133420 162812
rect 133472 162800 133478 162852
rect 209038 162800 209044 162852
rect 209096 162840 209102 162852
rect 320910 162840 320916 162852
rect 209096 162812 320916 162840
rect 209096 162800 209102 162812
rect 320910 162800 320916 162812
rect 320968 162800 320974 162852
rect 356698 162800 356704 162852
rect 356756 162840 356762 162852
rect 356974 162840 356980 162852
rect 356756 162812 356980 162840
rect 356756 162800 356762 162812
rect 356974 162800 356980 162812
rect 357032 162800 357038 162852
rect 415302 162800 415308 162852
rect 415360 162840 415366 162852
rect 418154 162840 418160 162852
rect 415360 162812 418160 162840
rect 415360 162800 415366 162812
rect 418154 162800 418160 162812
rect 418212 162800 418218 162852
rect 517606 162800 517612 162852
rect 517664 162840 517670 162852
rect 517974 162840 517980 162852
rect 517664 162812 517980 162840
rect 517664 162800 517670 162812
rect 517974 162800 517980 162812
rect 518032 162800 518038 162852
rect 56226 162732 56232 162784
rect 56284 162772 56290 162784
rect 130838 162772 130844 162784
rect 56284 162744 130844 162772
rect 56284 162732 56290 162744
rect 130838 162732 130844 162744
rect 130896 162732 130902 162784
rect 204898 162732 204904 162784
rect 204956 162772 204962 162784
rect 308582 162772 308588 162784
rect 204956 162744 308588 162772
rect 204956 162732 204962 162744
rect 308582 162732 308588 162744
rect 308640 162732 308646 162784
rect 365254 162732 365260 162784
rect 365312 162772 365318 162784
rect 455782 162772 455788 162784
rect 365312 162744 455788 162772
rect 365312 162732 365318 162744
rect 455782 162732 455788 162744
rect 455840 162732 455846 162784
rect 54846 162664 54852 162716
rect 54904 162704 54910 162716
rect 128354 162704 128360 162716
rect 54904 162676 128360 162704
rect 54904 162664 54910 162676
rect 128354 162664 128360 162676
rect 128412 162664 128418 162716
rect 207658 162664 207664 162716
rect 207716 162704 207722 162716
rect 303430 162704 303436 162716
rect 207716 162676 303436 162704
rect 207716 162664 207722 162676
rect 303430 162664 303436 162676
rect 303488 162664 303494 162716
rect 370682 162664 370688 162716
rect 370740 162704 370746 162716
rect 458358 162704 458364 162716
rect 370740 162676 458364 162704
rect 370740 162664 370746 162676
rect 458358 162664 458364 162676
rect 458416 162664 458422 162716
rect 56134 162596 56140 162648
rect 56192 162636 56198 162648
rect 125870 162636 125876 162648
rect 56192 162608 125876 162636
rect 56192 162596 56198 162608
rect 125870 162596 125876 162608
rect 125928 162596 125934 162648
rect 218882 162596 218888 162648
rect 218940 162636 218946 162648
rect 293310 162636 293316 162648
rect 218940 162608 293316 162636
rect 218940 162596 218946 162608
rect 293310 162596 293316 162608
rect 293368 162596 293374 162648
rect 363874 162596 363880 162648
rect 363932 162636 363938 162648
rect 448238 162636 448244 162648
rect 363932 162608 448244 162636
rect 363932 162596 363938 162608
rect 448238 162596 448244 162608
rect 448296 162596 448302 162648
rect 55030 162528 55036 162580
rect 55088 162568 55094 162580
rect 122834 162568 122840 162580
rect 55088 162540 122840 162568
rect 55088 162528 55094 162540
rect 122834 162528 122840 162540
rect 122892 162528 122898 162580
rect 211798 162528 211804 162580
rect 211856 162568 211862 162580
rect 283742 162568 283748 162580
rect 211856 162540 283748 162568
rect 211856 162528 211862 162540
rect 283742 162528 283748 162540
rect 283800 162528 283806 162580
rect 371970 162528 371976 162580
rect 372028 162568 372034 162580
rect 445846 162568 445852 162580
rect 372028 162540 445852 162568
rect 372028 162528 372034 162540
rect 445846 162528 445852 162540
rect 445904 162528 445910 162580
rect 53374 162460 53380 162512
rect 53432 162500 53438 162512
rect 120718 162500 120724 162512
rect 53432 162472 120724 162500
rect 53432 162460 53438 162472
rect 120718 162460 120724 162472
rect 120776 162460 120782 162512
rect 215938 162460 215944 162512
rect 215996 162500 216002 162512
rect 285950 162500 285956 162512
rect 215996 162472 285956 162500
rect 215996 162460 216002 162472
rect 285950 162460 285956 162472
rect 286008 162460 286014 162512
rect 369210 162460 369216 162512
rect 369268 162500 369274 162512
rect 440878 162500 440884 162512
rect 369268 162472 440884 162500
rect 369268 162460 369274 162472
rect 440878 162460 440884 162472
rect 440936 162460 440942 162512
rect 53282 162392 53288 162444
rect 53340 162432 53346 162444
rect 115934 162432 115940 162444
rect 53340 162404 115940 162432
rect 53340 162392 53346 162404
rect 115934 162392 115940 162404
rect 115992 162392 115998 162444
rect 210510 162392 210516 162444
rect 210568 162432 210574 162444
rect 278406 162432 278412 162444
rect 210568 162404 278412 162432
rect 210568 162392 210574 162404
rect 278406 162392 278412 162404
rect 278464 162392 278470 162444
rect 368014 162392 368020 162444
rect 368072 162432 368078 162444
rect 438486 162432 438492 162444
rect 368072 162404 438492 162432
rect 368072 162392 368078 162404
rect 438486 162392 438492 162404
rect 438544 162392 438550 162444
rect 56410 162324 56416 162376
rect 56468 162364 56474 162376
rect 118326 162364 118332 162376
rect 56468 162336 118332 162364
rect 56468 162324 56474 162336
rect 118326 162324 118332 162336
rect 118384 162324 118390 162376
rect 206462 162324 206468 162376
rect 206520 162364 206526 162376
rect 268286 162364 268292 162376
rect 206520 162336 268292 162364
rect 206520 162324 206526 162336
rect 268286 162324 268292 162336
rect 268344 162324 268350 162376
rect 374822 162324 374828 162376
rect 374880 162364 374886 162376
rect 443454 162364 443460 162376
rect 374880 162336 443460 162364
rect 374880 162324 374886 162336
rect 443454 162324 443460 162336
rect 443512 162324 443518 162376
rect 54938 162256 54944 162308
rect 54996 162296 55002 162308
rect 113542 162296 113548 162308
rect 54996 162268 113548 162296
rect 54996 162256 55002 162268
rect 113542 162256 113548 162268
rect 113600 162256 113606 162308
rect 183462 162256 183468 162308
rect 183520 162296 183526 162308
rect 197354 162296 197360 162308
rect 183520 162268 197360 162296
rect 183520 162256 183526 162268
rect 197354 162256 197360 162268
rect 197412 162256 197418 162308
rect 218974 162256 218980 162308
rect 219032 162296 219038 162308
rect 280798 162296 280804 162308
rect 219032 162268 280804 162296
rect 219032 162256 219038 162268
rect 280798 162256 280804 162268
rect 280856 162256 280862 162308
rect 343450 162256 343456 162308
rect 343508 162296 343514 162308
rect 356698 162296 356704 162308
rect 343508 162268 356704 162296
rect 343508 162256 343514 162268
rect 356698 162256 356704 162268
rect 356756 162256 356762 162308
rect 366542 162256 366548 162308
rect 366600 162296 366606 162308
rect 433518 162296 433524 162308
rect 366600 162268 433524 162296
rect 366600 162256 366606 162268
rect 433518 162256 433524 162268
rect 433576 162256 433582 162308
rect 503254 162256 503260 162308
rect 503312 162296 503318 162308
rect 517606 162296 517612 162308
rect 503312 162268 517612 162296
rect 503312 162256 503318 162268
rect 517606 162256 517612 162268
rect 517664 162256 517670 162308
rect 53558 162188 53564 162240
rect 53616 162228 53622 162240
rect 110966 162228 110972 162240
rect 53616 162200 110972 162228
rect 53616 162188 53622 162200
rect 110966 162188 110972 162200
rect 111024 162188 111030 162240
rect 216030 162188 216036 162240
rect 216088 162228 216094 162240
rect 273438 162228 273444 162240
rect 216088 162200 273444 162228
rect 216088 162188 216094 162200
rect 273438 162188 273444 162200
rect 273496 162188 273502 162240
rect 370590 162188 370596 162240
rect 370648 162228 370654 162240
rect 435910 162228 435916 162240
rect 370648 162200 435916 162228
rect 370648 162188 370654 162200
rect 435910 162188 435916 162200
rect 435968 162188 435974 162240
rect 48222 162120 48228 162172
rect 48280 162160 48286 162172
rect 93670 162160 93676 162172
rect 48280 162132 93676 162160
rect 48280 162120 48286 162132
rect 93670 162120 93676 162132
rect 93728 162120 93734 162172
rect 183186 162120 183192 162172
rect 183244 162160 183250 162172
rect 197446 162160 197452 162172
rect 183244 162132 197452 162160
rect 183244 162120 183250 162132
rect 197446 162120 197452 162132
rect 197504 162120 197510 162172
rect 210418 162120 210424 162172
rect 210476 162160 210482 162172
rect 265434 162160 265440 162172
rect 210476 162132 265440 162160
rect 210476 162120 210482 162132
rect 265434 162120 265440 162132
rect 265492 162120 265498 162172
rect 343358 162120 343364 162172
rect 343416 162160 343422 162172
rect 357526 162160 357532 162172
rect 343416 162132 357532 162160
rect 343416 162120 343422 162132
rect 357526 162120 357532 162132
rect 357584 162120 357590 162172
rect 358078 162120 358084 162172
rect 358136 162160 358142 162172
rect 413646 162160 413652 162172
rect 358136 162132 413652 162160
rect 358136 162120 358142 162132
rect 413646 162120 413652 162132
rect 413704 162120 413710 162172
rect 503622 162120 503628 162172
rect 503680 162160 503686 162172
rect 517514 162160 517520 162172
rect 503680 162132 517520 162160
rect 503680 162120 503686 162132
rect 517514 162120 517520 162132
rect 517572 162120 517578 162172
rect 49326 162052 49332 162104
rect 49384 162092 49390 162104
rect 90726 162092 90732 162104
rect 49384 162064 90732 162092
rect 49384 162052 49390 162064
rect 90726 162052 90732 162064
rect 90784 162052 90790 162104
rect 202138 162052 202144 162104
rect 202196 162092 202202 162104
rect 255958 162092 255964 162104
rect 202196 162064 255964 162092
rect 202196 162052 202202 162064
rect 255958 162052 255964 162064
rect 256016 162052 256022 162104
rect 358262 162052 358268 162104
rect 358320 162092 358326 162104
rect 408310 162092 408316 162104
rect 358320 162064 408316 162092
rect 358320 162052 358326 162064
rect 408310 162052 408316 162064
rect 408368 162052 408374 162104
rect 56502 161984 56508 162036
rect 56560 162024 56566 162036
rect 88334 162024 88340 162036
rect 56560 161996 88340 162024
rect 56560 161984 56566 161996
rect 88334 161984 88340 161996
rect 88392 161984 88398 162036
rect 213270 161984 213276 162036
rect 213328 162024 213334 162036
rect 263686 162024 263692 162036
rect 213328 161996 263692 162024
rect 213328 161984 213334 161996
rect 263686 161984 263692 161996
rect 263744 161984 263750 162036
rect 378778 161984 378784 162036
rect 378836 162024 378842 162036
rect 418430 162024 418436 162036
rect 378836 161996 418436 162024
rect 378836 161984 378842 161996
rect 418430 161984 418436 161996
rect 418488 161984 418494 162036
rect 218790 161916 218796 161968
rect 218848 161956 218854 161968
rect 247862 161956 247868 161968
rect 218848 161928 247868 161956
rect 218848 161916 218854 161928
rect 247862 161916 247868 161928
rect 247920 161916 247926 161968
rect 376294 161916 376300 161968
rect 376352 161956 376358 161968
rect 410610 161956 410616 161968
rect 376352 161928 410616 161956
rect 376352 161916 376358 161928
rect 410610 161916 410616 161928
rect 410668 161916 410674 161968
rect 360930 161848 360936 161900
rect 360988 161888 360994 161900
rect 453206 161888 453212 161900
rect 360988 161860 453212 161888
rect 360988 161848 360994 161860
rect 453206 161848 453212 161860
rect 453264 161848 453270 161900
rect 421558 161576 421564 161628
rect 421616 161616 421622 161628
rect 439038 161616 439044 161628
rect 421616 161588 439044 161616
rect 421616 161576 421622 161588
rect 439038 161576 439044 161588
rect 439096 161576 439102 161628
rect 435358 161548 435364 161560
rect 429120 161520 435364 161548
rect 87598 161440 87604 161492
rect 87656 161480 87662 161492
rect 96890 161480 96896 161492
rect 87656 161452 96896 161480
rect 87656 161440 87662 161452
rect 96890 161440 96896 161452
rect 96948 161440 96954 161492
rect 55950 161372 55956 161424
rect 56008 161412 56014 161424
rect 117314 161412 117320 161424
rect 56008 161384 117320 161412
rect 56008 161372 56014 161384
rect 117314 161372 117320 161384
rect 117372 161372 117378 161424
rect 219526 161372 219532 161424
rect 219584 161412 219590 161424
rect 267734 161412 267740 161424
rect 219584 161384 267740 161412
rect 219584 161372 219590 161384
rect 267734 161372 267740 161384
rect 267792 161372 267798 161424
rect 372246 161372 372252 161424
rect 372304 161412 372310 161424
rect 429120 161412 429148 161520
rect 435358 161508 435364 161520
rect 435416 161508 435422 161560
rect 434714 161480 434720 161492
rect 434686 161440 434720 161480
rect 434772 161440 434778 161492
rect 434686 161424 434714 161440
rect 372304 161384 429148 161412
rect 372304 161372 372310 161384
rect 434622 161372 434628 161424
rect 434680 161384 434714 161424
rect 434680 161372 434686 161384
rect 54662 161304 54668 161356
rect 54720 161344 54726 161356
rect 114738 161344 114744 161356
rect 54720 161316 114744 161344
rect 54720 161304 54726 161316
rect 114738 161304 114744 161316
rect 114796 161304 114802 161356
rect 216030 161304 216036 161356
rect 216088 161344 216094 161356
rect 263594 161344 263600 161356
rect 216088 161316 263600 161344
rect 216088 161304 216094 161316
rect 263594 161304 263600 161316
rect 263652 161304 263658 161356
rect 379514 161304 379520 161356
rect 379572 161344 379578 161356
rect 426434 161344 426440 161356
rect 379572 161316 426440 161344
rect 379572 161304 379578 161316
rect 426434 161304 426440 161316
rect 426492 161304 426498 161356
rect 59170 161236 59176 161288
rect 59228 161276 59234 161288
rect 106366 161276 106372 161288
rect 59228 161248 106372 161276
rect 59228 161236 59234 161248
rect 106366 161236 106372 161248
rect 106424 161236 106430 161288
rect 219802 161236 219808 161288
rect 219860 161276 219866 161288
rect 266354 161276 266360 161288
rect 219860 161248 266360 161276
rect 219860 161236 219866 161248
rect 266354 161236 266360 161248
rect 266412 161236 266418 161288
rect 379330 161236 379336 161288
rect 379388 161276 379394 161288
rect 422294 161276 422300 161288
rect 379388 161248 422300 161276
rect 379388 161236 379394 161248
rect 422294 161236 422300 161248
rect 422352 161236 422358 161288
rect 59722 161168 59728 161220
rect 59780 161208 59786 161220
rect 106274 161208 106280 161220
rect 59780 161180 106280 161208
rect 59780 161168 59786 161180
rect 106274 161168 106280 161180
rect 106332 161168 106338 161220
rect 219618 161168 219624 161220
rect 219676 161208 219682 161220
rect 264974 161208 264980 161220
rect 219676 161180 264980 161208
rect 219676 161168 219682 161180
rect 264974 161168 264980 161180
rect 265032 161168 265038 161220
rect 59078 161100 59084 161152
rect 59136 161140 59142 161152
rect 59136 161112 64874 161140
rect 59136 161100 59142 161112
rect 53006 161032 53012 161084
rect 53064 161072 53070 161084
rect 56502 161072 56508 161084
rect 53064 161044 56508 161072
rect 53064 161032 53070 161044
rect 56502 161032 56508 161044
rect 56560 161072 56566 161084
rect 64846 161072 64874 161112
rect 219342 161100 219348 161152
rect 219400 161140 219406 161152
rect 260834 161140 260840 161152
rect 219400 161112 260840 161140
rect 219400 161100 219406 161112
rect 260834 161100 260840 161112
rect 260892 161100 260898 161152
rect 95234 161072 95240 161084
rect 56560 161044 59308 161072
rect 64846 161044 95240 161072
rect 56560 161032 56566 161044
rect 58526 160964 58532 161016
rect 58584 161004 58590 161016
rect 59170 161004 59176 161016
rect 58584 160976 59176 161004
rect 58584 160964 58590 160976
rect 59170 160964 59176 160976
rect 59228 160964 59234 161016
rect 59280 161004 59308 161044
rect 95234 161032 95240 161044
rect 95292 161032 95298 161084
rect 217778 161032 217784 161084
rect 217836 161072 217842 161084
rect 258074 161072 258080 161084
rect 217836 161044 258080 161072
rect 217836 161032 217842 161044
rect 258074 161032 258080 161044
rect 258132 161032 258138 161084
rect 97994 161004 98000 161016
rect 59280 160976 98000 161004
rect 97994 160964 98000 160976
rect 98052 160964 98058 161016
rect 47394 160896 47400 160948
rect 47452 160936 47458 160948
rect 53466 160936 53472 160948
rect 47452 160908 53472 160936
rect 47452 160896 47458 160908
rect 53466 160896 53472 160908
rect 53524 160936 53530 160948
rect 109034 160936 109040 160948
rect 53524 160908 109040 160936
rect 53524 160896 53530 160908
rect 109034 160896 109040 160908
rect 109092 160896 109098 160948
rect 47302 160828 47308 160880
rect 47360 160868 47366 160880
rect 52086 160868 52092 160880
rect 47360 160840 52092 160868
rect 47360 160828 47366 160840
rect 52086 160828 52092 160840
rect 52144 160868 52150 160880
rect 110414 160868 110420 160880
rect 52144 160840 110420 160868
rect 52144 160828 52150 160840
rect 110414 160828 110420 160840
rect 110472 160828 110478 160880
rect 211522 160828 211528 160880
rect 211580 160868 211586 160880
rect 213362 160868 213368 160880
rect 211580 160840 213368 160868
rect 211580 160828 211586 160840
rect 213362 160828 213368 160840
rect 213420 160828 213426 160880
rect 52362 160760 52368 160812
rect 52420 160800 52426 160812
rect 59078 160800 59084 160812
rect 52420 160772 59084 160800
rect 52420 160760 52426 160772
rect 59078 160760 59084 160772
rect 59136 160760 59142 160812
rect 59354 160760 59360 160812
rect 59412 160800 59418 160812
rect 118694 160800 118700 160812
rect 59412 160772 118700 160800
rect 59412 160760 59418 160772
rect 118694 160760 118700 160772
rect 118752 160760 118758 160812
rect 262214 160800 262220 160812
rect 216140 160772 262220 160800
rect 216140 160744 216168 160772
rect 262214 160760 262220 160772
rect 262272 160760 262278 160812
rect 373442 160760 373448 160812
rect 373500 160800 373506 160812
rect 376294 160800 376300 160812
rect 373500 160772 376300 160800
rect 373500 160760 373506 160772
rect 376294 160760 376300 160772
rect 376352 160800 376358 160812
rect 429286 160800 429292 160812
rect 376352 160772 429292 160800
rect 376352 160760 376358 160772
rect 429286 160760 429292 160772
rect 429344 160760 429350 160812
rect 47486 160692 47492 160744
rect 47544 160732 47550 160744
rect 52178 160732 52184 160744
rect 47544 160704 52184 160732
rect 47544 160692 47550 160704
rect 52178 160692 52184 160704
rect 52236 160732 52242 160744
rect 111794 160732 111800 160744
rect 52236 160704 111800 160732
rect 52236 160692 52242 160704
rect 111794 160692 111800 160704
rect 111852 160692 111858 160744
rect 214650 160692 214656 160744
rect 214708 160732 214714 160744
rect 216122 160732 216128 160744
rect 214708 160704 216128 160732
rect 214708 160692 214714 160704
rect 216122 160692 216128 160704
rect 216180 160692 216186 160744
rect 273254 160732 273260 160744
rect 219406 160704 273260 160732
rect 213362 160624 213368 160676
rect 213420 160664 213426 160676
rect 219406 160664 219434 160704
rect 273254 160692 273260 160704
rect 273312 160692 273318 160744
rect 373534 160692 373540 160744
rect 373592 160732 373598 160744
rect 374822 160732 374828 160744
rect 373592 160704 374828 160732
rect 373592 160692 373598 160704
rect 374822 160692 374828 160704
rect 374880 160732 374886 160744
rect 430574 160732 430580 160744
rect 374880 160704 430580 160732
rect 374880 160692 374886 160704
rect 430574 160692 430580 160704
rect 430632 160692 430638 160744
rect 213420 160636 219434 160664
rect 213420 160624 213426 160636
rect 59722 160284 59728 160336
rect 59780 160324 59786 160336
rect 59998 160324 60004 160336
rect 59780 160296 60004 160324
rect 59780 160284 59786 160296
rect 59998 160284 60004 160296
rect 60056 160284 60062 160336
rect 53558 160080 53564 160132
rect 53616 160120 53622 160132
rect 54662 160120 54668 160132
rect 53616 160092 54668 160120
rect 53616 160080 53622 160092
rect 54662 160080 54668 160092
rect 54720 160080 54726 160132
rect 58434 160080 58440 160132
rect 58492 160120 58498 160132
rect 59354 160120 59360 160132
rect 58492 160092 59360 160120
rect 58492 160080 58498 160092
rect 59354 160080 59360 160092
rect 59412 160080 59418 160132
rect 218422 160080 218428 160132
rect 218480 160120 218486 160132
rect 219342 160120 219348 160132
rect 218480 160092 219348 160120
rect 218480 160080 218486 160092
rect 219342 160080 219348 160092
rect 219400 160080 219406 160132
rect 379514 160080 379520 160132
rect 379572 160120 379578 160132
rect 379882 160120 379888 160132
rect 379572 160092 379888 160120
rect 379572 160080 379578 160092
rect 379882 160080 379888 160092
rect 379940 160080 379946 160132
rect 215754 160012 215760 160064
rect 215812 160052 215818 160064
rect 259454 160052 259460 160064
rect 215812 160024 259460 160052
rect 215812 160012 215818 160024
rect 259454 160012 259460 160024
rect 259512 160012 259518 160064
rect 376662 160012 376668 160064
rect 376720 160052 376726 160064
rect 420914 160052 420920 160064
rect 376720 160024 420920 160052
rect 376720 160012 376726 160024
rect 420914 160012 420920 160024
rect 420972 160012 420978 160064
rect 215662 159944 215668 159996
rect 215720 159984 215726 159996
rect 259546 159984 259552 159996
rect 215720 159956 259552 159984
rect 215720 159944 215726 159956
rect 259546 159944 259552 159956
rect 259604 159944 259610 159996
rect 375374 159944 375380 159996
rect 375432 159984 375438 159996
rect 419534 159984 419540 159996
rect 375432 159956 419540 159984
rect 375432 159944 375438 159956
rect 419534 159944 419540 159956
rect 419592 159944 419598 159996
rect 378042 159876 378048 159928
rect 378100 159916 378106 159928
rect 418154 159916 418160 159928
rect 378100 159888 418160 159916
rect 378100 159876 378106 159888
rect 418154 159876 418160 159888
rect 418212 159876 418218 159928
rect 214742 159332 214748 159384
rect 214800 159372 214806 159384
rect 218882 159372 218888 159384
rect 214800 159344 218888 159372
rect 214800 159332 214806 159344
rect 218882 159332 218888 159344
rect 218940 159372 218946 159384
rect 256694 159372 256700 159384
rect 218940 159344 256700 159372
rect 218940 159332 218946 159344
rect 256694 159332 256700 159344
rect 256752 159332 256758 159384
rect 215754 159196 215760 159248
rect 215812 159236 215818 159248
rect 216398 159236 216404 159248
rect 215812 159208 216404 159236
rect 215812 159196 215818 159208
rect 216398 159196 216404 159208
rect 216456 159196 216462 159248
rect 215202 158720 215208 158772
rect 215260 158760 215266 158772
rect 215662 158760 215668 158772
rect 215260 158732 215668 158760
rect 215260 158720 215266 158732
rect 215662 158720 215668 158732
rect 215720 158720 215726 158772
rect 377122 156612 377128 156664
rect 377180 156652 377186 156664
rect 378042 156652 378048 156664
rect 377180 156624 378048 156652
rect 377180 156612 377186 156624
rect 378042 156612 378048 156624
rect 378100 156612 378106 156664
rect 53006 148996 53012 149048
rect 53064 149036 53070 149048
rect 53190 149036 53196 149048
rect 53064 149008 53196 149036
rect 53064 148996 53070 149008
rect 53190 148996 53196 149008
rect 53248 149036 53254 149048
rect 114554 149036 114560 149048
rect 53248 149008 114560 149036
rect 53248 148996 53254 149008
rect 114554 148996 114560 149008
rect 114612 148996 114618 149048
rect 213546 148996 213552 149048
rect 213604 149036 213610 149048
rect 276106 149036 276112 149048
rect 213604 149008 276112 149036
rect 213604 148996 213610 149008
rect 276106 148996 276112 149008
rect 276164 148996 276170 149048
rect 374270 148996 374276 149048
rect 374328 149036 374334 149048
rect 434714 149036 434720 149048
rect 374328 149008 434720 149036
rect 374328 148996 374334 149008
rect 434714 148996 434720 149008
rect 434772 148996 434778 149048
rect 214834 148928 214840 148980
rect 214892 148968 214898 148980
rect 274726 148968 274732 148980
rect 214892 148940 274732 148968
rect 214892 148928 214898 148940
rect 274726 148928 274732 148940
rect 274784 148928 274790 148980
rect 372338 148928 372344 148980
rect 372396 148968 372402 148980
rect 401594 148968 401600 148980
rect 372396 148940 401600 148968
rect 372396 148928 372402 148940
rect 401594 148928 401600 148940
rect 401652 148928 401658 148980
rect 212166 148860 212172 148912
rect 212224 148900 212230 148912
rect 241514 148900 241520 148912
rect 212224 148872 241520 148900
rect 212224 148860 212230 148872
rect 241514 148860 241520 148872
rect 241572 148860 241578 148912
rect 372154 148860 372160 148912
rect 372212 148900 372218 148912
rect 373626 148900 373632 148912
rect 372212 148872 373632 148900
rect 372212 148860 372218 148872
rect 373626 148860 373632 148872
rect 373684 148900 373690 148912
rect 400214 148900 400220 148912
rect 373684 148872 400220 148900
rect 373684 148860 373690 148872
rect 400214 148860 400220 148872
rect 400272 148860 400278 148912
rect 213270 148792 213276 148844
rect 213328 148832 213334 148844
rect 240134 148832 240140 148844
rect 213328 148804 240140 148832
rect 213328 148792 213334 148804
rect 240134 148792 240140 148804
rect 240192 148792 240198 148844
rect 49050 148588 49056 148640
rect 49108 148628 49114 148640
rect 54938 148628 54944 148640
rect 49108 148600 54944 148628
rect 49108 148588 49114 148600
rect 54938 148588 54944 148600
rect 54996 148628 55002 148640
rect 81434 148628 81440 148640
rect 54996 148600 81440 148628
rect 54996 148588 55002 148600
rect 81434 148588 81440 148600
rect 81492 148588 81498 148640
rect 47762 148520 47768 148572
rect 47820 148560 47826 148572
rect 53374 148560 53380 148572
rect 47820 148532 53380 148560
rect 47820 148520 47826 148532
rect 53374 148520 53380 148532
rect 53432 148560 53438 148572
rect 80054 148560 80060 148572
rect 53432 148532 80060 148560
rect 53432 148520 53438 148532
rect 80054 148520 80060 148532
rect 80112 148520 80118 148572
rect 46474 148452 46480 148504
rect 46532 148492 46538 148504
rect 51902 148492 51908 148504
rect 46532 148464 51908 148492
rect 46532 148452 46538 148464
rect 51902 148452 51908 148464
rect 51960 148492 51966 148504
rect 78674 148492 78680 148504
rect 51960 148464 78680 148492
rect 51960 148452 51966 148464
rect 78674 148452 78680 148464
rect 78732 148452 78738 148504
rect 212902 148452 212908 148504
rect 212960 148492 212966 148504
rect 213546 148492 213552 148504
rect 212960 148464 213552 148492
rect 212960 148452 212966 148464
rect 213546 148452 213552 148464
rect 213604 148452 213610 148504
rect 372522 148452 372528 148504
rect 372580 148492 372586 148504
rect 374730 148492 374736 148504
rect 372580 148464 374736 148492
rect 372580 148452 372586 148464
rect 374730 148452 374736 148464
rect 374788 148492 374794 148504
rect 397454 148492 397460 148504
rect 374788 148464 397460 148492
rect 374788 148452 374794 148464
rect 397454 148452 397460 148464
rect 397512 148452 397518 148504
rect 56226 148384 56232 148436
rect 56284 148424 56290 148436
rect 116210 148424 116216 148436
rect 56284 148396 116216 148424
rect 56284 148384 56290 148396
rect 116210 148384 116216 148396
rect 116268 148384 116274 148436
rect 376570 148384 376576 148436
rect 376628 148424 376634 148436
rect 398834 148424 398840 148436
rect 376628 148396 398840 148424
rect 376628 148384 376634 148396
rect 398834 148384 398840 148396
rect 398892 148384 398898 148436
rect 53282 148316 53288 148368
rect 53340 148356 53346 148368
rect 114646 148356 114652 148368
rect 53340 148328 114652 148356
rect 53340 148316 53346 148328
rect 114646 148316 114652 148328
rect 114704 148316 114710 148368
rect 215846 148316 215852 148368
rect 215904 148356 215910 148368
rect 238754 148356 238760 148368
rect 215904 148328 238760 148356
rect 215904 148316 215910 148328
rect 238754 148316 238760 148328
rect 238812 148316 238818 148368
rect 371786 148316 371792 148368
rect 371844 148356 371850 148368
rect 379974 148356 379980 148368
rect 371844 148328 379980 148356
rect 371844 148316 371850 148328
rect 379974 148316 379980 148328
rect 380032 148356 380038 148368
rect 429194 148356 429200 148368
rect 380032 148328 429200 148356
rect 380032 148316 380038 148328
rect 429194 148316 429200 148328
rect 429252 148316 429258 148368
rect 374270 148180 374276 148232
rect 374328 148220 374334 148232
rect 375006 148220 375012 148232
rect 374328 148192 375012 148220
rect 374328 148180 374334 148192
rect 375006 148180 375012 148192
rect 375064 148180 375070 148232
rect 57790 147568 57796 147620
rect 57848 147608 57854 147620
rect 104894 147608 104900 147620
rect 57848 147580 104900 147608
rect 57848 147568 57854 147580
rect 104894 147568 104900 147580
rect 104952 147568 104958 147620
rect 212074 147568 212080 147620
rect 212132 147608 212138 147620
rect 215846 147608 215852 147620
rect 212132 147580 215852 147608
rect 212132 147568 212138 147580
rect 215846 147568 215852 147580
rect 215904 147568 215910 147620
rect 370958 147568 370964 147620
rect 371016 147608 371022 147620
rect 376018 147608 376024 147620
rect 371016 147580 376024 147608
rect 371016 147568 371022 147580
rect 376018 147568 376024 147580
rect 376076 147608 376082 147620
rect 376570 147608 376576 147620
rect 376076 147580 376576 147608
rect 376076 147568 376082 147580
rect 376570 147568 376576 147580
rect 376628 147568 376634 147620
rect 378962 147568 378968 147620
rect 379020 147608 379026 147620
rect 379422 147608 379428 147620
rect 379020 147580 379428 147608
rect 379020 147568 379026 147580
rect 379422 147568 379428 147580
rect 379480 147608 379486 147620
rect 426526 147608 426532 147620
rect 379480 147580 426532 147608
rect 379480 147568 379486 147580
rect 426526 147568 426532 147580
rect 426584 147568 426590 147620
rect 58618 147500 58624 147552
rect 58676 147540 58682 147552
rect 103514 147540 103520 147552
rect 58676 147512 103520 147540
rect 58676 147500 58682 147512
rect 103514 147500 103520 147512
rect 103572 147500 103578 147552
rect 56134 147160 56140 147212
rect 56192 147200 56198 147212
rect 58618 147200 58624 147212
rect 56192 147172 58624 147200
rect 56192 147160 56198 147172
rect 58618 147160 58624 147172
rect 58676 147160 58682 147212
rect 59906 146888 59912 146940
rect 59964 146928 59970 146940
rect 107654 146928 107660 146940
rect 59964 146900 107660 146928
rect 59964 146888 59970 146900
rect 107654 146888 107660 146900
rect 107712 146888 107718 146940
rect 54202 146208 54208 146260
rect 54260 146248 54266 146260
rect 58802 146248 58808 146260
rect 54260 146220 58808 146248
rect 54260 146208 54266 146220
rect 58802 146208 58808 146220
rect 58860 146248 58866 146260
rect 99374 146248 99380 146260
rect 58860 146220 99380 146248
rect 58860 146208 58866 146220
rect 99374 146208 99380 146220
rect 99432 146208 99438 146260
rect 179046 146208 179052 146260
rect 179104 146248 179110 146260
rect 197538 146248 197544 146260
rect 179104 146220 197544 146248
rect 179104 146208 179110 146220
rect 197538 146208 197544 146220
rect 197596 146208 197602 146260
rect 217134 146208 217140 146260
rect 217192 146248 217198 146260
rect 255406 146248 255412 146260
rect 217192 146220 255412 146248
rect 217192 146208 217198 146220
rect 255406 146208 255412 146220
rect 255464 146208 255470 146260
rect 276014 146208 276020 146260
rect 276072 146248 276078 146260
rect 356606 146248 356612 146260
rect 276072 146220 356612 146248
rect 276072 146208 276078 146220
rect 356606 146208 356612 146220
rect 356664 146208 356670 146260
rect 358722 146208 358728 146260
rect 358780 146248 358786 146260
rect 510614 146248 510620 146260
rect 358780 146220 510620 146248
rect 358780 146208 358786 146220
rect 510614 146208 510620 146220
rect 510672 146208 510678 146260
rect 56962 146140 56968 146192
rect 57020 146180 57026 146192
rect 57238 146180 57244 146192
rect 57020 146152 57244 146180
rect 57020 146140 57026 146152
rect 57238 146140 57244 146152
rect 57296 146140 57302 146192
rect 59814 146140 59820 146192
rect 59872 146180 59878 146192
rect 93854 146180 93860 146192
rect 59872 146152 93860 146180
rect 59872 146140 59878 146152
rect 93854 146140 93860 146152
rect 93912 146140 93918 146192
rect 179690 146140 179696 146192
rect 179748 146180 179754 146192
rect 197630 146180 197636 146192
rect 179748 146152 197636 146180
rect 179748 146140 179754 146152
rect 197630 146140 197636 146152
rect 197688 146140 197694 146192
rect 219894 146140 219900 146192
rect 219952 146180 219958 146192
rect 253934 146180 253940 146192
rect 219952 146152 253940 146180
rect 219952 146140 219958 146152
rect 253934 146140 253940 146152
rect 253992 146140 253998 146192
rect 338482 146140 338488 146192
rect 338540 146180 338546 146192
rect 356882 146180 356888 146192
rect 338540 146152 356888 146180
rect 338540 146140 338546 146152
rect 356882 146140 356888 146152
rect 356940 146140 356946 146192
rect 374546 146140 374552 146192
rect 374604 146180 374610 146192
rect 375650 146180 375656 146192
rect 374604 146152 375656 146180
rect 374604 146140 374610 146152
rect 375650 146140 375656 146152
rect 375708 146140 375714 146192
rect 377214 146140 377220 146192
rect 377272 146180 377278 146192
rect 377950 146180 377956 146192
rect 377272 146152 377956 146180
rect 377272 146140 377278 146152
rect 377950 146140 377956 146152
rect 378008 146140 378014 146192
rect 378594 146140 378600 146192
rect 378652 146180 378658 146192
rect 378962 146180 378968 146192
rect 378652 146152 378968 146180
rect 378652 146140 378658 146152
rect 378962 146140 378968 146152
rect 379020 146140 379026 146192
rect 379606 146140 379612 146192
rect 379664 146180 379670 146192
rect 379790 146180 379796 146192
rect 379664 146152 379796 146180
rect 379664 146140 379670 146152
rect 379790 146140 379796 146152
rect 379848 146180 379854 146192
rect 414014 146180 414020 146192
rect 379848 146152 414020 146180
rect 379848 146140 379854 146152
rect 414014 146140 414020 146152
rect 414072 146140 414078 146192
rect 498654 146140 498660 146192
rect 498712 146180 498718 146192
rect 517790 146180 517796 146192
rect 498712 146152 517796 146180
rect 498712 146140 498718 146152
rect 517790 146140 517796 146152
rect 517848 146180 517854 146192
rect 518066 146180 518072 146192
rect 517848 146152 518072 146180
rect 517848 146140 517854 146152
rect 518066 146140 518072 146152
rect 518124 146140 518130 146192
rect 57256 146112 57284 146140
rect 91186 146112 91192 146124
rect 57256 146084 91192 146112
rect 91186 146072 91192 146084
rect 91244 146072 91250 146124
rect 218790 146072 218796 146124
rect 218848 146112 218854 146124
rect 219158 146112 219164 146124
rect 218848 146084 219164 146112
rect 218848 146072 218854 146084
rect 219158 146072 219164 146084
rect 219216 146112 219222 146124
rect 252554 146112 252560 146124
rect 219216 146084 252560 146112
rect 219216 146072 219222 146084
rect 252554 146072 252560 146084
rect 252612 146072 252618 146124
rect 340230 146072 340236 146124
rect 340288 146112 340294 146124
rect 357434 146112 357440 146124
rect 340288 146084 357440 146112
rect 340288 146072 340294 146084
rect 357434 146072 357440 146084
rect 357492 146072 357498 146124
rect 374454 146072 374460 146124
rect 374512 146112 374518 146124
rect 375098 146112 375104 146124
rect 374512 146084 375104 146112
rect 374512 146072 374518 146084
rect 375098 146072 375104 146084
rect 375156 146072 375162 146124
rect 53190 146004 53196 146056
rect 53248 146044 53254 146056
rect 53834 146044 53840 146056
rect 53248 146016 53840 146044
rect 53248 146004 53254 146016
rect 53834 146004 53840 146016
rect 53892 146044 53898 146056
rect 86954 146044 86960 146056
rect 53892 146016 86960 146044
rect 53892 146004 53898 146016
rect 86954 146004 86960 146016
rect 87012 146004 87018 146056
rect 216766 146004 216772 146056
rect 216824 146044 216830 146056
rect 251174 146044 251180 146056
rect 216824 146016 251180 146044
rect 216824 146004 216830 146016
rect 56042 145936 56048 145988
rect 56100 145976 56106 145988
rect 88426 145976 88432 145988
rect 56100 145948 88432 145976
rect 56100 145936 56106 145948
rect 88426 145936 88432 145948
rect 88484 145936 88490 145988
rect 54570 145868 54576 145920
rect 54628 145908 54634 145920
rect 54846 145908 54852 145920
rect 54628 145880 54852 145908
rect 54628 145868 54634 145880
rect 54846 145868 54852 145880
rect 54904 145908 54910 145920
rect 85574 145908 85580 145920
rect 54904 145880 85580 145908
rect 54904 145868 54910 145880
rect 85574 145868 85580 145880
rect 85632 145868 85638 145920
rect 58894 145800 58900 145852
rect 58952 145840 58958 145852
rect 89806 145840 89812 145852
rect 58952 145812 89812 145840
rect 58952 145800 58958 145812
rect 89806 145800 89812 145812
rect 89864 145800 89870 145852
rect 47578 145732 47584 145784
rect 47636 145772 47642 145784
rect 52362 145772 52368 145784
rect 47636 145744 52368 145772
rect 47636 145732 47642 145744
rect 52362 145732 52368 145744
rect 52420 145772 52426 145784
rect 77294 145772 77300 145784
rect 52420 145744 77300 145772
rect 52420 145732 52426 145744
rect 77294 145732 77300 145744
rect 77352 145732 77358 145784
rect 217796 145772 217824 146016
rect 251174 146004 251180 146016
rect 251232 146004 251238 146056
rect 377968 146044 377996 146140
rect 396718 146072 396724 146124
rect 396776 146112 396782 146124
rect 416774 146112 416780 146124
rect 396776 146084 416780 146112
rect 396776 146072 396782 146084
rect 416774 146072 416780 146084
rect 416832 146072 416838 146124
rect 499850 146072 499856 146124
rect 499908 146112 499914 146124
rect 517882 146112 517888 146124
rect 499908 146084 517888 146112
rect 499908 146072 499914 146084
rect 517882 146072 517888 146084
rect 517940 146112 517946 146124
rect 518434 146112 518440 146124
rect 517940 146084 518440 146112
rect 517940 146072 517946 146084
rect 518434 146072 518440 146084
rect 518492 146072 518498 146124
rect 409966 146044 409972 146056
rect 377968 146016 409972 146044
rect 409966 146004 409972 146016
rect 410024 146004 410030 146056
rect 219066 145936 219072 145988
rect 219124 145976 219130 145988
rect 251266 145976 251272 145988
rect 219124 145948 251272 145976
rect 219124 145936 219130 145948
rect 251266 145936 251272 145948
rect 251324 145936 251330 145988
rect 374362 145936 374368 145988
rect 374420 145976 374426 145988
rect 378686 145976 378692 145988
rect 374420 145948 378692 145976
rect 374420 145936 374426 145948
rect 378686 145936 378692 145948
rect 378744 145936 378750 145988
rect 379238 145936 379244 145988
rect 379296 145976 379302 145988
rect 411346 145976 411352 145988
rect 379296 145948 411352 145976
rect 379296 145936 379302 145948
rect 411346 145936 411352 145948
rect 411404 145936 411410 145988
rect 217870 145868 217876 145920
rect 217928 145908 217934 145920
rect 249794 145908 249800 145920
rect 217928 145880 249800 145908
rect 217928 145868 217934 145880
rect 249794 145868 249800 145880
rect 249852 145868 249858 145920
rect 375742 145868 375748 145920
rect 375800 145908 375806 145920
rect 407206 145908 407212 145920
rect 375800 145880 407212 145908
rect 375800 145868 375806 145880
rect 407206 145868 407212 145880
rect 407264 145868 407270 145920
rect 219406 145812 224264 145840
rect 217870 145772 217876 145784
rect 217796 145744 217876 145772
rect 217870 145732 217876 145744
rect 217928 145732 217934 145784
rect 218606 145732 218612 145784
rect 218664 145772 218670 145784
rect 219250 145772 219256 145784
rect 218664 145744 219256 145772
rect 218664 145732 218670 145744
rect 219250 145732 219256 145744
rect 219308 145772 219314 145784
rect 219406 145772 219434 145812
rect 219308 145744 219434 145772
rect 224236 145772 224264 145812
rect 224310 145800 224316 145852
rect 224368 145840 224374 145852
rect 247126 145840 247132 145852
rect 224368 145812 247132 145840
rect 224368 145800 224374 145812
rect 247126 145800 247132 145812
rect 247184 145800 247190 145852
rect 375098 145800 375104 145852
rect 375156 145800 375162 145852
rect 378962 145800 378968 145852
rect 379020 145840 379026 145852
rect 408494 145840 408500 145852
rect 379020 145812 408500 145840
rect 379020 145800 379026 145812
rect 408494 145800 408500 145812
rect 408552 145800 408558 145852
rect 248414 145772 248420 145784
rect 224236 145744 248420 145772
rect 219308 145732 219314 145744
rect 248414 145732 248420 145744
rect 248472 145732 248478 145784
rect 375116 145772 375144 145800
rect 402974 145772 402980 145784
rect 375116 145744 402980 145772
rect 402974 145732 402980 145744
rect 403032 145732 403038 145784
rect 49234 145664 49240 145716
rect 49292 145704 49298 145716
rect 54662 145704 54668 145716
rect 49292 145676 54668 145704
rect 49292 145664 49298 145676
rect 54662 145664 54668 145676
rect 54720 145704 54726 145716
rect 82814 145704 82820 145716
rect 54720 145676 82820 145704
rect 54720 145664 54726 145676
rect 82814 145664 82820 145676
rect 82872 145664 82878 145716
rect 216214 145664 216220 145716
rect 216272 145704 216278 145716
rect 224126 145704 224132 145716
rect 216272 145676 224132 145704
rect 216272 145664 216278 145676
rect 224126 145664 224132 145676
rect 224184 145664 224190 145716
rect 224218 145664 224224 145716
rect 224276 145704 224282 145716
rect 244274 145704 244280 145716
rect 224276 145676 244280 145704
rect 224276 145664 224282 145676
rect 244274 145664 244280 145676
rect 244332 145664 244338 145716
rect 375650 145664 375656 145716
rect 375708 145704 375714 145716
rect 403066 145704 403072 145716
rect 375708 145676 403072 145704
rect 375708 145664 375714 145676
rect 403066 145664 403072 145676
rect 403124 145664 403130 145716
rect 56318 145596 56324 145648
rect 56376 145636 56382 145648
rect 84286 145636 84292 145648
rect 56376 145608 84292 145636
rect 56376 145596 56382 145608
rect 84286 145596 84292 145608
rect 84344 145596 84350 145648
rect 216306 145596 216312 145648
rect 216364 145636 216370 145648
rect 244366 145636 244372 145648
rect 216364 145608 244372 145636
rect 216364 145596 216370 145608
rect 244366 145596 244372 145608
rect 244424 145596 244430 145648
rect 280062 145596 280068 145648
rect 280120 145636 280126 145648
rect 356606 145636 356612 145648
rect 280120 145608 356612 145636
rect 280120 145596 280126 145608
rect 356606 145596 356612 145608
rect 356664 145636 356670 145648
rect 357618 145636 357624 145648
rect 356664 145608 357624 145636
rect 356664 145596 356670 145608
rect 357618 145596 357624 145608
rect 357676 145596 357682 145648
rect 376570 145596 376576 145648
rect 376628 145636 376634 145648
rect 404354 145636 404360 145648
rect 376628 145608 404360 145636
rect 376628 145596 376634 145608
rect 404354 145596 404360 145608
rect 404412 145596 404418 145648
rect 518434 145596 518440 145648
rect 518492 145636 518498 145648
rect 580258 145636 580264 145648
rect 518492 145608 580264 145636
rect 518492 145596 518498 145608
rect 580258 145596 580264 145608
rect 580316 145596 580322 145648
rect 58802 145528 58808 145580
rect 58860 145568 58866 145580
rect 91094 145568 91100 145580
rect 58860 145540 91100 145568
rect 58860 145528 58866 145540
rect 91094 145528 91100 145540
rect 91152 145528 91158 145580
rect 191742 145528 191748 145580
rect 191800 145568 191806 145580
rect 197998 145568 198004 145580
rect 191800 145540 198004 145568
rect 191800 145528 191806 145540
rect 197998 145528 198004 145540
rect 198056 145568 198062 145580
rect 204898 145568 204904 145580
rect 198056 145540 204904 145568
rect 198056 145528 198062 145540
rect 204898 145528 204904 145540
rect 204956 145528 204962 145580
rect 214742 145528 214748 145580
rect 214800 145568 214806 145580
rect 245654 145568 245660 145580
rect 214800 145540 245660 145568
rect 214800 145528 214806 145540
rect 245654 145528 245660 145540
rect 245712 145528 245718 145580
rect 351638 145528 351644 145580
rect 351696 145568 351702 145580
rect 358722 145568 358728 145580
rect 351696 145540 358728 145568
rect 351696 145528 351702 145540
rect 358722 145528 358728 145540
rect 358780 145528 358786 145580
rect 375190 145528 375196 145580
rect 375248 145568 375254 145580
rect 405734 145568 405740 145580
rect 375248 145540 405740 145568
rect 375248 145528 375254 145540
rect 405734 145528 405740 145540
rect 405792 145528 405798 145580
rect 518066 145528 518072 145580
rect 518124 145568 518130 145580
rect 580350 145568 580356 145580
rect 518124 145540 580356 145568
rect 518124 145528 518130 145540
rect 580350 145528 580356 145540
rect 580408 145528 580414 145580
rect 58710 145460 58716 145512
rect 58768 145500 58774 145512
rect 84194 145500 84200 145512
rect 58768 145472 84200 145500
rect 58768 145460 58774 145472
rect 84194 145460 84200 145472
rect 84252 145460 84258 145512
rect 214466 145460 214472 145512
rect 214524 145500 214530 145512
rect 242894 145500 242900 145512
rect 214524 145472 242900 145500
rect 214524 145460 214530 145472
rect 242894 145460 242900 145472
rect 242952 145460 242958 145512
rect 375742 145460 375748 145512
rect 375800 145500 375806 145512
rect 376478 145500 376484 145512
rect 375800 145472 376484 145500
rect 375800 145460 375806 145472
rect 376478 145460 376484 145472
rect 376536 145460 376542 145512
rect 378594 145460 378600 145512
rect 378652 145500 378658 145512
rect 396074 145500 396080 145512
rect 378652 145472 396080 145500
rect 378652 145460 378658 145472
rect 396074 145460 396080 145472
rect 396132 145460 396138 145512
rect 47210 145392 47216 145444
rect 47268 145432 47274 145444
rect 55030 145432 55036 145444
rect 47268 145404 55036 145432
rect 47268 145392 47274 145404
rect 55030 145392 55036 145404
rect 55088 145432 55094 145444
rect 76006 145432 76012 145444
rect 55088 145404 76012 145432
rect 55088 145392 55094 145404
rect 76006 145392 76012 145404
rect 76064 145392 76070 145444
rect 215570 145392 215576 145444
rect 215628 145432 215634 145444
rect 218514 145432 218520 145444
rect 215628 145404 218520 145432
rect 215628 145392 215634 145404
rect 218514 145392 218520 145404
rect 218572 145432 218578 145444
rect 236086 145432 236092 145444
rect 218572 145404 236092 145432
rect 218572 145392 218578 145404
rect 236086 145392 236092 145404
rect 236144 145392 236150 145444
rect 378686 145392 378692 145444
rect 378744 145432 378750 145444
rect 396166 145432 396172 145444
rect 378744 145404 396172 145432
rect 378744 145392 378750 145404
rect 396166 145392 396172 145404
rect 396224 145392 396230 145444
rect 46658 145324 46664 145376
rect 46716 145364 46722 145376
rect 54754 145364 54760 145376
rect 46716 145336 54760 145364
rect 46716 145324 46722 145336
rect 54754 145324 54760 145336
rect 54812 145364 54818 145376
rect 75914 145364 75920 145376
rect 54812 145336 75920 145364
rect 54812 145324 54818 145336
rect 75914 145324 75920 145336
rect 75972 145324 75978 145376
rect 215110 145324 215116 145376
rect 215168 145364 215174 145376
rect 219158 145364 219164 145376
rect 215168 145336 219164 145364
rect 215168 145324 215174 145336
rect 219158 145324 219164 145336
rect 219216 145364 219222 145376
rect 235994 145364 236000 145376
rect 219216 145336 236000 145364
rect 219216 145324 219222 145336
rect 235994 145324 236000 145336
rect 236052 145324 236058 145376
rect 378778 145324 378784 145376
rect 378836 145364 378842 145376
rect 393314 145364 393320 145376
rect 378836 145336 393320 145364
rect 378836 145324 378842 145336
rect 393314 145324 393320 145336
rect 393372 145324 393378 145376
rect 49142 145256 49148 145308
rect 49200 145296 49206 145308
rect 59906 145296 59912 145308
rect 49200 145268 59912 145296
rect 49200 145256 49206 145268
rect 59906 145256 59912 145268
rect 59964 145256 59970 145308
rect 377030 145256 377036 145308
rect 377088 145296 377094 145308
rect 411254 145296 411260 145308
rect 377088 145268 411260 145296
rect 377088 145256 377094 145268
rect 411254 145256 411260 145268
rect 411312 145256 411318 145308
rect 215018 145188 215024 145240
rect 215076 145228 215082 145240
rect 224218 145228 224224 145240
rect 215076 145200 224224 145228
rect 215076 145188 215082 145200
rect 224218 145188 224224 145200
rect 224276 145188 224282 145240
rect 54478 144848 54484 144900
rect 54536 144888 54542 144900
rect 55950 144888 55956 144900
rect 54536 144860 55956 144888
rect 54536 144848 54542 144860
rect 55950 144848 55956 144860
rect 56008 144888 56014 144900
rect 56318 144888 56324 144900
rect 56008 144860 56324 144888
rect 56008 144848 56014 144860
rect 56318 144848 56324 144860
rect 56376 144848 56382 144900
rect 213638 144848 213644 144900
rect 213696 144888 213702 144900
rect 214742 144888 214748 144900
rect 213696 144860 214748 144888
rect 213696 144848 213702 144860
rect 214742 144848 214748 144860
rect 214800 144848 214806 144900
rect 373166 144848 373172 144900
rect 373224 144888 373230 144900
rect 375190 144888 375196 144900
rect 373224 144860 375196 144888
rect 373224 144848 373230 144860
rect 375190 144848 375196 144860
rect 375248 144848 375254 144900
rect 377950 144848 377956 144900
rect 378008 144888 378014 144900
rect 421558 144888 421564 144900
rect 378008 144860 421564 144888
rect 378008 144848 378014 144860
rect 421558 144848 421564 144860
rect 421616 144848 421622 144900
rect 53098 144780 53104 144832
rect 53156 144820 53162 144832
rect 55858 144820 55864 144832
rect 53156 144792 55864 144820
rect 53156 144780 53162 144792
rect 55858 144780 55864 144792
rect 55916 144820 55922 144832
rect 56410 144820 56416 144832
rect 55916 144792 56416 144820
rect 55916 144780 55922 144792
rect 56410 144780 56416 144792
rect 56468 144780 56474 144832
rect 213454 144780 213460 144832
rect 213512 144820 213518 144832
rect 214650 144820 214656 144832
rect 213512 144792 214656 144820
rect 213512 144780 213518 144792
rect 214650 144780 214656 144792
rect 214708 144780 214714 144832
rect 375098 144780 375104 144832
rect 375156 144820 375162 144832
rect 378594 144820 378600 144832
rect 375156 144792 378600 144820
rect 375156 144780 375162 144792
rect 378594 144780 378600 144792
rect 378652 144780 378658 144832
rect 51994 144712 52000 144764
rect 52052 144752 52058 144764
rect 58710 144752 58716 144764
rect 52052 144724 58716 144752
rect 52052 144712 52058 144724
rect 58710 144712 58716 144724
rect 58768 144712 58774 144764
rect 212350 144712 212356 144764
rect 212408 144752 212414 144764
rect 215846 144752 215852 144764
rect 212408 144724 215852 144752
rect 212408 144712 212414 144724
rect 215846 144712 215852 144724
rect 215904 144712 215910 144764
rect 373718 144712 373724 144764
rect 373776 144752 373782 144764
rect 376202 144752 376208 144764
rect 373776 144724 376208 144752
rect 373776 144712 373782 144724
rect 376202 144712 376208 144724
rect 376260 144752 376266 144764
rect 376570 144752 376576 144764
rect 376260 144724 376576 144752
rect 376260 144712 376266 144724
rect 376570 144712 376576 144724
rect 376628 144712 376634 144764
rect 47946 144644 47952 144696
rect 48004 144684 48010 144696
rect 58618 144684 58624 144696
rect 48004 144656 58624 144684
rect 48004 144644 48010 144656
rect 58618 144644 58624 144656
rect 58676 144644 58682 144696
rect 210694 144644 210700 144696
rect 210752 144684 210758 144696
rect 214558 144684 214564 144696
rect 210752 144656 214564 144684
rect 210752 144644 210758 144656
rect 214558 144644 214564 144656
rect 214616 144644 214622 144696
rect 50338 144576 50344 144628
rect 50396 144616 50402 144628
rect 58802 144616 58808 144628
rect 50396 144588 58808 144616
rect 50396 144576 50402 144588
rect 58802 144576 58808 144588
rect 58860 144576 58866 144628
rect 56134 144508 56140 144560
rect 56192 144548 56198 144560
rect 56410 144548 56416 144560
rect 56192 144520 56416 144548
rect 56192 144508 56198 144520
rect 56410 144508 56416 144520
rect 56468 144508 56474 144560
rect 56226 144440 56232 144492
rect 56284 144440 56290 144492
rect 56244 144288 56272 144440
rect 56226 144236 56232 144288
rect 56284 144236 56290 144288
rect 520182 79976 520188 80028
rect 520240 80016 520246 80028
rect 580442 80016 580448 80028
rect 520240 79988 580448 80016
rect 520240 79976 520246 79988
rect 580442 79976 580448 79988
rect 580500 79976 580506 80028
rect 364978 70320 364984 70372
rect 365036 70360 365042 70372
rect 376938 70360 376944 70372
rect 365036 70332 376944 70360
rect 365036 70320 365042 70332
rect 376938 70320 376944 70332
rect 376996 70320 377002 70372
rect 374638 68960 374644 69012
rect 374696 69000 374702 69012
rect 377306 69000 377312 69012
rect 374696 68972 377312 69000
rect 374696 68960 374702 68972
rect 377306 68960 377312 68972
rect 377364 68960 377370 69012
rect 358722 68280 358728 68332
rect 358780 68320 358786 68332
rect 376938 68320 376944 68332
rect 358780 68292 376944 68320
rect 358780 68280 358786 68292
rect 376938 68280 376944 68292
rect 376996 68280 377002 68332
rect 358078 68144 358084 68196
rect 358136 68184 358142 68196
rect 358722 68184 358728 68196
rect 358136 68156 358728 68184
rect 358136 68144 358142 68156
rect 358722 68144 358728 68156
rect 358780 68144 358786 68196
rect 204898 67600 204904 67652
rect 204956 67640 204962 67652
rect 216674 67640 216680 67652
rect 204956 67612 216680 67640
rect 204956 67600 204962 67612
rect 216674 67600 216680 67612
rect 216732 67600 216738 67652
rect 378686 59780 378692 59832
rect 378744 59820 378750 59832
rect 397086 59820 397092 59832
rect 378744 59792 397092 59820
rect 378744 59780 378750 59792
rect 397086 59780 397092 59792
rect 397144 59780 397150 59832
rect 218514 59712 218520 59764
rect 218572 59752 218578 59764
rect 237098 59752 237104 59764
rect 218572 59724 237104 59752
rect 218572 59712 218578 59724
rect 237098 59712 237104 59724
rect 237156 59712 237162 59764
rect 378594 59712 378600 59764
rect 378652 59752 378658 59764
rect 396074 59752 396080 59764
rect 378652 59724 396080 59752
rect 378652 59712 378658 59724
rect 396074 59712 396080 59724
rect 396132 59712 396138 59764
rect 55030 59644 55036 59696
rect 55088 59684 55094 59696
rect 77110 59684 77116 59696
rect 55088 59656 77116 59684
rect 55088 59644 55094 59656
rect 77110 59644 77116 59656
rect 77168 59644 77174 59696
rect 217134 59644 217140 59696
rect 217192 59684 217198 59696
rect 255866 59684 255872 59696
rect 217192 59656 255872 59684
rect 217192 59644 217198 59656
rect 255866 59644 255872 59656
rect 255924 59644 255930 59696
rect 378042 59644 378048 59696
rect 378100 59684 378106 59696
rect 416958 59684 416964 59696
rect 378100 59656 416964 59684
rect 378100 59644 378106 59656
rect 416958 59644 416964 59656
rect 417016 59644 417022 59696
rect 54662 59576 54668 59628
rect 54720 59616 54726 59628
rect 83090 59616 83096 59628
rect 54720 59588 83096 59616
rect 54720 59576 54726 59588
rect 83090 59576 83096 59588
rect 83148 59576 83154 59628
rect 218422 59576 218428 59628
rect 218480 59616 218486 59628
rect 261754 59616 261760 59628
rect 218480 59588 261760 59616
rect 218480 59576 218486 59588
rect 261754 59576 261760 59588
rect 261812 59576 261818 59628
rect 378778 59576 378784 59628
rect 378836 59616 378842 59628
rect 418154 59616 418160 59628
rect 378836 59588 418160 59616
rect 378836 59576 378842 59588
rect 418154 59576 418160 59588
rect 418212 59576 418218 59628
rect 54202 59508 54208 59560
rect 54260 59548 54266 59560
rect 99466 59548 99472 59560
rect 54260 59520 99472 59548
rect 54260 59508 54266 59520
rect 99466 59508 99472 59520
rect 99524 59508 99530 59560
rect 216398 59508 216404 59560
rect 216456 59548 216462 59560
rect 260650 59548 260656 59560
rect 216456 59520 260656 59548
rect 216456 59508 216462 59520
rect 260650 59508 260656 59520
rect 260708 59508 260714 59560
rect 379330 59508 379336 59560
rect 379388 59548 379394 59560
rect 422846 59548 422852 59560
rect 379388 59520 422852 59548
rect 379388 59508 379394 59520
rect 422846 59508 422852 59520
rect 422904 59508 422910 59560
rect 49602 59440 49608 59492
rect 49660 59480 49666 59492
rect 113542 59480 113548 59492
rect 49660 59452 113548 59480
rect 49660 59440 49666 59452
rect 113542 59440 113548 59452
rect 113600 59440 113606 59492
rect 215202 59440 215208 59492
rect 215260 59480 215266 59492
rect 259454 59480 259460 59492
rect 215260 59452 259460 59480
rect 215260 59440 215266 59452
rect 259454 59440 259460 59452
rect 259512 59440 259518 59492
rect 375926 59440 375932 59492
rect 375984 59480 375990 59492
rect 423950 59480 423956 59492
rect 375984 59452 423956 59480
rect 375984 59440 375990 59452
rect 423950 59440 423956 59452
rect 424008 59440 424014 59492
rect 50890 59372 50896 59424
rect 50948 59412 50954 59424
rect 120902 59412 120908 59424
rect 50948 59384 120908 59412
rect 50948 59372 50954 59384
rect 120902 59372 120908 59384
rect 120960 59372 120966 59424
rect 216030 59372 216036 59424
rect 216088 59412 216094 59424
rect 263870 59412 263876 59424
rect 216088 59384 263876 59412
rect 216088 59372 216094 59384
rect 263870 59372 263876 59384
rect 263928 59372 263934 59424
rect 358170 59372 358176 59424
rect 358228 59412 358234 59424
rect 418430 59412 418436 59424
rect 358228 59384 418436 59412
rect 358228 59372 358234 59384
rect 418430 59372 418436 59384
rect 418488 59372 418494 59424
rect 55950 59304 55956 59356
rect 56008 59344 56014 59356
rect 84194 59344 84200 59356
rect 56008 59316 84200 59344
rect 56008 59304 56014 59316
rect 84194 59304 84200 59316
rect 84252 59304 84258 59356
rect 217962 59304 217968 59356
rect 218020 59344 218026 59356
rect 358078 59344 358084 59356
rect 218020 59316 358084 59344
rect 218020 59304 218026 59316
rect 358078 59304 358084 59316
rect 358136 59304 358142 59356
rect 59814 59236 59820 59288
rect 59872 59276 59878 59288
rect 94498 59276 94504 59288
rect 59872 59248 94504 59276
rect 59872 59236 59878 59248
rect 94498 59236 94504 59248
rect 94556 59236 94562 59288
rect 218882 59236 218888 59288
rect 218940 59276 218946 59288
rect 256970 59276 256976 59288
rect 218940 59248 256976 59276
rect 218940 59236 218946 59248
rect 256970 59236 256976 59248
rect 257028 59236 257034 59288
rect 374546 59236 374552 59288
rect 374604 59276 374610 59288
rect 403066 59276 403072 59288
rect 374604 59248 403072 59276
rect 374604 59236 374610 59248
rect 403066 59236 403072 59248
rect 403124 59236 403130 59288
rect 59078 59168 59084 59220
rect 59136 59208 59142 59220
rect 95878 59208 95884 59220
rect 59136 59180 95884 59208
rect 59136 59168 59142 59180
rect 95878 59168 95884 59180
rect 95936 59168 95942 59220
rect 217778 59168 217784 59220
rect 217836 59208 217842 59220
rect 258074 59208 258080 59220
rect 217836 59180 258080 59208
rect 217836 59168 217842 59180
rect 258074 59168 258080 59180
rect 258132 59168 258138 59220
rect 376662 59168 376668 59220
rect 376720 59208 376726 59220
rect 421742 59208 421748 59220
rect 376720 59180 421748 59208
rect 376720 59168 376726 59180
rect 421742 59168 421748 59180
rect 421800 59168 421806 59220
rect 56502 59100 56508 59152
rect 56560 59140 56566 59152
rect 98086 59140 98092 59152
rect 56560 59112 98092 59140
rect 56560 59100 56566 59112
rect 98086 59100 98092 59112
rect 98144 59100 98150 59152
rect 219618 59100 219624 59152
rect 219676 59140 219682 59152
rect 265250 59140 265256 59152
rect 219676 59112 265256 59140
rect 219676 59100 219682 59112
rect 265250 59100 265256 59112
rect 265308 59100 265314 59152
rect 375282 59100 375288 59152
rect 375340 59140 375346 59152
rect 420638 59140 420644 59152
rect 375340 59112 420644 59140
rect 375340 59100 375346 59112
rect 420638 59100 420644 59112
rect 420696 59100 420702 59152
rect 55858 59032 55864 59084
rect 55916 59072 55922 59084
rect 100754 59072 100760 59084
rect 55916 59044 100760 59072
rect 55916 59032 55922 59044
rect 100754 59032 100760 59044
rect 100812 59032 100818 59084
rect 216122 59032 216128 59084
rect 216180 59072 216186 59084
rect 262766 59072 262772 59084
rect 216180 59044 262772 59072
rect 216180 59032 216186 59044
rect 262766 59032 262772 59044
rect 262824 59032 262830 59084
rect 373258 59032 373264 59084
rect 373316 59072 373322 59084
rect 425974 59072 425980 59084
rect 373316 59044 425980 59072
rect 373316 59032 373322 59044
rect 425974 59032 425980 59044
rect 426032 59032 426038 59084
rect 58526 58964 58532 59016
rect 58584 59004 58590 59016
rect 102778 59004 102784 59016
rect 58584 58976 102784 59004
rect 58584 58964 58590 58976
rect 102778 58964 102784 58976
rect 102836 58964 102842 59016
rect 206922 58964 206928 59016
rect 206980 59004 206986 59016
rect 295886 59004 295892 59016
rect 206980 58976 295892 59004
rect 206980 58964 206986 58976
rect 295886 58964 295892 58976
rect 295944 58964 295950 59016
rect 362218 58964 362224 59016
rect 362276 59004 362282 59016
rect 423490 59004 423496 59016
rect 362276 58976 423496 59004
rect 362276 58964 362282 58976
rect 423490 58964 423496 58976
rect 423548 58964 423554 59016
rect 54386 58896 54392 58948
rect 54444 58936 54450 58948
rect 101766 58936 101772 58948
rect 54444 58908 101772 58936
rect 54444 58896 54450 58908
rect 101766 58896 101772 58908
rect 101824 58896 101830 58948
rect 211614 58896 211620 58948
rect 211672 58936 211678 58948
rect 303430 58936 303436 58948
rect 211672 58908 303436 58936
rect 211672 58896 211678 58908
rect 303430 58896 303436 58908
rect 303488 58896 303494 58948
rect 366358 58896 366364 58948
rect 366416 58936 366422 58948
rect 453390 58936 453396 58948
rect 366416 58908 453396 58936
rect 366416 58896 366422 58908
rect 453390 58896 453396 58908
rect 453448 58896 453454 58948
rect 56226 58828 56232 58880
rect 56284 58868 56290 58880
rect 116946 58868 116952 58880
rect 56284 58840 116952 58868
rect 56284 58828 56290 58840
rect 116946 58828 116952 58840
rect 117004 58828 117010 58880
rect 201402 58828 201408 58880
rect 201460 58868 201466 58880
rect 298462 58868 298468 58880
rect 201460 58840 298468 58868
rect 201460 58828 201466 58840
rect 298462 58828 298468 58840
rect 298520 58828 298526 58880
rect 360838 58828 360844 58880
rect 360896 58868 360902 58880
rect 463510 58868 463516 58880
rect 360896 58840 463516 58868
rect 360896 58828 360902 58840
rect 463510 58828 463516 58840
rect 463568 58828 463574 58880
rect 53006 58760 53012 58812
rect 53064 58800 53070 58812
rect 113266 58800 113272 58812
rect 53064 58772 113272 58800
rect 53064 58760 53070 58772
rect 113266 58760 113272 58772
rect 113324 58760 113330 58812
rect 198642 58760 198648 58812
rect 198700 58800 198706 58812
rect 315850 58800 315856 58812
rect 198700 58772 315856 58800
rect 198700 58760 198706 58772
rect 315850 58760 315856 58772
rect 315908 58760 315914 58812
rect 366450 58760 366456 58812
rect 366508 58800 366514 58812
rect 480898 58800 480904 58812
rect 366508 58772 480904 58800
rect 366508 58760 366514 58772
rect 480898 58760 480904 58772
rect 480956 58760 480962 58812
rect 50062 58692 50068 58744
rect 50120 58732 50126 58744
rect 148502 58732 148508 58744
rect 50120 58704 148508 58732
rect 50120 58692 50126 58704
rect 148502 58692 148508 58704
rect 148560 58692 148566 58744
rect 206830 58692 206836 58744
rect 206888 58732 206894 58744
rect 323302 58732 323308 58744
rect 206888 58704 323308 58732
rect 206888 58692 206894 58704
rect 323302 58692 323308 58704
rect 323360 58692 323366 58744
rect 361482 58692 361488 58744
rect 361540 58732 361546 58744
rect 485958 58732 485964 58744
rect 361540 58704 485964 58732
rect 361540 58692 361546 58704
rect 485958 58692 485964 58704
rect 486016 58692 486022 58744
rect 52822 58624 52828 58676
rect 52880 58664 52886 58676
rect 150894 58664 150900 58676
rect 52880 58636 150900 58664
rect 52880 58624 52886 58636
rect 150894 58624 150900 58636
rect 150952 58624 150958 58676
rect 219250 58624 219256 58676
rect 219308 58664 219314 58676
rect 428182 58664 428188 58676
rect 219308 58636 428188 58664
rect 219308 58624 219314 58636
rect 428182 58624 428188 58636
rect 428240 58624 428246 58676
rect 374454 58556 374460 58608
rect 374512 58596 374518 58608
rect 404170 58596 404176 58608
rect 374512 58568 404176 58596
rect 374512 58556 374518 58568
rect 404170 58556 404176 58568
rect 404228 58556 404234 58608
rect 57882 57876 57888 57928
rect 57940 57916 57946 57928
rect 204898 57916 204904 57928
rect 57940 57888 204904 57916
rect 57940 57876 57946 57888
rect 204898 57876 204904 57888
rect 204956 57876 204962 57928
rect 208302 57876 208308 57928
rect 208360 57916 208366 57928
rect 325878 57916 325884 57928
rect 208360 57888 325884 57916
rect 208360 57876 208366 57888
rect 325878 57876 325884 57888
rect 325936 57876 325942 57928
rect 343174 57876 343180 57928
rect 343232 57916 343238 57928
rect 357526 57916 357532 57928
rect 343232 57888 357532 57916
rect 343232 57876 343238 57888
rect 357526 57876 357532 57888
rect 357584 57876 357590 57928
rect 364242 57876 364248 57928
rect 364300 57916 364306 57928
rect 478414 57916 478420 57928
rect 364300 57888 478420 57916
rect 364300 57876 364306 57888
rect 478414 57876 478420 57888
rect 478472 57876 478478 57928
rect 503254 57876 503260 57928
rect 503312 57916 503318 57928
rect 517606 57916 517612 57928
rect 503312 57888 517612 57916
rect 503312 57876 503318 57888
rect 517606 57876 517612 57888
rect 517664 57876 517670 57928
rect 51442 57808 51448 57860
rect 51500 57848 51506 57860
rect 145558 57848 145564 57860
rect 51500 57820 145564 57848
rect 51500 57808 51506 57820
rect 145558 57808 145564 57820
rect 145616 57808 145622 57860
rect 183278 57808 183284 57860
rect 183336 57848 183342 57860
rect 197446 57848 197452 57860
rect 183336 57820 197452 57848
rect 183336 57808 183342 57820
rect 197446 57808 197452 57820
rect 197504 57808 197510 57860
rect 211062 57808 211068 57860
rect 211120 57848 211126 57860
rect 318334 57848 318340 57860
rect 211120 57820 318340 57848
rect 211120 57808 211126 57820
rect 318334 57808 318340 57820
rect 318392 57808 318398 57860
rect 343450 57808 343456 57860
rect 343508 57848 343514 57860
rect 356698 57848 356704 57860
rect 343508 57820 356704 57848
rect 343508 57808 343514 57820
rect 356698 57808 356704 57820
rect 356756 57808 356762 57860
rect 378502 57808 378508 57860
rect 378560 57848 378566 57860
rect 470870 57848 470876 57860
rect 378560 57820 470876 57848
rect 378560 57808 378566 57820
rect 470870 57808 470876 57820
rect 470928 57808 470934 57860
rect 503530 57808 503536 57860
rect 503588 57848 503594 57860
rect 517514 57848 517520 57860
rect 503588 57820 517520 57848
rect 503588 57808 503594 57820
rect 517514 57808 517520 57820
rect 517572 57808 517578 57860
rect 41230 57740 41236 57792
rect 41288 57780 41294 57792
rect 133414 57780 133420 57792
rect 41288 57752 133420 57780
rect 41288 57740 41294 57752
rect 133414 57740 133420 57752
rect 133472 57740 133478 57792
rect 183462 57740 183468 57792
rect 183520 57780 183526 57792
rect 197354 57780 197360 57792
rect 183520 57752 197360 57780
rect 183520 57740 183526 57752
rect 197354 57740 197360 57752
rect 197412 57740 197418 57792
rect 205542 57740 205548 57792
rect 205600 57780 205606 57792
rect 310974 57780 310980 57792
rect 205600 57752 310980 57780
rect 205600 57740 205606 57752
rect 310974 57740 310980 57752
rect 311032 57740 311038 57792
rect 363598 57740 363604 57792
rect 363656 57780 363662 57792
rect 443454 57780 443460 57792
rect 363656 57752 443460 57780
rect 363656 57740 363662 57752
rect 443454 57740 443460 57752
rect 443512 57740 443518 57792
rect 41138 57672 41144 57724
rect 41196 57712 41202 57724
rect 123478 57712 123484 57724
rect 41196 57684 123484 57712
rect 41196 57672 41202 57684
rect 123478 57672 123484 57684
rect 123536 57672 123542 57724
rect 218974 57672 218980 57724
rect 219032 57712 219038 57724
rect 320910 57712 320916 57724
rect 219032 57684 320916 57712
rect 219032 57672 219038 57684
rect 320910 57672 320916 57684
rect 320968 57672 320974 57724
rect 367922 57672 367928 57724
rect 367980 57712 367986 57724
rect 448238 57712 448244 57724
rect 367980 57684 448244 57712
rect 367980 57672 367986 57684
rect 448238 57672 448244 57684
rect 448296 57672 448302 57724
rect 53742 57604 53748 57656
rect 53800 57644 53806 57656
rect 130838 57644 130844 57656
rect 53800 57616 130844 57644
rect 53800 57604 53806 57616
rect 130838 57604 130844 57616
rect 130896 57604 130902 57656
rect 213730 57604 213736 57656
rect 213788 57644 213794 57656
rect 313366 57644 313372 57656
rect 213788 57616 313372 57644
rect 213788 57604 213794 57616
rect 313366 57604 313372 57616
rect 313424 57604 313430 57656
rect 367830 57604 367836 57656
rect 367888 57644 367894 57656
rect 440878 57644 440884 57656
rect 367888 57616 440884 57644
rect 367888 57604 367894 57616
rect 440878 57604 440884 57616
rect 440936 57604 440942 57656
rect 57238 57536 57244 57588
rect 57296 57576 57302 57588
rect 57882 57576 57888 57588
rect 57296 57548 57888 57576
rect 57296 57536 57302 57548
rect 57882 57536 57888 57548
rect 57940 57536 57946 57588
rect 128354 57576 128360 57588
rect 58820 57548 128360 57576
rect 55122 57468 55128 57520
rect 55180 57508 55186 57520
rect 58820 57508 58848 57548
rect 128354 57536 128360 57548
rect 128412 57536 128418 57588
rect 209682 57536 209688 57588
rect 209740 57576 209746 57588
rect 305822 57576 305828 57588
rect 209740 57548 305828 57576
rect 209740 57536 209746 57548
rect 305822 57536 305828 57548
rect 305880 57536 305886 57588
rect 363690 57536 363696 57588
rect 363748 57576 363754 57588
rect 433610 57576 433616 57588
rect 363748 57548 433616 57576
rect 363748 57536 363754 57548
rect 433610 57536 433616 57548
rect 433668 57536 433674 57588
rect 55180 57480 58848 57508
rect 55180 57468 55186 57480
rect 58986 57468 58992 57520
rect 59044 57508 59050 57520
rect 125870 57508 125876 57520
rect 59044 57480 125876 57508
rect 59044 57468 59050 57480
rect 125870 57468 125876 57480
rect 125928 57468 125934 57520
rect 218330 57468 218336 57520
rect 218388 57508 218394 57520
rect 300854 57508 300860 57520
rect 218388 57480 300860 57508
rect 218388 57468 218394 57480
rect 300854 57468 300860 57480
rect 300912 57468 300918 57520
rect 370498 57468 370504 57520
rect 370556 57508 370562 57520
rect 438486 57508 438492 57520
rect 370556 57480 438492 57508
rect 370556 57468 370562 57480
rect 438486 57468 438492 57480
rect 438544 57468 438550 57520
rect 52086 57400 52092 57452
rect 52144 57440 52150 57452
rect 111150 57440 111156 57452
rect 52144 57412 111156 57440
rect 52144 57400 52150 57412
rect 111150 57400 111156 57412
rect 111208 57400 111214 57452
rect 279050 57400 279056 57452
rect 279108 57440 279114 57452
rect 356606 57440 356612 57452
rect 279108 57412 356612 57440
rect 279108 57400 279114 57412
rect 356606 57400 356612 57412
rect 356664 57400 356670 57452
rect 371878 57400 371884 57452
rect 371936 57440 371942 57452
rect 435910 57440 435916 57452
rect 371936 57412 435916 57440
rect 371936 57400 371942 57412
rect 435910 57400 435916 57412
rect 435968 57400 435974 57452
rect 51534 57332 51540 57384
rect 51592 57372 51598 57384
rect 88334 57372 88340 57384
rect 51592 57344 88340 57372
rect 51592 57332 51598 57344
rect 88334 57332 88340 57344
rect 88392 57332 88398 57384
rect 216490 57332 216496 57384
rect 216548 57372 216554 57384
rect 293310 57372 293316 57384
rect 216548 57344 293316 57372
rect 216548 57332 216554 57344
rect 293310 57332 293316 57344
rect 293368 57332 293374 57384
rect 376110 57332 376116 57384
rect 376168 57372 376174 57384
rect 430942 57372 430948 57384
rect 376168 57344 430948 57372
rect 376168 57332 376174 57344
rect 430942 57332 430948 57344
rect 431000 57332 431006 57384
rect 58342 57264 58348 57316
rect 58400 57304 58406 57316
rect 58986 57304 58992 57316
rect 58400 57276 58992 57304
rect 58400 57264 58406 57276
rect 58986 57264 58992 57276
rect 59044 57264 59050 57316
rect 59262 57264 59268 57316
rect 59320 57304 59326 57316
rect 90726 57304 90732 57316
rect 59320 57276 90732 57304
rect 59320 57264 59326 57276
rect 90726 57264 90732 57276
rect 90784 57264 90790 57316
rect 216582 57264 216588 57316
rect 216640 57304 216646 57316
rect 287606 57304 287612 57316
rect 216640 57276 287612 57304
rect 216640 57264 216646 57276
rect 287606 57264 287612 57276
rect 287664 57264 287670 57316
rect 365070 57264 365076 57316
rect 365128 57304 365134 57316
rect 416038 57304 416044 57316
rect 365128 57276 416044 57304
rect 365128 57264 365134 57276
rect 416038 57264 416044 57276
rect 416096 57264 416102 57316
rect 52362 57196 52368 57248
rect 52420 57236 52426 57248
rect 78214 57236 78220 57248
rect 52420 57208 78220 57236
rect 52420 57196 52426 57208
rect 78214 57196 78220 57208
rect 78272 57196 78278 57248
rect 218698 57196 218704 57248
rect 218756 57236 218762 57248
rect 265342 57236 265348 57248
rect 218756 57208 265348 57236
rect 218756 57196 218762 57208
rect 265342 57196 265348 57208
rect 265400 57196 265406 57248
rect 379698 57196 379704 57248
rect 379756 57236 379762 57248
rect 415486 57236 415492 57248
rect 379756 57208 415492 57236
rect 379756 57196 379762 57208
rect 415486 57196 415492 57208
rect 415544 57196 415550 57248
rect 54754 57128 54760 57180
rect 54812 57168 54818 57180
rect 76006 57168 76012 57180
rect 54812 57140 76012 57168
rect 54812 57128 54818 57140
rect 76006 57128 76012 57140
rect 76064 57128 76070 57180
rect 213822 57128 213828 57180
rect 213880 57168 213886 57180
rect 283650 57168 283656 57180
rect 213880 57140 283656 57168
rect 213880 57128 213886 57140
rect 283650 57128 283656 57140
rect 283708 57128 283714 57180
rect 54938 56516 54944 56568
rect 54996 56556 55002 56568
rect 81802 56556 81808 56568
rect 54996 56528 81808 56556
rect 54996 56516 55002 56528
rect 81802 56516 81808 56528
rect 81860 56516 81866 56568
rect 214466 56516 214472 56568
rect 214524 56556 214530 56568
rect 242894 56556 242900 56568
rect 214524 56528 242900 56556
rect 214524 56516 214530 56528
rect 242894 56516 242900 56528
rect 242952 56516 242958 56568
rect 376018 56516 376024 56568
rect 376076 56556 376082 56568
rect 399478 56556 399484 56568
rect 376076 56528 399484 56556
rect 376076 56516 376082 56528
rect 399478 56516 399484 56528
rect 399536 56516 399542 56568
rect 53466 56448 53472 56500
rect 53524 56488 53530 56500
rect 109218 56488 109224 56500
rect 53524 56460 109224 56488
rect 53524 56448 53530 56460
rect 109218 56448 109224 56460
rect 109276 56448 109282 56500
rect 215938 56448 215944 56500
rect 215996 56488 216002 56500
rect 239214 56488 239220 56500
rect 215996 56460 239220 56488
rect 215996 56448 216002 56460
rect 239214 56448 239220 56460
rect 239272 56448 239278 56500
rect 372246 56448 372252 56500
rect 372304 56488 372310 56500
rect 435726 56488 435732 56500
rect 372304 56460 435732 56488
rect 372304 56448 372310 56460
rect 435726 56448 435732 56460
rect 435784 56448 435790 56500
rect 59906 56380 59912 56432
rect 59964 56420 59970 56432
rect 108022 56420 108028 56432
rect 59964 56392 108028 56420
rect 59964 56380 59970 56392
rect 108022 56380 108028 56392
rect 108080 56380 108086 56432
rect 219158 56380 219164 56432
rect 219216 56420 219222 56432
rect 235994 56420 236000 56432
rect 219216 56392 236000 56420
rect 219216 56380 219222 56392
rect 235994 56380 236000 56392
rect 236052 56380 236058 56432
rect 378410 56380 378416 56432
rect 378468 56420 378474 56432
rect 438210 56420 438216 56432
rect 378468 56392 438216 56420
rect 378468 56380 378474 56392
rect 438210 56380 438216 56392
rect 438268 56380 438274 56432
rect 57790 56312 57796 56364
rect 57848 56352 57854 56364
rect 104986 56352 104992 56364
rect 57848 56324 104992 56352
rect 57848 56312 57854 56324
rect 104986 56312 104992 56324
rect 105044 56312 105050 56364
rect 214926 56312 214932 56364
rect 214984 56352 214990 56364
rect 269758 56352 269764 56364
rect 214984 56324 269764 56352
rect 214984 56312 214990 56324
rect 269758 56312 269764 56324
rect 269816 56312 269822 56364
rect 374914 56312 374920 56364
rect 374972 56352 374978 56364
rect 432230 56352 432236 56364
rect 374972 56324 432236 56352
rect 374972 56312 374978 56324
rect 432230 56312 432236 56324
rect 432288 56312 432294 56364
rect 59170 56244 59176 56296
rect 59228 56284 59234 56296
rect 106734 56284 106740 56296
rect 59228 56256 106740 56284
rect 59228 56244 59234 56256
rect 106734 56244 106740 56256
rect 106792 56244 106798 56296
rect 218238 56244 218244 56296
rect 218296 56284 218302 56296
rect 266998 56284 267004 56296
rect 218296 56256 267004 56284
rect 218296 56244 218302 56256
rect 266998 56244 267004 56256
rect 267056 56244 267062 56296
rect 379422 56244 379428 56296
rect 379480 56284 379486 56296
rect 427630 56284 427636 56296
rect 379480 56256 427636 56284
rect 379480 56244 379486 56256
rect 427630 56244 427636 56256
rect 427688 56244 427694 56296
rect 56410 56176 56416 56228
rect 56468 56216 56474 56228
rect 103790 56216 103796 56228
rect 56468 56188 103796 56216
rect 56468 56176 56474 56188
rect 103790 56176 103796 56188
rect 103848 56176 103854 56228
rect 219802 56176 219808 56228
rect 219860 56216 219866 56228
rect 266354 56216 266360 56228
rect 219860 56188 266360 56216
rect 219860 56176 219866 56188
rect 266354 56176 266360 56188
rect 266412 56176 266418 56228
rect 379882 56176 379888 56228
rect 379940 56216 379946 56228
rect 426434 56216 426440 56228
rect 379940 56188 426440 56216
rect 379940 56176 379946 56188
rect 426434 56176 426440 56188
rect 426492 56176 426498 56228
rect 59998 56108 60004 56160
rect 60056 56148 60062 56160
rect 106366 56148 106372 56160
rect 60056 56120 106372 56148
rect 60056 56108 60062 56120
rect 106366 56108 106372 56120
rect 106424 56108 106430 56160
rect 218790 56108 218796 56160
rect 218848 56148 218854 56160
rect 253382 56148 253388 56160
rect 218848 56120 253388 56148
rect 218848 56108 218854 56120
rect 253382 56108 253388 56120
rect 253440 56108 253446 56160
rect 379790 56108 379796 56160
rect 379848 56148 379854 56160
rect 414566 56148 414572 56160
rect 379848 56120 414572 56148
rect 379848 56108 379854 56120
rect 414566 56108 414572 56120
rect 414624 56108 414630 56160
rect 58802 56040 58808 56092
rect 58860 56080 58866 56092
rect 92106 56080 92112 56092
rect 58860 56052 92112 56080
rect 58860 56040 58866 56052
rect 92106 56040 92112 56052
rect 92164 56040 92170 56092
rect 219066 56040 219072 56092
rect 219124 56080 219130 56092
rect 251174 56080 251180 56092
rect 219124 56052 251180 56080
rect 219124 56040 219130 56052
rect 251174 56040 251180 56052
rect 251232 56040 251238 56092
rect 378870 56040 378876 56092
rect 378928 56080 378934 56092
rect 412634 56080 412640 56092
rect 378928 56052 412640 56080
rect 378928 56040 378934 56052
rect 412634 56040 412640 56052
rect 412692 56040 412698 56092
rect 56318 55972 56324 56024
rect 56376 56012 56382 56024
rect 88702 56012 88708 56024
rect 56376 55984 88708 56012
rect 56376 55972 56382 55984
rect 88702 55972 88708 55984
rect 88760 55972 88766 56024
rect 214742 55972 214748 56024
rect 214800 56012 214806 56024
rect 246390 56012 246396 56024
rect 214800 55984 246396 56012
rect 214800 55972 214806 55984
rect 246390 55972 246396 55984
rect 246448 55972 246454 56024
rect 379146 55972 379152 56024
rect 379204 56012 379210 56024
rect 411254 56012 411260 56024
rect 379204 55984 411260 56012
rect 379204 55972 379210 55984
rect 411254 55972 411260 55984
rect 411312 55972 411318 56024
rect 54846 55904 54852 55956
rect 54904 55944 54910 55956
rect 86494 55944 86500 55956
rect 54904 55916 86500 55944
rect 54904 55904 54910 55916
rect 86494 55904 86500 55916
rect 86552 55904 86558 55956
rect 218606 55904 218612 55956
rect 218664 55944 218670 55956
rect 248598 55944 248604 55956
rect 218664 55916 248604 55944
rect 218664 55904 218670 55916
rect 248598 55904 248604 55916
rect 248656 55904 248662 55956
rect 378962 55904 378968 55956
rect 379020 55944 379026 55956
rect 408678 55944 408684 55956
rect 379020 55916 408684 55944
rect 379020 55904 379026 55916
rect 408678 55904 408684 55916
rect 408736 55904 408742 55956
rect 58710 55836 58716 55888
rect 58768 55876 58774 55888
rect 85390 55876 85396 55888
rect 58768 55848 85396 55876
rect 58768 55836 58774 55848
rect 85390 55836 85396 55848
rect 85448 55836 85454 55888
rect 213362 55836 213368 55888
rect 213420 55876 213426 55888
rect 273622 55876 273628 55888
rect 213420 55848 273628 55876
rect 213420 55836 213426 55848
rect 273622 55836 273628 55848
rect 273680 55836 273686 55888
rect 372338 55836 372344 55888
rect 372396 55876 372402 55888
rect 401686 55876 401692 55888
rect 372396 55848 401692 55876
rect 372396 55836 372402 55848
rect 401686 55836 401692 55848
rect 401744 55836 401750 55888
rect 53558 55768 53564 55820
rect 53616 55808 53622 55820
rect 115750 55808 115756 55820
rect 53616 55780 115756 55808
rect 53616 55768 53622 55780
rect 115750 55768 115756 55780
rect 115808 55768 115814 55820
rect 219986 55768 219992 55820
rect 220044 55808 220050 55820
rect 408310 55808 408316 55820
rect 220044 55780 408316 55808
rect 220044 55768 220050 55780
rect 408310 55768 408316 55780
rect 408368 55768 408374 55820
rect 51902 55700 51908 55752
rect 51960 55740 51966 55752
rect 79502 55740 79508 55752
rect 51960 55712 79508 55740
rect 51960 55700 51966 55712
rect 79502 55700 79508 55712
rect 79560 55700 79566 55752
rect 215846 55700 215852 55752
rect 215904 55740 215910 55752
rect 272150 55740 272156 55752
rect 215904 55712 272156 55740
rect 215904 55700 215910 55712
rect 272150 55700 272156 55712
rect 272208 55700 272214 55752
rect 44082 55156 44088 55208
rect 44140 55196 44146 55208
rect 115934 55196 115940 55208
rect 44140 55168 115940 55196
rect 44140 55156 44146 55168
rect 115934 55156 115940 55168
rect 115992 55156 115998 55208
rect 213546 55156 213552 55208
rect 213604 55196 213610 55208
rect 274634 55196 274640 55208
rect 213604 55168 274640 55196
rect 213604 55156 213610 55168
rect 274634 55156 274640 55168
rect 274692 55156 274698 55208
rect 376386 55156 376392 55208
rect 376444 55196 376450 55208
rect 436094 55196 436100 55208
rect 376444 55168 436100 55196
rect 376444 55156 376450 55168
rect 436094 55156 436100 55168
rect 436152 55156 436158 55208
rect 53282 55088 53288 55140
rect 53340 55128 53346 55140
rect 113174 55128 113180 55140
rect 53340 55100 113180 55128
rect 53340 55088 53346 55100
rect 113174 55088 113180 55100
rect 113232 55088 113238 55140
rect 214834 55088 214840 55140
rect 214892 55128 214898 55140
rect 273346 55128 273352 55140
rect 214892 55100 273352 55128
rect 214892 55088 214898 55100
rect 273346 55088 273352 55100
rect 273404 55088 273410 55140
rect 375006 55088 375012 55140
rect 375064 55128 375070 55140
rect 433334 55128 433340 55140
rect 375064 55100 433340 55128
rect 375064 55088 375070 55100
rect 433334 55088 433340 55100
rect 433392 55088 433398 55140
rect 52178 55020 52184 55072
rect 52236 55060 52242 55072
rect 111794 55060 111800 55072
rect 52236 55032 111800 55060
rect 52236 55020 52242 55032
rect 111794 55020 111800 55032
rect 111852 55020 111858 55072
rect 214650 55020 214656 55072
rect 214708 55060 214714 55072
rect 270494 55060 270500 55072
rect 214708 55032 270500 55060
rect 214708 55020 214714 55032
rect 270494 55020 270500 55032
rect 270552 55020 270558 55072
rect 375558 55020 375564 55072
rect 375616 55060 375622 55072
rect 433426 55060 433432 55072
rect 375616 55032 433432 55060
rect 375616 55020 375622 55032
rect 433426 55020 433432 55032
rect 433484 55020 433490 55072
rect 58618 54952 58624 55004
rect 58676 54992 58682 55004
rect 92474 54992 92480 55004
rect 58676 54964 92480 54992
rect 58676 54952 58682 54964
rect 92474 54952 92480 54964
rect 92532 54952 92538 55004
rect 219526 54952 219532 55004
rect 219584 54992 219590 55004
rect 267734 54992 267740 55004
rect 219584 54964 267740 54992
rect 219584 54952 219590 54964
rect 267734 54952 267740 54964
rect 267792 54952 267798 55004
rect 374822 54952 374828 55004
rect 374880 54992 374886 55004
rect 430574 54992 430580 55004
rect 374880 54964 430580 54992
rect 374880 54952 374886 54964
rect 430574 54952 430580 54964
rect 430632 54952 430638 55004
rect 56962 54884 56968 54936
rect 57020 54924 57026 54936
rect 91186 54924 91192 54936
rect 57020 54896 91192 54924
rect 57020 54884 57026 54896
rect 91186 54884 91192 54896
rect 91244 54884 91250 54936
rect 219894 54884 219900 54936
rect 219952 54924 219958 54936
rect 253934 54924 253940 54936
rect 219952 54896 253940 54924
rect 219952 54884 219958 54896
rect 253934 54884 253940 54896
rect 253992 54884 253998 54936
rect 376294 54884 376300 54936
rect 376352 54924 376358 54936
rect 429194 54924 429200 54936
rect 376352 54896 429200 54924
rect 376352 54884 376358 54896
rect 429194 54884 429200 54896
rect 429252 54884 429258 54936
rect 53190 54816 53196 54868
rect 53248 54856 53254 54868
rect 86954 54856 86960 54868
rect 53248 54828 86960 54856
rect 53248 54816 53254 54828
rect 86954 54816 86960 54828
rect 87012 54816 87018 54868
rect 217870 54816 217876 54868
rect 217928 54856 217934 54868
rect 251358 54856 251364 54868
rect 217928 54828 251364 54856
rect 217928 54816 217934 54828
rect 251358 54816 251364 54828
rect 251416 54816 251422 54868
rect 379974 54816 379980 54868
rect 380032 54856 380038 54868
rect 427814 54856 427820 54868
rect 380032 54828 427820 54856
rect 380032 54816 380038 54828
rect 427814 54816 427820 54828
rect 427872 54816 427878 54868
rect 58894 54748 58900 54800
rect 58952 54788 58958 54800
rect 89714 54788 89720 54800
rect 58952 54760 89720 54788
rect 58952 54748 58958 54760
rect 89714 54748 89720 54760
rect 89772 54748 89778 54800
rect 216214 54748 216220 54800
rect 216272 54788 216278 54800
rect 247034 54788 247040 54800
rect 216272 54760 247040 54788
rect 216272 54748 216278 54760
rect 247034 54748 247040 54760
rect 247092 54748 247098 54800
rect 377030 54748 377036 54800
rect 377088 54788 377094 54800
rect 411346 54788 411352 54800
rect 377088 54760 411352 54788
rect 377088 54748 377094 54760
rect 411346 54748 411352 54760
rect 411404 54748 411410 54800
rect 53374 54680 53380 54732
rect 53432 54720 53438 54732
rect 80054 54720 80060 54732
rect 53432 54692 80060 54720
rect 53432 54680 53438 54692
rect 80054 54680 80060 54692
rect 80112 54680 80118 54732
rect 212166 54680 212172 54732
rect 212224 54720 212230 54732
rect 241514 54720 241520 54732
rect 212224 54692 241520 54720
rect 212224 54680 212230 54692
rect 241514 54680 241520 54692
rect 241572 54680 241578 54732
rect 377214 54680 377220 54732
rect 377272 54720 377278 54732
rect 409874 54720 409880 54732
rect 377272 54692 409880 54720
rect 377272 54680 377278 54692
rect 409874 54680 409880 54692
rect 409932 54680 409938 54732
rect 215018 54612 215024 54664
rect 215076 54652 215082 54664
rect 244274 54652 244280 54664
rect 215076 54624 244280 54652
rect 215076 54612 215082 54624
rect 244274 54612 244280 54624
rect 244332 54612 244338 54664
rect 375098 54612 375104 54664
rect 375156 54652 375162 54664
rect 405826 54652 405832 54664
rect 375156 54624 405832 54652
rect 375156 54612 375162 54624
rect 405826 54612 405832 54624
rect 405884 54612 405890 54664
rect 216306 54544 216312 54596
rect 216364 54584 216370 54596
rect 244366 54584 244372 54596
rect 216364 54556 244372 54584
rect 216364 54544 216370 54556
rect 244366 54544 244372 54556
rect 244424 54544 244430 54596
rect 376570 54544 376576 54596
rect 376628 54584 376634 54596
rect 407206 54584 407212 54596
rect 376628 54556 407212 54584
rect 376628 54544 376634 54556
rect 407206 54544 407212 54556
rect 407264 54544 407270 54596
rect 213270 54476 213276 54528
rect 213328 54516 213334 54528
rect 240134 54516 240140 54528
rect 213328 54488 240140 54516
rect 213328 54476 213334 54488
rect 240134 54476 240140 54488
rect 240192 54476 240198 54528
rect 376202 54476 376208 54528
rect 376260 54516 376266 54528
rect 404354 54516 404360 54528
rect 376260 54488 404360 54516
rect 376260 54476 376266 54488
rect 404354 54476 404360 54488
rect 404412 54476 404418 54528
rect 214558 54408 214564 54460
rect 214616 54448 214622 54460
rect 237374 54448 237380 54460
rect 214616 54420 237380 54448
rect 214616 54408 214622 54420
rect 237374 54408 237380 54420
rect 237432 54408 237438 54460
rect 372154 54408 372160 54460
rect 372212 54448 372218 54460
rect 400214 54448 400220 54460
rect 372212 54420 400220 54448
rect 372212 54408 372218 54420
rect 400214 54408 400220 54420
rect 400272 54408 400278 54460
rect 374730 54340 374736 54392
rect 374788 54380 374794 54392
rect 397454 54380 397460 54392
rect 374788 54352 397460 54380
rect 374788 54340 374794 54352
rect 397454 54340 397460 54352
rect 397512 54340 397518 54392
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 4798 20380 4804 20392
rect 2832 20352 4804 20380
rect 2832 20340 2838 20352
rect 4798 20340 4804 20352
rect 4856 20340 4862 20392
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 57238 3448 57244 3460
rect 624 3420 57244 3448
rect 624 3408 630 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
<< via1 >>
rect 235172 700340 235224 700392
rect 305644 700340 305696 700392
rect 57888 700272 57940 700324
rect 543464 700272 543516 700324
rect 137928 683136 137980 683188
rect 580172 683136 580224 683188
rect 169760 640976 169812 641028
rect 430948 640976 431000 641028
rect 3424 639548 3476 639600
rect 317052 639548 317104 639600
rect 104900 638188 104952 638240
rect 429292 638188 429344 638240
rect 299480 636828 299532 636880
rect 401140 636828 401192 636880
rect 364340 635468 364392 635520
rect 423680 635468 423732 635520
rect 316960 634924 317012 634976
rect 430580 634924 430632 634976
rect 316868 634856 316920 634908
rect 430856 634856 430908 634908
rect 291200 634788 291252 634840
rect 457444 634788 457496 634840
rect 318800 634040 318852 634092
rect 494060 634040 494112 634092
rect 280988 633632 281040 633684
rect 383108 633632 383160 633684
rect 281080 633564 281132 633616
rect 430764 633564 430816 633616
rect 289820 633496 289872 633548
rect 489920 633496 489972 633548
rect 288440 633428 288492 633480
rect 512000 633428 512052 633480
rect 313924 632952 313976 633004
rect 337384 632952 337436 633004
rect 309784 632884 309836 632936
rect 332876 632884 332928 632936
rect 295984 632816 296036 632868
rect 378600 632816 378652 632868
rect 291292 632748 291344 632800
rect 432604 632748 432656 632800
rect 319536 632680 319588 632732
rect 355416 632680 355468 632732
rect 311164 632612 311216 632664
rect 350908 632612 350960 632664
rect 319720 632544 319772 632596
rect 364432 632544 364484 632596
rect 312544 632476 312596 632528
rect 359924 632476 359976 632528
rect 319812 632408 319864 632460
rect 373448 632408 373500 632460
rect 316776 632340 316828 632392
rect 387616 632340 387668 632392
rect 316684 632272 316736 632324
rect 396632 632272 396684 632324
rect 320824 632204 320876 632256
rect 341892 632204 341944 632256
rect 318248 632136 318300 632188
rect 428188 632136 428240 632188
rect 319904 632068 319956 632120
rect 323860 632068 323912 632120
rect 284944 631320 284996 631372
rect 368940 631320 368992 631372
rect 318064 631252 318116 631304
rect 430672 631252 430724 631304
rect 298100 631184 298152 631236
rect 429844 631184 429896 631236
rect 296812 631116 296864 631168
rect 435364 631116 435416 631168
rect 293960 631048 294012 631100
rect 432696 631048 432748 631100
rect 288532 630980 288584 631032
rect 428464 630980 428516 631032
rect 319444 630912 319496 630964
rect 466736 630912 466788 630964
rect 296720 630844 296772 630896
rect 510620 630844 510672 630896
rect 319076 630776 319128 630828
rect 580172 630776 580224 630828
rect 18604 630708 18656 630760
rect 409880 630708 409932 630760
rect 218704 630640 218756 630692
rect 414388 630640 414440 630692
rect 280712 629960 280764 630012
rect 320824 630436 320876 630488
rect 217784 629892 217836 629944
rect 319076 629892 319128 629944
rect 314016 629280 314068 629332
rect 317788 629280 317840 629332
rect 214012 625744 214064 625796
rect 225420 625744 225472 625796
rect 100576 625676 100628 625728
rect 124312 625676 124364 625728
rect 137836 625676 137888 625728
rect 186504 625676 186556 625728
rect 206468 625676 206520 625728
rect 231308 625676 231360 625728
rect 112168 625608 112220 625660
rect 122840 625608 122892 625660
rect 135168 625608 135220 625660
rect 160284 625608 160336 625660
rect 212540 625608 212592 625660
rect 271880 625608 271932 625660
rect 94780 625540 94832 625592
rect 122288 625540 122340 625592
rect 136456 625540 136508 625592
rect 162860 625540 162912 625592
rect 217876 625540 217928 625592
rect 242900 625540 242952 625592
rect 83188 625472 83240 625524
rect 124404 625472 124456 625524
rect 139216 625472 139268 625524
rect 166172 625472 166224 625524
rect 218888 625472 218940 625524
rect 251916 625472 251968 625524
rect 109592 625404 109644 625456
rect 120908 625404 120960 625456
rect 139124 625404 139176 625456
rect 174452 625404 174504 625456
rect 218796 625404 218848 625456
rect 263600 625404 263652 625456
rect 103796 625336 103848 625388
rect 121644 625336 121696 625388
rect 137744 625336 137796 625388
rect 180340 625336 180392 625388
rect 190000 625336 190052 625388
rect 204536 625336 204588 625388
rect 209780 625336 209832 625388
rect 260196 625336 260248 625388
rect 54852 625268 54904 625320
rect 88984 625268 89036 625320
rect 124220 625268 124272 625320
rect 171876 625268 171928 625320
rect 213920 625268 213972 625320
rect 269212 625268 269264 625320
rect 55128 625200 55180 625252
rect 92204 625200 92256 625252
rect 115388 625200 115440 625252
rect 124680 625200 124732 625252
rect 135260 625200 135312 625252
rect 183652 625200 183704 625252
rect 192576 625200 192628 625252
rect 204444 625200 204496 625252
rect 219348 625200 219400 625252
rect 275100 625200 275152 625252
rect 56508 625132 56560 625184
rect 77392 625132 77444 625184
rect 133880 625132 133932 625184
rect 139860 625132 139912 625184
rect 157524 625132 157576 625184
rect 195704 625132 195756 625184
rect 201684 625132 201736 625184
rect 140136 625064 140188 625116
rect 215300 624044 215352 624096
rect 234620 624044 234672 624096
rect 219624 623976 219676 624028
rect 246028 623976 246080 624028
rect 59360 623908 59412 623960
rect 98000 623908 98052 623960
rect 210424 623908 210476 623960
rect 237564 623908 237616 623960
rect 57796 623840 57848 623892
rect 80612 623840 80664 623892
rect 86408 623840 86460 623892
rect 124588 623840 124640 623892
rect 133144 623840 133196 623892
rect 151268 623840 151320 623892
rect 206284 623840 206336 623892
rect 254492 623840 254544 623892
rect 69020 623772 69072 623824
rect 124496 623772 124548 623824
rect 136640 623772 136692 623824
rect 168748 623772 168800 623824
rect 204260 623772 204312 623824
rect 277676 623772 277728 623824
rect 217968 622820 218020 622872
rect 228732 622820 228784 622872
rect 126244 622752 126296 622804
rect 177856 622752 177908 622804
rect 214564 622752 214616 622804
rect 257620 622752 257672 622804
rect 136364 622684 136416 622736
rect 145564 622684 145616 622736
rect 204352 622684 204404 622736
rect 222844 622684 222896 622736
rect 56324 622616 56376 622668
rect 74632 622616 74684 622668
rect 135076 622616 135128 622668
rect 149152 622616 149204 622668
rect 208400 622616 208452 622668
rect 240324 622616 240376 622668
rect 54944 622548 54996 622600
rect 65524 622548 65576 622600
rect 134892 622548 134944 622600
rect 154580 622548 154632 622600
rect 206376 622548 206428 622600
rect 248696 622548 248748 622600
rect 56416 622480 56468 622532
rect 71228 622480 71280 622532
rect 134984 622480 135036 622532
rect 142988 622480 143040 622532
rect 211804 622480 211856 622532
rect 266268 622480 266320 622532
rect 280712 622480 280764 622532
rect 55036 622412 55088 622464
rect 62948 622412 63000 622464
rect 136548 622412 136600 622464
rect 218704 622412 218756 622464
rect 118240 622344 118292 622396
rect 121552 622344 121604 622396
rect 198280 622344 198332 622396
rect 201500 622344 201552 622396
rect 217324 622344 217376 622396
rect 219716 622344 219768 622396
rect 280712 622276 280764 622328
rect 435364 621800 435416 621852
rect 474832 621800 474884 621852
rect 432696 621732 432748 621784
rect 498016 621732 498068 621784
rect 429844 621664 429896 621716
rect 505744 621664 505796 621716
rect 482560 620984 482612 621036
rect 509884 620984 509936 621036
rect 213184 619624 213236 619676
rect 216680 619624 216732 619676
rect 302884 619624 302936 619676
rect 317972 619624 318024 619676
rect 432604 619556 432656 619608
rect 456800 619556 456852 619608
rect 208492 616836 208544 616888
rect 216680 616836 216732 616888
rect 286324 615476 286376 615528
rect 317972 615476 318024 615528
rect 428464 611260 428516 611312
rect 456800 611260 456852 611312
rect 307024 609968 307076 610020
rect 317880 609968 317932 610020
rect 132500 607180 132552 607232
rect 136732 607180 136784 607232
rect 204904 607180 204956 607232
rect 216680 607180 216732 607232
rect 304264 605820 304316 605872
rect 317972 605820 318024 605872
rect 289084 600312 289136 600364
rect 317604 600312 317656 600364
rect 286416 596164 286468 596216
rect 317604 596164 317656 596216
rect 134524 594804 134576 594856
rect 136548 594804 136600 594856
rect 207020 593376 207072 593428
rect 216680 593376 216732 593428
rect 210516 589364 210568 589416
rect 216680 589364 216732 589416
rect 124128 589296 124180 589348
rect 131764 589296 131816 589348
rect 134616 589296 134668 589348
rect 136916 589296 136968 589348
rect 204168 589296 204220 589348
rect 216772 589296 216824 589348
rect 283564 589296 283616 589348
rect 302240 589296 302292 589348
rect 211160 586848 211212 586900
rect 216680 586848 216732 586900
rect 300124 586508 300176 586560
rect 317420 586508 317472 586560
rect 57520 583720 57572 583772
rect 58624 583720 58676 583772
rect 291844 582360 291896 582412
rect 317972 582360 318024 582412
rect 217692 581680 217744 581732
rect 218704 581680 218756 581732
rect 509884 578144 509936 578196
rect 580172 578144 580224 578196
rect 125600 576852 125652 576904
rect 136732 576852 136784 576904
rect 287704 576852 287756 576904
rect 317880 576852 317932 576904
rect 206560 574064 206612 574116
rect 216680 574064 216732 574116
rect 57336 572296 57388 572348
rect 58716 572296 58768 572348
rect 210608 571344 210660 571396
rect 216680 571344 216732 571396
rect 286508 571344 286560 571396
rect 317972 571344 318024 571396
rect 209044 562300 209096 562352
rect 217416 562300 217468 562352
rect 319352 562300 319404 562352
rect 319812 562300 319864 562352
rect 281540 562232 281592 562284
rect 282092 562232 282144 562284
rect 57888 561144 57940 561196
rect 134524 561144 134576 561196
rect 3424 561076 3476 561128
rect 291844 561076 291896 561128
rect 217692 560260 217744 560312
rect 220176 560260 220228 560312
rect 57152 560192 57204 560244
rect 62120 560192 62172 560244
rect 131764 560192 131816 560244
rect 216772 560192 216824 560244
rect 302240 560192 302292 560244
rect 137652 560124 137704 560176
rect 140780 560124 140832 560176
rect 106280 560056 106332 560108
rect 124680 560056 124732 560108
rect 98092 559988 98144 560040
rect 120908 559988 120960 560040
rect 182364 559988 182416 560040
rect 218888 559988 218940 560040
rect 255964 559988 256016 560040
rect 282920 559988 282972 560040
rect 96804 559920 96856 559972
rect 122840 559920 122892 559972
rect 164332 559920 164384 559972
rect 201684 559920 201736 559972
rect 273260 559920 273312 559972
rect 318248 559920 318300 559972
rect 57060 559852 57112 559904
rect 67732 559852 67784 559904
rect 93860 559852 93912 559904
rect 124312 559852 124364 559904
rect 157984 559852 158036 559904
rect 203248 559852 203300 559904
rect 260840 559852 260892 559904
rect 316868 559852 316920 559904
rect 59084 559784 59136 559836
rect 82912 559784 82964 559836
rect 87052 559784 87104 559836
rect 121552 559784 121604 559836
rect 139032 559784 139084 559836
rect 150624 559784 150676 559836
rect 156144 559784 156196 559836
rect 204536 559784 204588 559836
rect 258080 559784 258132 559836
rect 316960 559784 317012 559836
rect 54852 559716 54904 559768
rect 78680 559716 78732 559768
rect 85580 559716 85632 559768
rect 121736 559716 121788 559768
rect 139308 559716 139360 559768
rect 160100 559716 160152 559768
rect 182272 559716 182324 559768
rect 281540 559716 281592 559768
rect 67640 559648 67692 559700
rect 121828 559648 121880 559700
rect 137744 559648 137796 559700
rect 151820 559648 151872 559700
rect 154580 559648 154632 559700
rect 204444 559648 204496 559700
rect 216128 559648 216180 559700
rect 283012 559648 283064 559700
rect 302240 559648 302292 559700
rect 302976 559648 303028 559700
rect 63500 559580 63552 559632
rect 123024 559580 123076 559632
rect 139216 559580 139268 559632
rect 161664 559580 161716 559632
rect 179696 559580 179748 559632
rect 282092 559580 282144 559632
rect 3424 559512 3476 559564
rect 286324 559512 286376 559564
rect 217876 559308 217928 559360
rect 222200 559308 222252 559360
rect 139124 559036 139176 559088
rect 142160 559036 142212 559088
rect 219348 559036 219400 559088
rect 223580 559036 223632 559088
rect 57428 558832 57480 558884
rect 60740 558832 60792 558884
rect 100760 558764 100812 558816
rect 102876 558764 102928 558816
rect 116584 558764 116636 558816
rect 120172 558764 120224 558816
rect 161572 558764 161624 558816
rect 168472 558764 168524 558816
rect 173900 558764 173952 558816
rect 179604 558764 179656 558816
rect 225144 558764 225196 558816
rect 227996 558764 228048 558816
rect 260104 558764 260156 558816
rect 262772 558764 262824 558816
rect 278044 558764 278096 558816
rect 280252 558764 280304 558816
rect 60280 558696 60332 558748
rect 62764 558696 62816 558748
rect 119344 558696 119396 558748
rect 120724 558696 120776 558748
rect 147680 558628 147732 558680
rect 162308 558628 162360 558680
rect 151360 558560 151412 558612
rect 164884 558560 164936 558612
rect 231952 558560 232004 558612
rect 259644 558560 259696 558612
rect 142896 558492 142948 558544
rect 160744 558492 160796 558544
rect 199384 558492 199436 558544
rect 202972 558492 203024 558544
rect 222292 558492 222344 558544
rect 253940 558492 253992 558544
rect 68744 558424 68796 558476
rect 71044 558424 71096 558476
rect 82728 558424 82780 558476
rect 88984 558424 89036 558476
rect 140320 558424 140372 558476
rect 159364 558424 159416 558476
rect 188344 558424 188396 558476
rect 200212 558424 200264 558476
rect 212632 558424 212684 558476
rect 251180 558424 251232 558476
rect 77024 558356 77076 558408
rect 85672 558356 85724 558408
rect 94504 558356 94556 558408
rect 104164 558356 104216 558408
rect 111892 558356 111944 558408
rect 123116 558356 123168 558408
rect 129740 558356 129792 558408
rect 153844 558356 153896 558408
rect 154672 558356 154724 558408
rect 171324 558356 171376 558408
rect 187884 558356 187936 558408
rect 233884 558356 233936 558408
rect 62856 558288 62908 558340
rect 80704 558288 80756 558340
rect 86040 558288 86092 558340
rect 108304 558288 108356 558340
rect 112444 558288 112496 558340
rect 117412 558288 117464 558340
rect 118700 558288 118752 558340
rect 144920 558288 144972 558340
rect 158720 558288 158772 558340
rect 182916 558288 182968 558340
rect 190460 558288 190512 558340
rect 257068 558288 257120 558340
rect 269120 558288 269172 558340
rect 287704 558288 287756 558340
rect 71320 558220 71372 558272
rect 93952 558220 94004 558272
rect 100208 558220 100260 558272
rect 115204 558220 115256 558272
rect 133972 558220 134024 558272
rect 197452 558220 197504 558272
rect 199476 558220 199528 558272
rect 203156 558220 203208 558272
rect 227720 558220 227772 558272
rect 245660 558220 245712 558272
rect 249800 558220 249852 558272
rect 319812 558220 319864 558272
rect 58900 558152 58952 558204
rect 74540 558152 74592 558204
rect 79876 558152 79928 558204
rect 114560 558152 114612 558204
rect 132592 558152 132644 558204
rect 177028 558152 177080 558204
rect 177304 558152 177356 558204
rect 188620 558152 188672 558204
rect 191840 558152 191892 558204
rect 276940 558152 276992 558204
rect 71780 557880 71832 557932
rect 73804 557880 73856 557932
rect 184204 557880 184256 557932
rect 185492 557880 185544 557932
rect 264244 557880 264296 557932
rect 265348 557880 265400 557932
rect 262864 557608 262916 557660
rect 268660 557608 268712 557660
rect 64144 557540 64196 557592
rect 65064 557540 65116 557592
rect 222936 557540 222988 557592
rect 224408 557540 224460 557592
rect 267740 557540 267792 557592
rect 317420 557540 317472 557592
rect 219256 557472 219308 557524
rect 223672 557472 223724 557524
rect 178040 557064 178092 557116
rect 206560 557064 206612 557116
rect 57336 556996 57388 557048
rect 81716 556996 81768 557048
rect 122840 556996 122892 557048
rect 202236 556996 202288 557048
rect 78864 556928 78916 556980
rect 121460 556928 121512 556980
rect 137468 556928 137520 556980
rect 149060 556928 149112 556980
rect 194600 556928 194652 556980
rect 283564 556928 283616 556980
rect 63776 556860 63828 556912
rect 122932 556860 122984 556912
rect 138480 556860 138532 556912
rect 159088 556860 159140 556912
rect 159824 556860 159876 556912
rect 173440 556860 173492 556912
rect 179512 556860 179564 556912
rect 281632 556860 281684 556912
rect 4804 556792 4856 556844
rect 318340 556792 318392 556844
rect 193220 555704 193272 555756
rect 218796 555704 218848 555756
rect 143540 555636 143592 555688
rect 201868 555636 201920 555688
rect 228640 555636 228692 555688
rect 281724 555636 281776 555688
rect 59268 555568 59320 555620
rect 92572 555568 92624 555620
rect 100392 555568 100444 555620
rect 123484 555568 123536 555620
rect 126152 555568 126204 555620
rect 200764 555568 200816 555620
rect 242900 555568 242952 555620
rect 316776 555568 316828 555620
rect 64880 555500 64932 555552
rect 122196 555500 122248 555552
rect 138664 555500 138716 555552
rect 174912 555500 174964 555552
rect 181352 555500 181404 555552
rect 281816 555500 281868 555552
rect 3516 555432 3568 555484
rect 319812 555432 319864 555484
rect 171324 554208 171376 554260
rect 203340 554208 203392 554260
rect 266544 554208 266596 554260
rect 311164 554208 311216 554260
rect 73252 554140 73304 554192
rect 108580 554140 108632 554192
rect 124312 554140 124364 554192
rect 201132 554140 201184 554192
rect 229284 554140 229336 554192
rect 281264 554140 281316 554192
rect 58532 554072 58584 554124
rect 110420 554072 110472 554124
rect 198004 554072 198056 554124
rect 283104 554072 283156 554124
rect 66720 554004 66772 554056
rect 121184 554004 121236 554056
rect 138848 554004 138900 554056
rect 160560 554004 160612 554056
rect 186320 554004 186372 554056
rect 283196 554004 283248 554056
rect 219532 553596 219584 553648
rect 219900 553596 219952 553648
rect 3516 553392 3568 553444
rect 317972 553392 318024 553444
rect 226432 552916 226484 552968
rect 280804 552916 280856 552968
rect 59452 552848 59504 552900
rect 75920 552848 75972 552900
rect 88616 552848 88668 552900
rect 103520 552848 103572 552900
rect 106924 552848 106976 552900
rect 123392 552848 123444 552900
rect 129004 552848 129056 552900
rect 203064 552848 203116 552900
rect 255320 552848 255372 552900
rect 315304 552848 315356 552900
rect 75276 552780 75328 552832
rect 96988 552780 97040 552832
rect 121460 552780 121512 552832
rect 201040 552780 201092 552832
rect 247960 552780 248012 552832
rect 319352 552780 319404 552832
rect 57704 552712 57756 552764
rect 77392 552712 77444 552764
rect 80060 552712 80112 552764
rect 120816 552712 120868 552764
rect 195980 552712 196032 552764
rect 283288 552712 283340 552764
rect 69020 552644 69072 552696
rect 114652 552644 114704 552696
rect 138940 552644 138992 552696
rect 166264 552644 166316 552696
rect 179144 552644 179196 552696
rect 271236 552644 271288 552696
rect 279516 552644 279568 552696
rect 302884 552644 302936 552696
rect 192116 551556 192168 551608
rect 217324 551556 217376 551608
rect 259460 551556 259512 551608
rect 314016 551556 314068 551608
rect 80980 551488 81032 551540
rect 122104 551488 122156 551540
rect 176660 551488 176712 551540
rect 210516 551488 210568 551540
rect 253664 551488 253716 551540
rect 316684 551488 316736 551540
rect 57520 551420 57572 551472
rect 89812 551420 89864 551472
rect 93952 551420 94004 551472
rect 114652 551420 114704 551472
rect 121552 551420 121604 551472
rect 201592 551420 201644 551472
rect 211620 551420 211672 551472
rect 280896 551420 280948 551472
rect 58992 551352 59044 551404
rect 102508 551352 102560 551404
rect 144736 551352 144788 551404
rect 156420 551352 156472 551404
rect 200212 551352 200264 551404
rect 283472 551352 283524 551404
rect 65984 551284 66036 551336
rect 123208 551284 123260 551336
rect 137192 551284 137244 551336
rect 169116 551284 169168 551336
rect 186412 551284 186464 551336
rect 281908 551284 281960 551336
rect 69112 550128 69164 550180
rect 121000 550128 121052 550180
rect 193496 550128 193548 550180
rect 213184 550128 213236 550180
rect 246488 550128 246540 550180
rect 307024 550128 307076 550180
rect 80704 550060 80756 550112
rect 109684 550060 109736 550112
rect 177764 550060 177816 550112
rect 225052 550060 225104 550112
rect 245108 550060 245160 550112
rect 312544 550060 312596 550112
rect 59544 549992 59596 550044
rect 101036 549992 101088 550044
rect 142620 549992 142672 550044
rect 202144 549992 202196 550044
rect 210332 549992 210384 550044
rect 281172 549992 281224 550044
rect 70952 549924 71004 549976
rect 121920 549924 121972 549976
rect 131212 549924 131264 549976
rect 177304 549924 177356 549976
rect 189080 549924 189132 549976
rect 262864 549924 262916 549976
rect 120264 549856 120316 549908
rect 190552 549856 190604 549908
rect 197084 549856 197136 549908
rect 283380 549856 283432 549908
rect 40040 549176 40092 549228
rect 317512 549176 317564 549228
rect 199200 548700 199252 548752
rect 215944 548700 215996 548752
rect 88432 548632 88484 548684
rect 104900 548632 104952 548684
rect 189908 548632 189960 548684
rect 206468 548632 206520 548684
rect 76748 548564 76800 548616
rect 112444 548564 112496 548616
rect 138756 548564 138808 548616
rect 153384 548564 153436 548616
rect 157892 548564 157944 548616
rect 200948 548564 201000 548616
rect 205640 548564 205692 548616
rect 264244 548564 264296 548616
rect 59176 548496 59228 548548
rect 108212 548496 108264 548548
rect 136916 548496 136968 548548
rect 202328 548496 202380 548548
rect 251548 548496 251600 548548
rect 319720 548496 319772 548548
rect 283748 547476 283800 547528
rect 304264 547476 304316 547528
rect 260196 547408 260248 547460
rect 286508 547408 286560 547460
rect 57612 547340 57664 547392
rect 91744 547340 91796 547392
rect 140504 547340 140556 547392
rect 188344 547340 188396 547392
rect 190644 547340 190696 547392
rect 204904 547340 204956 547392
rect 211068 547340 211120 547392
rect 236000 547340 236052 547392
rect 263692 547340 263744 547392
rect 309784 547340 309836 547392
rect 84568 547272 84620 547324
rect 122012 547272 122064 547324
rect 124036 547272 124088 547324
rect 201776 547272 201828 547324
rect 235080 547272 235132 547324
rect 319628 547272 319680 547324
rect 62764 547204 62816 547256
rect 105360 547204 105412 547256
rect 185584 547204 185636 547256
rect 274640 547204 274692 547256
rect 282368 547204 282420 547256
rect 300124 547204 300176 547256
rect 63132 547136 63184 547188
rect 110512 547136 110564 547188
rect 122656 547136 122708 547188
rect 137284 547136 137336 547188
rect 147864 547136 147916 547188
rect 184204 547136 184256 547188
rect 187792 547136 187844 547188
rect 283656 547136 283708 547188
rect 139860 546456 139912 546508
rect 141884 546456 141936 546508
rect 184940 545980 184992 546032
rect 216036 545980 216088 546032
rect 138296 545912 138348 545964
rect 200856 545912 200908 545964
rect 206376 545912 206428 545964
rect 241520 545912 241572 545964
rect 250076 545912 250128 545964
rect 289084 545912 289136 545964
rect 82452 545844 82504 545896
rect 116584 545844 116636 545896
rect 139032 545844 139084 545896
rect 202052 545844 202104 545896
rect 217876 545844 217928 545896
rect 260104 545844 260156 545896
rect 275192 545844 275244 545896
rect 313924 545844 313976 545896
rect 57244 545776 57296 545828
rect 103244 545776 103296 545828
rect 198556 545776 198608 545828
rect 278044 545776 278096 545828
rect 71688 545708 71740 545760
rect 123576 545708 123628 545760
rect 127624 545708 127676 545760
rect 194692 545708 194744 545760
rect 197820 545708 197872 545760
rect 210608 545708 210660 545760
rect 234344 545708 234396 545760
rect 319536 545708 319588 545760
rect 288072 545232 288124 545284
rect 314200 545232 314252 545284
rect 286692 545164 286744 545216
rect 314016 545164 314068 545216
rect 242256 545096 242308 545148
rect 316776 545096 316828 545148
rect 168380 544552 168432 544604
rect 200672 544552 200724 544604
rect 270132 544552 270184 544604
rect 286416 544552 286468 544604
rect 137928 544484 137980 544536
rect 149796 544484 149848 544536
rect 152648 544484 152700 544536
rect 201960 544484 202012 544536
rect 219164 544484 219216 544536
rect 227168 544484 227220 544536
rect 267280 544484 267332 544536
rect 295984 544484 296036 544536
rect 94596 544416 94648 544468
rect 123300 544416 123352 544468
rect 129740 544416 129792 544468
rect 202880 544416 202932 544468
rect 220728 544416 220780 544468
rect 247040 544416 247092 544468
rect 271604 544416 271656 544468
rect 318156 544416 318208 544468
rect 71044 544348 71096 544400
rect 108948 544348 109000 544400
rect 147772 544348 147824 544400
rect 167000 544348 167052 544400
rect 184204 544348 184256 544400
rect 282000 544348 282052 544400
rect 69112 544008 69164 544060
rect 70308 544008 70360 544060
rect 104164 544008 104216 544060
rect 113272 544008 113324 544060
rect 121092 544008 121144 544060
rect 121552 544008 121604 544060
rect 122564 544008 122616 544060
rect 290924 544008 290976 544060
rect 63500 543872 63552 543924
rect 64512 543872 64564 543924
rect 78680 543872 78732 543924
rect 79600 543872 79652 543924
rect 88432 543872 88484 543924
rect 89628 543872 89680 543924
rect 89812 543872 89864 543924
rect 91008 543872 91060 543924
rect 100760 543872 100812 543924
rect 101772 543872 101824 543924
rect 61660 543668 61712 543720
rect 64144 543668 64196 543720
rect 88984 543668 89036 543720
rect 90364 543668 90416 543720
rect 179512 543940 179564 543992
rect 180616 543940 180668 543992
rect 293960 543940 294012 543992
rect 295248 543940 295300 543992
rect 314108 543940 314160 543992
rect 106280 543872 106332 543924
rect 107568 543872 107620 543924
rect 114560 543872 114612 543924
rect 115388 543872 115440 543924
rect 124220 543872 124272 543924
rect 125416 543872 125468 543924
rect 125600 543872 125652 543924
rect 126888 543872 126940 543924
rect 136640 543872 136692 543924
rect 137652 543872 137704 543924
rect 142160 543872 142212 543924
rect 143356 543872 143408 543924
rect 147680 543872 147732 543924
rect 148324 543872 148376 543924
rect 154580 543872 154632 543924
rect 155500 543872 155552 543924
rect 158720 543872 158772 543924
rect 159824 543872 159876 543924
rect 160100 543872 160152 543924
rect 161296 543872 161348 543924
rect 161572 543872 161624 543924
rect 162676 543872 162728 543924
rect 164332 543872 164384 543924
rect 165528 543872 165580 543924
rect 186320 543872 186372 543924
rect 187056 543872 187108 543924
rect 191840 543872 191892 543924
rect 192760 543872 192812 543924
rect 193220 543872 193272 543924
rect 194232 543872 194284 543924
rect 208400 543872 208452 543924
rect 209228 543872 209280 543924
rect 212540 543872 212592 543924
rect 213552 543872 213604 543924
rect 222200 543872 222252 543924
rect 222844 543872 222896 543924
rect 255320 543872 255372 543924
rect 256516 543872 256568 543924
rect 273260 543872 273312 543924
rect 274456 543872 274508 543924
rect 285220 543872 285272 543924
rect 313924 543872 313976 543924
rect 137560 543804 137612 543856
rect 139768 543804 139820 543856
rect 252284 543804 252336 543856
rect 317972 543804 318024 543856
rect 237932 543736 237984 543788
rect 316684 543736 316736 543788
rect 106096 543668 106148 543720
rect 108304 543668 108356 543720
rect 111800 543668 111852 543720
rect 115204 543668 115256 543720
rect 116124 543668 116176 543720
rect 135444 543668 135496 543720
rect 137376 543668 137428 543720
rect 159364 543668 159416 543720
rect 163412 543668 163464 543720
rect 165620 543668 165672 543720
rect 169852 543668 169904 543720
rect 201408 543668 201460 543720
rect 206284 543668 206336 543720
rect 207112 543668 207164 543720
rect 209044 543668 209096 543720
rect 217232 543668 217284 543720
rect 218612 543668 218664 543720
rect 219532 543668 219584 543720
rect 221464 543668 221516 543720
rect 224408 543668 224460 543720
rect 225788 543668 225840 543720
rect 55128 543600 55180 543652
rect 67364 543600 67416 543652
rect 137836 543600 137888 543652
rect 145472 543600 145524 543652
rect 164884 543600 164936 543652
rect 172704 543600 172756 543652
rect 217600 543600 217652 543652
rect 219256 543600 219308 543652
rect 55036 543532 55088 543584
rect 88892 543532 88944 543584
rect 91100 543532 91152 543584
rect 96804 543532 96856 543584
rect 110420 543532 110472 543584
rect 119344 543532 119396 543584
rect 120448 543532 120500 543584
rect 122656 543532 122708 543584
rect 131856 543532 131908 543584
rect 133144 543532 133196 543584
rect 134984 543532 135036 543584
rect 146944 543532 146996 543584
rect 57796 543464 57848 543516
rect 93216 543464 93268 543516
rect 118240 543464 118292 543516
rect 126244 543464 126296 543516
rect 136364 543464 136416 543516
rect 156972 543464 157024 543516
rect 58716 543396 58768 543448
rect 95332 543396 95384 543448
rect 96068 543396 96120 543448
rect 106924 543396 106976 543448
rect 114008 543396 114060 543448
rect 124496 543396 124548 543448
rect 134892 543396 134944 543448
rect 157708 543396 157760 543448
rect 164148 543396 164200 543448
rect 173992 543396 174044 543448
rect 199936 543396 199988 543448
rect 210424 543396 210476 543448
rect 56508 543328 56560 543380
rect 83924 543328 83976 543380
rect 85304 543328 85356 543380
rect 122288 543328 122340 543380
rect 136456 543328 136508 543380
rect 164884 543328 164936 543380
rect 195612 543328 195664 543380
rect 206468 543328 206520 543380
rect 257252 543328 257304 543380
rect 300584 543328 300636 543380
rect 56324 543260 56376 543312
rect 99656 543260 99708 543312
rect 106832 543260 106884 543312
rect 124404 543260 124456 543312
rect 128268 543260 128320 543312
rect 157984 543260 158036 543312
rect 160744 543260 160796 543312
rect 167736 543260 167788 543312
rect 170588 543260 170640 543312
rect 199384 543260 199436 543312
rect 252928 543260 252980 543312
rect 300216 543260 300268 543312
rect 54944 543192 54996 543244
rect 98920 543192 98972 543244
rect 103980 543192 104032 543244
rect 124772 543192 124824 543244
rect 138572 543192 138624 543244
rect 175556 543192 175608 543244
rect 181996 543192 182048 543244
rect 198004 543192 198056 543244
rect 202144 543192 202196 543244
rect 216128 543192 216180 543244
rect 217968 543192 218020 543244
rect 230020 543192 230072 543244
rect 231492 543192 231544 543244
rect 238760 543192 238812 543244
rect 276572 543192 276624 543244
rect 318340 543192 318392 543244
rect 56416 543124 56468 543176
rect 73804 543124 73856 543176
rect 78128 543124 78180 543176
rect 121920 543124 121972 543176
rect 135076 543124 135128 543176
rect 171968 543124 172020 543176
rect 176292 543124 176344 543176
rect 214564 543124 214616 543176
rect 216404 543124 216456 543176
rect 255964 543124 256016 543176
rect 257988 543124 258040 543176
rect 280988 543124 281040 543176
rect 298100 543124 298152 543176
rect 317052 543124 317104 543176
rect 58808 543056 58860 543108
rect 116860 543056 116912 543108
rect 135168 543056 135220 543108
rect 151268 543056 151320 543108
rect 154120 543056 154172 543108
rect 199476 543056 199528 543108
rect 203524 543056 203576 543108
rect 211804 543056 211856 543108
rect 220084 543056 220136 543108
rect 232872 543056 232924 543108
rect 239404 543056 239456 543108
rect 281080 543056 281132 543108
rect 295984 543056 296036 543108
rect 304264 543056 304316 543108
rect 58624 542988 58676 543040
rect 117596 542988 117648 543040
rect 118976 542988 119028 543040
rect 134800 542988 134852 543040
rect 146208 542988 146260 543040
rect 201500 542988 201552 543040
rect 202788 542988 202840 543040
rect 211068 542988 211120 543040
rect 218704 542988 218756 543040
rect 233608 542988 233660 543040
rect 240784 542988 240836 543040
rect 284944 542988 284996 543040
rect 299572 542988 299624 543040
rect 319444 542988 319496 543040
rect 280160 542920 280212 542972
rect 301688 542920 301740 542972
rect 278044 542852 278096 542904
rect 300400 542852 300452 542904
rect 277308 542784 277360 542836
rect 301964 542784 302016 542836
rect 275928 542716 275980 542768
rect 301872 542716 301924 542768
rect 270868 542648 270920 542700
rect 300308 542648 300360 542700
rect 273720 542580 273772 542632
rect 304356 542580 304408 542632
rect 285956 542512 286008 542564
rect 300124 542512 300176 542564
rect 281632 542444 281684 542496
rect 302884 542444 302936 542496
rect 237196 542376 237248 542428
rect 282920 542376 282972 542428
rect 284484 542376 284536 542428
rect 301412 542376 301464 542428
rect 236460 541832 236512 541884
rect 304448 541832 304500 541884
rect 235816 541764 235868 541816
rect 319444 541764 319496 541816
rect 268752 541696 268804 541748
rect 301780 541696 301832 541748
rect 263048 541628 263100 541680
rect 302056 541628 302108 541680
rect 260840 541560 260892 541612
rect 317144 541560 317196 541612
rect 243636 541492 243688 541544
rect 300676 541492 300728 541544
rect 244372 541424 244424 541476
rect 303068 541424 303120 541476
rect 255872 541356 255924 541408
rect 318156 541356 318208 541408
rect 240048 541288 240100 541340
rect 303160 541288 303212 541340
rect 254400 541220 254452 541272
rect 319720 541220 319772 541272
rect 283104 541152 283156 541204
rect 316960 541152 317012 541204
rect 249432 541084 249484 541136
rect 317972 541084 318024 541136
rect 247224 541016 247276 541068
rect 319628 541016 319680 541068
rect 272340 540948 272392 541000
rect 300492 540948 300544 541000
rect 293776 540608 293828 540660
rect 314292 540540 314344 540592
rect 287336 540472 287388 540524
rect 314384 540472 314436 540524
rect 278780 540404 278832 540456
rect 301504 540404 301556 540456
rect 265900 540336 265952 540388
rect 307024 540336 307076 540388
rect 265164 540268 265216 540320
rect 312544 540268 312596 540320
rect 273076 540200 273128 540252
rect 319812 540200 319864 540252
rect 262312 540132 262364 540184
rect 318432 540132 318484 540184
rect 3608 540064 3660 540116
rect 319352 540064 319404 540116
rect 301504 539520 301556 539572
rect 318064 539520 318116 539572
rect 304448 535372 304500 535424
rect 317604 535372 317656 535424
rect 302240 532176 302292 532228
rect 304448 532176 304500 532228
rect 300676 529864 300728 529916
rect 317604 529864 317656 529916
rect 303160 525716 303212 525768
rect 317604 525716 317656 525768
rect 431224 525376 431276 525428
rect 431408 525376 431460 525428
rect 430948 525240 431000 525292
rect 431224 525240 431276 525292
rect 430580 524968 430632 525020
rect 430856 524968 430908 525020
rect 319260 523676 319312 523728
rect 319628 523676 319680 523728
rect 314200 520208 314252 520260
rect 512000 520208 512052 520260
rect 302976 520140 303028 520192
rect 457628 520140 457680 520192
rect 317236 520072 317288 520124
rect 457536 520072 457588 520124
rect 300308 520004 300360 520056
rect 430948 520004 431000 520056
rect 300400 519936 300452 519988
rect 430856 519936 430908 519988
rect 300584 519868 300636 519920
rect 431316 519868 431368 519920
rect 301964 519800 302016 519852
rect 431224 519800 431276 519852
rect 301688 519732 301740 519784
rect 430580 519732 430632 519784
rect 319536 519664 319588 519716
rect 431408 519664 431460 519716
rect 301872 519188 301924 519240
rect 351276 519188 351328 519240
rect 305644 519120 305696 519172
rect 369308 519120 369360 519172
rect 304356 519052 304408 519104
rect 396908 519052 396960 519104
rect 318340 518984 318392 519036
rect 414940 518984 414992 519036
rect 312544 518848 312596 518900
rect 320088 518916 320140 518968
rect 324872 518916 324924 518968
rect 429200 518916 429252 518968
rect 319720 518848 319772 518900
rect 346676 518848 346728 518900
rect 319444 518780 319496 518832
rect 333244 518780 333296 518832
rect 318432 518712 318484 518764
rect 328736 518712 328788 518764
rect 318064 518644 318116 518696
rect 423956 518644 424008 518696
rect 302056 518576 302108 518628
rect 401600 518576 401652 518628
rect 318156 518508 318208 518560
rect 406016 518508 406068 518560
rect 301780 518440 301832 518492
rect 387892 518440 387944 518492
rect 307024 518372 307076 518424
rect 383660 518372 383712 518424
rect 319812 518304 319864 518356
rect 364708 518304 364760 518356
rect 319260 518236 319312 518288
rect 360292 518236 360344 518288
rect 317144 518168 317196 518220
rect 342260 518168 342312 518220
rect 300216 518100 300268 518152
rect 431132 518100 431184 518152
rect 303068 518032 303120 518084
rect 419540 518032 419592 518084
rect 300492 517964 300544 518016
rect 410524 517964 410576 518016
rect 304264 517420 304316 517472
rect 505100 517420 505152 517472
rect 318248 517352 318300 517404
rect 512184 517352 512236 517404
rect 300124 517284 300176 517336
rect 483020 517284 483072 517336
rect 317052 517216 317104 517268
rect 457444 517216 457496 517268
rect 301504 517148 301556 517200
rect 430764 517148 430816 517200
rect 302792 517080 302844 517132
rect 431040 517080 431092 517132
rect 302884 516128 302936 516180
rect 519544 516128 519596 516180
rect 314016 516060 314068 516112
rect 512092 516060 512144 516112
rect 314108 515992 314160 516044
rect 489920 515992 489972 516044
rect 314384 515924 314436 515976
rect 474740 515924 474792 515976
rect 313924 515856 313976 515908
rect 466460 515856 466512 515908
rect 314292 515788 314344 515840
rect 459560 515788 459612 515840
rect 316776 515720 316828 515772
rect 429568 515720 429620 515772
rect 316960 515652 317012 515704
rect 429476 515652 429528 515704
rect 304448 515380 304500 515432
rect 580264 515380 580316 515432
rect 316684 514700 316736 514752
rect 428372 514700 428424 514752
rect 316868 514632 316920 514684
rect 427820 514632 427872 514684
rect 498200 511912 498252 511964
rect 580172 511912 580224 511964
rect 41328 509872 41380 509924
rect 57704 509872 57756 509924
rect 302884 487160 302936 487212
rect 520924 487160 520976 487212
rect 189080 480020 189132 480072
rect 189356 480020 189408 480072
rect 160116 479816 160168 479868
rect 160284 479816 160336 479868
rect 197560 479816 197612 479868
rect 198280 479816 198332 479868
rect 50804 479136 50856 479188
rect 84384 479136 84436 479188
rect 52000 479068 52052 479120
rect 99380 479068 99432 479120
rect 50344 479000 50396 479052
rect 98920 479000 98972 479052
rect 140780 479000 140832 479052
rect 199108 479000 199160 479052
rect 51724 478932 51776 478984
rect 100208 478932 100260 478984
rect 109040 478932 109092 478984
rect 206100 478932 206152 478984
rect 45376 478864 45428 478916
rect 105084 478864 105136 478916
rect 109500 478864 109552 478916
rect 207112 478864 207164 478916
rect 53748 478796 53800 478848
rect 74264 478796 74316 478848
rect 75368 478796 75420 478848
rect 107292 478796 107344 478848
rect 149520 478796 149572 478848
rect 208400 478796 208452 478848
rect 60004 478728 60056 478780
rect 91836 478728 91888 478780
rect 152188 478728 152240 478780
rect 210240 478728 210292 478780
rect 52184 478660 52236 478712
rect 84844 478660 84896 478712
rect 154396 478660 154448 478712
rect 211344 478660 211396 478712
rect 238944 478660 238996 478712
rect 356704 478660 356756 478712
rect 50712 478592 50764 478644
rect 68928 478592 68980 478644
rect 71320 478592 71372 478644
rect 106372 478592 106424 478644
rect 153108 478592 153160 478644
rect 205640 478592 205692 478644
rect 239864 478592 239916 478644
rect 362316 478592 362368 478644
rect 68284 478524 68336 478576
rect 104624 478524 104676 478576
rect 149152 478524 149204 478576
rect 200764 478524 200816 478576
rect 240232 478524 240284 478576
rect 365168 478524 365220 478576
rect 68376 478456 68428 478508
rect 105544 478456 105596 478508
rect 151268 478456 151320 478508
rect 201592 478456 201644 478508
rect 232320 478456 232372 478508
rect 360844 478456 360896 478508
rect 54760 478388 54812 478440
rect 102416 478388 102468 478440
rect 157892 478388 157944 478440
rect 205640 478388 205692 478440
rect 235448 478388 235500 478440
rect 366456 478388 366508 478440
rect 48044 478320 48096 478372
rect 97540 478320 97592 478372
rect 153476 478320 153528 478372
rect 200488 478320 200540 478372
rect 209412 478320 209464 478372
rect 216680 478320 216732 478372
rect 224408 478320 224460 478372
rect 358176 478320 358228 478372
rect 51908 478252 51960 478304
rect 99748 478252 99800 478304
rect 138940 478252 138992 478304
rect 193864 478252 193916 478304
rect 209596 478252 209648 478304
rect 221740 478252 221792 478304
rect 230572 478252 230624 478304
rect 366364 478252 366416 478304
rect 47952 478184 48004 478236
rect 97172 478184 97224 478236
rect 109868 478184 109920 478236
rect 169024 478184 169076 478236
rect 200212 478184 200264 478236
rect 212264 478184 212316 478236
rect 225328 478184 225380 478236
rect 362224 478184 362276 478236
rect 55128 478116 55180 478168
rect 89628 478116 89680 478168
rect 95332 478116 95384 478168
rect 182824 478116 182876 478168
rect 186504 478116 186556 478168
rect 198188 478116 198240 478168
rect 201960 478116 202012 478168
rect 217324 478116 217376 478168
rect 225696 478116 225748 478168
rect 373264 478116 373316 478168
rect 64144 478048 64196 478100
rect 69664 478048 69716 478100
rect 75276 478048 75328 478100
rect 102876 478048 102928 478100
rect 150440 478048 150492 478100
rect 197452 478048 197504 478100
rect 56508 477980 56560 478032
rect 81716 477980 81768 478032
rect 156604 477980 156656 478032
rect 197360 477980 197412 478032
rect 50896 477912 50948 477964
rect 75828 477912 75880 477964
rect 139400 477912 139452 477964
rect 178592 477912 178644 477964
rect 58440 477844 58492 477896
rect 81256 477844 81308 477896
rect 168932 477844 168984 477896
rect 206376 477844 206428 477896
rect 194876 477572 194928 477624
rect 196992 477572 197044 477624
rect 202420 477572 202472 477624
rect 209504 477572 209556 477624
rect 195796 477504 195848 477556
rect 196900 477504 196952 477556
rect 208584 477504 208636 477556
rect 210792 477504 210844 477556
rect 211160 477504 211212 477556
rect 214564 477504 214616 477556
rect 220176 477504 220228 477556
rect 222660 477504 222712 477556
rect 297088 477368 297140 477420
rect 372528 477368 372580 477420
rect 290924 477300 290976 477352
rect 365628 477300 365680 477352
rect 283012 477232 283064 477284
rect 359740 477232 359792 477284
rect 282552 477164 282604 477216
rect 363512 477164 363564 477216
rect 261852 477096 261904 477148
rect 374184 477096 374236 477148
rect 256608 477028 256660 477080
rect 376392 477028 376444 477080
rect 242900 476960 242952 477012
rect 368020 476960 368072 477012
rect 45468 476892 45520 476944
rect 117872 476892 117924 476944
rect 177764 476892 177816 476944
rect 211988 476892 212040 476944
rect 247316 476892 247368 476944
rect 374736 476892 374788 476944
rect 60556 476824 60608 476876
rect 120724 476824 120776 476876
rect 3608 476756 3660 476808
rect 159640 476824 159692 476876
rect 218704 476824 218756 476876
rect 236736 476824 236788 476876
rect 364984 476824 365036 476876
rect 429384 476756 429436 476808
rect 120724 476688 120776 476740
rect 133144 476620 133196 476672
rect 70400 476076 70452 476128
rect 70860 476076 70912 476128
rect 85764 476076 85816 476128
rect 85948 476076 86000 476128
rect 47768 476008 47820 476060
rect 111708 476008 111760 476060
rect 46664 475940 46716 475992
rect 111248 475940 111300 475992
rect 294052 475940 294104 475992
rect 294236 475940 294288 475992
rect 49240 475872 49292 475924
rect 115204 475872 115256 475924
rect 274732 475872 274784 475924
rect 274916 475872 274968 475924
rect 291844 475872 291896 475924
rect 373908 475872 373960 475924
rect 46388 475804 46440 475856
rect 112536 475804 112588 475856
rect 267556 475804 267608 475856
rect 359464 475804 359516 475856
rect 46480 475736 46532 475788
rect 112076 475736 112128 475788
rect 267096 475736 267148 475788
rect 359556 475736 359608 475788
rect 50252 475668 50304 475720
rect 116032 475668 116084 475720
rect 136364 475668 136416 475720
rect 141884 475668 141936 475720
rect 171140 475668 171192 475720
rect 171324 475668 171376 475720
rect 184296 475668 184348 475720
rect 216128 475668 216180 475720
rect 273260 475668 273312 475720
rect 369768 475668 369820 475720
rect 48136 475600 48188 475652
rect 115664 475600 115716 475652
rect 138112 475600 138164 475652
rect 200488 475600 200540 475652
rect 219532 475600 219584 475652
rect 272892 475600 272944 475652
rect 372436 475600 372488 475652
rect 47860 475532 47912 475584
rect 119620 475532 119672 475584
rect 136732 475532 136784 475584
rect 199384 475532 199436 475584
rect 57152 475464 57204 475516
rect 132408 475464 132460 475516
rect 137652 475464 137704 475516
rect 57336 475396 57388 475448
rect 135904 475396 135956 475448
rect 140780 475396 140832 475448
rect 141700 475396 141752 475448
rect 141884 475464 141936 475516
rect 201684 475464 201736 475516
rect 204444 475396 204496 475448
rect 62120 475328 62172 475380
rect 62948 475328 63000 475380
rect 63500 475328 63552 475380
rect 64236 475328 64288 475380
rect 64328 475328 64380 475380
rect 49148 475260 49200 475312
rect 98000 475260 98052 475312
rect 100852 475260 100904 475312
rect 101220 475260 101272 475312
rect 103612 475260 103664 475312
rect 103796 475260 103848 475312
rect 107660 475260 107712 475312
rect 107844 475260 107896 475312
rect 133972 475260 134024 475312
rect 134708 475260 134760 475312
rect 139400 475260 139452 475312
rect 140044 475260 140096 475312
rect 140872 475260 140924 475312
rect 141332 475260 141384 475312
rect 142252 475260 142304 475312
rect 142620 475260 142672 475312
rect 143540 475260 143592 475312
rect 143908 475260 143960 475312
rect 150440 475260 150492 475312
rect 151452 475260 151504 475312
rect 160100 475260 160152 475312
rect 160652 475260 160704 475312
rect 161572 475260 161624 475312
rect 161940 475260 161992 475312
rect 165620 475260 165672 475312
rect 166356 475260 166408 475312
rect 167000 475260 167052 475312
rect 167736 475260 167788 475312
rect 178132 475260 178184 475312
rect 178684 475260 178736 475312
rect 179420 475260 179472 475312
rect 180064 475260 180116 475312
rect 180892 475260 180944 475312
rect 181444 475260 181496 475312
rect 182364 475260 182416 475312
rect 182732 475260 182784 475312
rect 183560 475260 183612 475312
rect 184388 475260 184440 475312
rect 185032 475260 185084 475312
rect 185860 475260 185912 475312
rect 51816 475192 51868 475244
rect 98460 475192 98512 475244
rect 100760 475192 100812 475244
rect 101588 475192 101640 475244
rect 142160 475192 142212 475244
rect 142988 475192 143040 475244
rect 161480 475192 161532 475244
rect 161756 475192 161808 475244
rect 180800 475192 180852 475244
rect 181076 475192 181128 475244
rect 182180 475192 182232 475244
rect 182548 475192 182600 475244
rect 205732 475328 205784 475380
rect 206468 475328 206520 475380
rect 207204 475328 207256 475380
rect 207756 475328 207808 475380
rect 209780 475328 209832 475380
rect 209964 475328 210016 475380
rect 212540 475464 212592 475516
rect 253020 475532 253072 475584
rect 365444 475532 365496 475584
rect 243360 475464 243412 475516
rect 369216 475464 369268 475516
rect 219532 475396 219584 475448
rect 247776 475396 247828 475448
rect 376208 475396 376260 475448
rect 212540 475328 212592 475380
rect 213092 475328 213144 475380
rect 213920 475328 213972 475380
rect 214932 475328 214984 475380
rect 215300 475328 215352 475380
rect 216220 475328 216272 475380
rect 218060 475328 218112 475380
rect 218796 475328 218848 475380
rect 222200 475328 222252 475380
rect 374644 475328 374696 475380
rect 212724 475260 212776 475312
rect 244280 475260 244332 475312
rect 244556 475260 244608 475312
rect 245660 475260 245712 475312
rect 246580 475260 246632 475312
rect 248512 475260 248564 475312
rect 249156 475260 249208 475312
rect 251180 475260 251232 475312
rect 251364 475260 251416 475312
rect 252560 475260 252612 475312
rect 253204 475260 253256 475312
rect 259460 475260 259512 475312
rect 260196 475260 260248 475312
rect 262220 475260 262272 475312
rect 262404 475260 262456 475312
rect 276112 475260 276164 475312
rect 276572 475260 276624 475312
rect 277492 475260 277544 475312
rect 277860 475260 277912 475312
rect 284300 475260 284352 475312
rect 284852 475260 284904 475312
rect 285680 475260 285732 475312
rect 286692 475260 286744 475312
rect 291200 475260 291252 475312
rect 291936 475260 291988 475312
rect 296720 475260 296772 475312
rect 297732 475260 297784 475312
rect 199200 475192 199252 475244
rect 276020 475192 276072 475244
rect 276940 475192 276992 475244
rect 277400 475192 277452 475244
rect 278228 475192 278280 475244
rect 54668 475124 54720 475176
rect 96712 475124 96764 475176
rect 182272 475124 182324 475176
rect 183100 475124 183152 475176
rect 205640 475124 205692 475176
rect 205916 475124 205968 475176
rect 62764 475056 62816 475108
rect 64328 475056 64380 475108
rect 64972 475056 65024 475108
rect 65524 475056 65576 475108
rect 66260 475056 66312 475108
rect 66812 475056 66864 475108
rect 71872 475056 71924 475108
rect 72608 475056 72660 475108
rect 78680 475056 78732 475108
rect 79692 475056 79744 475108
rect 82820 475056 82872 475108
rect 83556 475056 83608 475108
rect 85672 475056 85724 475108
rect 86316 475056 86368 475108
rect 87052 475056 87104 475108
rect 87236 475056 87288 475108
rect 88432 475056 88484 475108
rect 88892 475056 88944 475108
rect 89812 475056 89864 475108
rect 90732 475056 90784 475108
rect 92480 475056 92532 475108
rect 92940 475056 92992 475108
rect 86960 474988 87012 475040
rect 87604 474988 87656 475040
rect 88524 474988 88576 475040
rect 88708 474988 88760 475040
rect 92572 474988 92624 475040
rect 93308 474988 93360 475040
rect 293592 474648 293644 474700
rect 379336 474648 379388 474700
rect 282092 474580 282144 474632
rect 379980 474580 380032 474632
rect 275928 474512 275980 474564
rect 373724 474512 373776 474564
rect 260932 474444 260984 474496
rect 362500 474444 362552 474496
rect 254768 474376 254820 474428
rect 366824 474376 366876 474428
rect 255228 474308 255280 474360
rect 369124 474308 369176 474360
rect 252192 474240 252244 474292
rect 366916 474240 366968 474292
rect 242440 474172 242492 474224
rect 370596 474172 370648 474224
rect 204996 474104 205048 474156
rect 217324 474104 217376 474156
rect 228824 474104 228876 474156
rect 363604 474104 363656 474156
rect 58808 473968 58860 474020
rect 96252 474036 96304 474088
rect 176016 474036 176068 474088
rect 210608 474036 210660 474088
rect 238116 474036 238168 474088
rect 376300 474036 376352 474088
rect 166264 473968 166316 474020
rect 215944 473968 215996 474020
rect 228364 473968 228416 474020
rect 367836 473968 367888 474020
rect 295340 473900 295392 473952
rect 375472 473900 375524 473952
rect 81532 473560 81584 473612
rect 82268 473560 82320 473612
rect 46848 473288 46900 473340
rect 116492 473288 116544 473340
rect 58624 473220 58676 473272
rect 130568 473220 130620 473272
rect 59728 473152 59780 473204
rect 132592 473152 132644 473204
rect 43996 473084 44048 473136
rect 118240 473084 118292 473136
rect 298560 473084 298612 473136
rect 374000 473084 374052 473136
rect 49056 473016 49108 473068
rect 131028 473016 131080 473068
rect 275468 473016 275520 473068
rect 356888 473016 356940 473068
rect 50160 472948 50212 473000
rect 131488 472948 131540 473000
rect 295800 472948 295852 473000
rect 377772 472948 377824 473000
rect 52276 472880 52328 472932
rect 134156 472880 134208 472932
rect 279240 472880 279292 472932
rect 364892 472880 364944 472932
rect 47584 472812 47636 472864
rect 129740 472812 129792 472864
rect 280804 472812 280856 472864
rect 369676 472812 369728 472864
rect 46112 472744 46164 472796
rect 129280 472744 129332 472796
rect 258816 472744 258868 472796
rect 372252 472744 372304 472796
rect 42340 472676 42392 472728
rect 131948 472676 132000 472728
rect 238484 472676 238536 472728
rect 358084 472676 358136 472728
rect 43260 472608 43312 472660
rect 132500 472608 132552 472660
rect 175556 472608 175608 472660
rect 213184 472608 213236 472660
rect 239404 472608 239456 472660
rect 378784 472608 378836 472660
rect 47676 472540 47728 472592
rect 116952 472540 117004 472592
rect 54576 472472 54628 472524
rect 117412 472472 117464 472524
rect 172520 472472 172572 472524
rect 173532 472472 173584 472524
rect 57888 472404 57940 472456
rect 114284 472404 114336 472456
rect 296168 471928 296220 471980
rect 373816 471928 373868 471980
rect 288716 471860 288768 471912
rect 375196 471860 375248 471912
rect 270684 471792 270736 471844
rect 358452 471792 358504 471844
rect 272432 471724 272484 471776
rect 360752 471724 360804 471776
rect 266268 471656 266320 471708
rect 356796 471656 356848 471708
rect 265808 471588 265860 471640
rect 361028 471588 361080 471640
rect 257436 471520 257488 471572
rect 358360 471520 358412 471572
rect 259644 471452 259696 471504
rect 369492 471452 369544 471504
rect 253940 471384 253992 471436
rect 369584 471384 369636 471436
rect 193220 471316 193272 471368
rect 194140 471316 194192 471368
rect 198740 471316 198792 471368
rect 199016 471316 199068 471368
rect 244464 471316 244516 471368
rect 371976 471316 372028 471368
rect 57704 471248 57756 471300
rect 113916 471248 113968 471300
rect 169392 471248 169444 471300
rect 207664 471248 207716 471300
rect 226800 471248 226852 471300
rect 376116 471248 376168 471300
rect 190460 471180 190512 471232
rect 190644 471180 190696 471232
rect 191840 471180 191892 471232
rect 192852 471180 192904 471232
rect 193312 471180 193364 471232
rect 193772 471180 193824 471232
rect 198832 471180 198884 471232
rect 199476 471180 199528 471232
rect 202880 471180 202932 471232
rect 203156 471180 203208 471232
rect 204352 471180 204404 471232
rect 205180 471180 205232 471232
rect 267740 471180 267792 471232
rect 268108 471180 268160 471232
rect 203156 471044 203208 471096
rect 203892 471044 203944 471096
rect 43628 470500 43680 470552
rect 120172 470500 120224 470552
rect 43812 470432 43864 470484
rect 121736 470432 121788 470484
rect 56048 470364 56100 470416
rect 133972 470364 134024 470416
rect 42708 470296 42760 470348
rect 121920 470296 121972 470348
rect 278872 470296 278924 470348
rect 356980 470296 357032 470348
rect 45192 470228 45244 470280
rect 124956 470228 125008 470280
rect 285956 470228 286008 470280
rect 379152 470228 379204 470280
rect 43536 470160 43588 470212
rect 122840 470160 122892 470212
rect 269948 470160 270000 470212
rect 371792 470160 371844 470212
rect 43720 470092 43772 470144
rect 124496 470092 124548 470144
rect 258172 470092 258224 470144
rect 364064 470092 364116 470144
rect 42248 470024 42300 470076
rect 123668 470024 123720 470076
rect 252652 470024 252704 470076
rect 376484 470024 376536 470076
rect 42524 469956 42576 470008
rect 124220 469956 124272 470008
rect 187148 469956 187200 470008
rect 209228 469956 209280 470008
rect 245844 469956 245896 470008
rect 370688 469956 370740 470008
rect 48964 469888 49016 469940
rect 132684 469888 132736 469940
rect 176752 469888 176804 469940
rect 204996 469888 205048 469940
rect 205916 469888 205968 469940
rect 217600 469888 217652 469940
rect 242900 469888 242952 469940
rect 374828 469888 374880 469940
rect 44732 469820 44784 469872
rect 143632 469820 143684 469872
rect 165712 469820 165764 469872
rect 211804 469820 211856 469872
rect 229192 469820 229244 469872
rect 367928 469820 367980 469872
rect 53656 469752 53708 469804
rect 127164 469752 127216 469804
rect 57060 469684 57112 469736
rect 128452 469684 128504 469736
rect 58532 469616 58584 469668
rect 128544 469616 128596 469668
rect 40960 469072 41012 469124
rect 62120 469072 62172 469124
rect 289912 469072 289964 469124
rect 362684 469072 362736 469124
rect 40868 469004 40920 469056
rect 62212 469004 62264 469056
rect 274732 469004 274784 469056
rect 363420 469004 363472 469056
rect 45100 468936 45152 468988
rect 71044 468936 71096 468988
rect 178224 468936 178276 468988
rect 202328 468936 202380 468988
rect 271236 468936 271288 468988
rect 361304 468936 361356 468988
rect 44088 468868 44140 468920
rect 70584 468868 70636 468920
rect 178684 468868 178736 468920
rect 205916 468868 205968 468920
rect 273352 468868 273404 468920
rect 368388 468868 368440 468920
rect 46572 468800 46624 468852
rect 75276 468800 75328 468852
rect 161756 468800 161808 468852
rect 210424 468800 210476 468852
rect 263784 468800 263836 468852
rect 362592 468800 362644 468852
rect 41052 468732 41104 468784
rect 93952 468732 94004 468784
rect 162952 468732 163004 468784
rect 216036 468732 216088 468784
rect 262404 468732 262456 468784
rect 368204 468732 368256 468784
rect 45008 468664 45060 468716
rect 104992 468664 105044 468716
rect 139492 468664 139544 468716
rect 207480 468664 207532 468716
rect 259552 468664 259604 468716
rect 370872 468664 370924 468716
rect 44916 468596 44968 468648
rect 106372 468596 106424 468648
rect 127716 468596 127768 468648
rect 197636 468596 197688 468648
rect 245752 468596 245804 468648
rect 365260 468596 365312 468648
rect 59360 468528 59412 468580
rect 179604 468528 179656 468580
rect 187884 468528 187936 468580
rect 209412 468528 209464 468580
rect 241612 468528 241664 468580
rect 366548 468528 366600 468580
rect 15844 468460 15896 468512
rect 378140 468460 378192 468512
rect 285864 467712 285916 467764
rect 357072 467712 357124 467764
rect 294144 467644 294196 467696
rect 376576 467644 376628 467696
rect 265072 467576 265124 467628
rect 365536 467576 365588 467628
rect 269212 467508 269264 467560
rect 375932 467508 375984 467560
rect 268660 467440 268712 467492
rect 375288 467440 375340 467492
rect 253940 467372 253992 467424
rect 364156 467372 364208 467424
rect 187976 467304 188028 467356
rect 200764 467304 200816 467356
rect 207296 467304 207348 467356
rect 217692 467304 217744 467356
rect 258080 467304 258132 467356
rect 373448 467304 373500 467356
rect 185124 467236 185176 467288
rect 214656 467236 214708 467288
rect 244464 467236 244516 467288
rect 360936 467236 360988 467288
rect 176660 467168 176712 467220
rect 207848 467168 207900 467220
rect 237380 467168 237432 467220
rect 358268 467168 358320 467220
rect 57520 467100 57572 467152
rect 114744 467100 114796 467152
rect 171416 467100 171468 467152
rect 209044 467100 209096 467152
rect 227720 467100 227772 467152
rect 370504 467100 370556 467152
rect 44824 466352 44876 466404
rect 68376 466352 68428 466404
rect 182456 466352 182508 466404
rect 206560 466352 206612 466404
rect 52092 466284 52144 466336
rect 82820 466284 82872 466336
rect 190644 466284 190696 466336
rect 214840 466284 214892 466336
rect 50528 466216 50580 466268
rect 82912 466216 82964 466268
rect 191932 466216 191984 466268
rect 216312 466216 216364 466268
rect 289820 466216 289872 466268
rect 361396 466216 361448 466268
rect 42432 466148 42484 466200
rect 75184 466148 75236 466200
rect 182364 466148 182416 466200
rect 207940 466148 207992 466200
rect 299480 466148 299532 466200
rect 371240 466148 371292 466200
rect 48228 466080 48280 466132
rect 81532 466080 81584 466132
rect 174084 466080 174136 466132
rect 200856 466080 200908 466132
rect 296812 466080 296864 466132
rect 369032 466080 369084 466132
rect 49424 466012 49476 466064
rect 83004 466012 83056 466064
rect 192024 466012 192076 466064
rect 219164 466012 219216 466064
rect 298192 466012 298244 466064
rect 373172 466012 373224 466064
rect 59820 465944 59872 465996
rect 102232 465944 102284 465996
rect 139400 465944 139452 465996
rect 197084 465944 197136 465996
rect 288532 465944 288584 465996
rect 371056 465944 371108 465996
rect 57244 465876 57296 465928
rect 103612 465876 103664 465928
rect 140964 465876 141016 465928
rect 200580 465876 200632 465928
rect 240232 465876 240284 465928
rect 366640 465876 366692 465928
rect 53196 465808 53248 465860
rect 100852 465808 100904 465860
rect 140780 465808 140832 465860
rect 201776 465808 201828 465860
rect 241520 465808 241572 465860
rect 369308 465808 369360 465860
rect 58716 465740 58768 465792
rect 110604 465740 110656 465792
rect 140872 465740 140924 465792
rect 204536 465740 204588 465792
rect 226340 465740 226392 465792
rect 363696 465740 363748 465792
rect 53104 465672 53156 465724
rect 100944 465672 100996 465724
rect 107844 465672 107896 465724
rect 202972 465672 203024 465724
rect 226432 465672 226484 465724
rect 371884 465672 371936 465724
rect 40776 465604 40828 465656
rect 60832 465604 60884 465656
rect 183652 465604 183704 465656
rect 205180 465604 205232 465656
rect 46296 465536 46348 465588
rect 64972 465536 65024 465588
rect 182272 465536 182324 465588
rect 202420 465536 202472 465588
rect 47492 465468 47544 465520
rect 65064 465468 65116 465520
rect 192116 465468 192168 465520
rect 208032 465468 208084 465520
rect 294052 464856 294104 464908
rect 358544 464856 358596 464908
rect 292672 464788 292724 464840
rect 367652 464788 367704 464840
rect 283012 464720 283064 464772
rect 357992 464720 358044 464772
rect 284392 464652 284444 464704
rect 359924 464652 359976 464704
rect 284484 464584 284536 464636
rect 360568 464584 360620 464636
rect 293960 464516 294012 464568
rect 377864 464516 377916 464568
rect 291292 464448 291344 464500
rect 378048 464448 378100 464500
rect 285772 464380 285824 464432
rect 377496 464380 377548 464432
rect 57612 464312 57664 464364
rect 111984 464312 112036 464364
rect 158720 464312 158772 464364
rect 203524 464312 203576 464364
rect 284300 464312 284352 464364
rect 377404 464312 377456 464364
rect 55864 463632 55916 463684
rect 87144 463632 87196 463684
rect 185032 463632 185084 463684
rect 212080 463632 212132 463684
rect 282920 463632 282972 463684
rect 359832 463632 359884 463684
rect 55036 463564 55088 463616
rect 86960 463564 87012 463616
rect 190460 463564 190512 463616
rect 217508 463564 217560 463616
rect 277584 463564 277636 463616
rect 360660 463564 360712 463616
rect 48872 463496 48924 463548
rect 81624 463496 81676 463548
rect 186320 463496 186372 463548
rect 213460 463496 213512 463548
rect 276204 463496 276256 463548
rect 364800 463496 364852 463548
rect 56232 463428 56284 463480
rect 88432 463428 88484 463480
rect 180984 463428 181036 463480
rect 210700 463428 210752 463480
rect 277400 463428 277452 463480
rect 367560 463428 367612 463480
rect 56140 463360 56192 463412
rect 88616 463360 88668 463412
rect 180892 463360 180944 463412
rect 212172 463360 212224 463412
rect 273260 463360 273312 463412
rect 366180 463360 366232 463412
rect 52920 463292 52972 463344
rect 85672 463292 85724 463344
rect 175280 463292 175332 463344
rect 206652 463292 206704 463344
rect 267832 463292 267884 463344
rect 362868 463292 362920 463344
rect 56416 463224 56468 463276
rect 89720 463224 89772 463276
rect 168380 463224 168432 463276
rect 209136 463224 209188 463276
rect 274640 463224 274692 463276
rect 370412 463224 370464 463276
rect 54852 463156 54904 463208
rect 88524 463156 88576 463208
rect 160100 463156 160152 463208
rect 202144 463156 202196 463208
rect 267740 463156 267792 463208
rect 367008 463156 367060 463208
rect 57428 463088 57480 463140
rect 113364 463088 113416 463140
rect 142344 463088 142396 463140
rect 208492 463088 208544 463140
rect 249984 463088 250036 463140
rect 370780 463088 370832 463140
rect 53288 463020 53340 463072
rect 87052 463020 87104 463072
rect 109040 463020 109092 463072
rect 200396 463020 200448 463072
rect 248604 463020 248656 463072
rect 372068 463020 372120 463072
rect 53380 462952 53432 463004
rect 92572 462952 92624 463004
rect 107660 462952 107712 463004
rect 200304 462952 200356 463004
rect 240140 462952 240192 463004
rect 363788 462952 363840 463004
rect 54944 462884 54996 462936
rect 85580 462884 85632 462936
rect 190552 462884 190604 462936
rect 203800 462884 203852 462936
rect 40592 462816 40644 462868
rect 60740 462816 60792 462868
rect 189264 462816 189316 462868
rect 199384 462816 199436 462868
rect 46204 462748 46256 462800
rect 64880 462748 64932 462800
rect 193404 462544 193456 462596
rect 202512 462544 202564 462596
rect 133144 462272 133196 462324
rect 178316 462272 178368 462324
rect 287152 462204 287204 462256
rect 362776 462204 362828 462256
rect 298100 462136 298152 462188
rect 375748 462136 375800 462188
rect 280160 462068 280212 462120
rect 363328 462068 363380 462120
rect 260840 462000 260892 462052
rect 361120 462000 361172 462052
rect 269120 461932 269172 461984
rect 370320 461932 370372 461984
rect 191840 461864 191892 461916
rect 205364 461864 205416 461916
rect 263600 461864 263652 461916
rect 372344 461864 372396 461916
rect 511264 461864 511316 461916
rect 517520 461864 517572 461916
rect 182180 461796 182232 461848
rect 203616 461796 203668 461848
rect 264980 461796 265032 461848
rect 375104 461796 375156 461848
rect 179604 461728 179656 461780
rect 201592 461728 201644 461780
rect 262312 461728 262364 461780
rect 373540 461728 373592 461780
rect 179512 461660 179564 461712
rect 206744 461660 206796 461712
rect 251272 461660 251324 461712
rect 365352 461660 365404 461712
rect 161572 461592 161624 461644
rect 213276 461592 213328 461644
rect 252560 461592 252612 461644
rect 375012 461592 375064 461644
rect 178316 461048 178368 461100
rect 210056 461048 210108 461100
rect 338304 461048 338356 461100
rect 357440 461048 357492 461100
rect 498384 461048 498436 461100
rect 201592 460980 201644 461032
rect 339776 460980 339828 461032
rect 358820 460980 358872 461032
rect 499856 460980 499908 461032
rect 517612 460980 517664 461032
rect 190920 460912 190972 460964
rect 207020 460912 207072 460964
rect 210056 460912 210108 460964
rect 338304 460912 338356 460964
rect 351000 460912 351052 460964
rect 367744 460912 367796 460964
rect 498384 460912 498436 460964
rect 517704 460912 517756 460964
rect 48688 460844 48740 460896
rect 78772 460844 78824 460896
rect 157340 460844 157392 460896
rect 218336 460844 218388 460896
rect 285680 460844 285732 460896
rect 377128 460844 377180 460896
rect 53380 460776 53432 460828
rect 78680 460776 78732 460828
rect 193864 460776 193916 460828
rect 203340 460776 203392 460828
rect 287060 460776 287112 460828
rect 379428 460776 379480 460828
rect 51632 460708 51684 460760
rect 76104 460708 76156 460760
rect 189172 460708 189224 460760
rect 202604 460708 202656 460760
rect 266360 460708 266412 460760
rect 368296 460708 368348 460760
rect 52368 460640 52420 460692
rect 76012 460640 76064 460692
rect 193312 460640 193364 460692
rect 208860 460640 208912 460692
rect 259460 460640 259512 460692
rect 370964 460640 371016 460692
rect 55956 460572 56008 460624
rect 77300 460572 77352 460624
rect 189080 460572 189132 460624
rect 210332 460572 210384 460624
rect 249892 460572 249944 460624
rect 362408 460572 362460 460624
rect 51540 460504 51592 460556
rect 66352 460504 66404 460556
rect 169024 460504 169076 460556
rect 197728 460504 197780 460556
rect 251180 460504 251232 460556
rect 363972 460504 364024 460556
rect 47400 460436 47452 460488
rect 63500 460436 63552 460488
rect 184940 460436 184992 460488
rect 216220 460436 216272 460488
rect 249800 460436 249852 460488
rect 368112 460436 368164 460488
rect 49608 460368 49660 460420
rect 70400 460368 70452 460420
rect 179420 460368 179472 460420
rect 214748 460368 214800 460420
rect 248420 460368 248472 460420
rect 369400 460368 369452 460420
rect 41144 460300 41196 460352
rect 71872 460300 71924 460352
rect 178132 460300 178184 460352
rect 213552 460300 213604 460352
rect 244372 460300 244424 460352
rect 366732 460300 366784 460352
rect 41236 460232 41288 460284
rect 74540 460232 74592 460284
rect 164332 460232 164384 460284
rect 218980 460232 219032 460284
rect 248512 460232 248564 460284
rect 373356 460232 373408 460284
rect 43352 460164 43404 460216
rect 68284 460164 68336 460216
rect 69664 460164 69716 460216
rect 199016 460164 199068 460216
rect 247040 460164 247092 460216
rect 378876 460164 378928 460216
rect 54484 460096 54536 460148
rect 63592 460096 63644 460148
rect 278780 460096 278832 460148
rect 362132 460096 362184 460148
rect 291200 460028 291252 460080
rect 374460 460028 374512 460080
rect 288440 459960 288492 460012
rect 357164 459960 357216 460012
rect 215208 459620 215260 459672
rect 221004 459620 221056 459672
rect 216588 459552 216640 459604
rect 220912 459552 220964 459604
rect 187700 459484 187752 459536
rect 200948 459484 201000 459536
rect 295340 459484 295392 459536
rect 370228 459484 370280 459536
rect 193220 459416 193272 459468
rect 211620 459416 211672 459468
rect 281540 459416 281592 459468
rect 359648 459416 359700 459468
rect 178040 459348 178092 459400
rect 203708 459348 203760 459400
rect 276020 459348 276072 459400
rect 358636 459348 358688 459400
rect 58900 459280 58952 459332
rect 92480 459280 92532 459332
rect 180800 459280 180852 459332
rect 209320 459280 209372 459332
rect 271880 459280 271932 459332
rect 358728 459280 358780 459332
rect 55772 459212 55824 459264
rect 103704 459212 103756 459264
rect 173900 459212 173952 459264
rect 205272 459212 205324 459264
rect 256792 459212 256844 459264
rect 361212 459212 361264 459264
rect 51632 459144 51684 459196
rect 99472 459144 99524 459196
rect 173992 459144 174044 459196
rect 219072 459144 219124 459196
rect 262220 459144 262272 459196
rect 378968 459144 379020 459196
rect 53012 459076 53064 459128
rect 100760 459076 100812 459128
rect 142252 459076 142304 459128
rect 197912 459076 197964 459128
rect 256700 459076 256752 459128
rect 373632 459076 373684 459128
rect 57796 459008 57848 459060
rect 118884 459008 118936 459060
rect 142160 459008 142212 459060
rect 199568 459008 199620 459060
rect 244280 459008 244332 459060
rect 363880 459008 363932 459060
rect 54392 458940 54444 458992
rect 121460 458940 121512 458992
rect 135444 458940 135496 458992
rect 197820 458940 197872 458992
rect 245660 458940 245712 458992
rect 379060 458940 379112 458992
rect 55956 458872 56008 458924
rect 130016 458872 130068 458924
rect 136640 458872 136692 458924
rect 199292 458872 199344 458924
rect 236000 458872 236052 458924
rect 372160 458872 372212 458924
rect 54300 458804 54352 458856
rect 134064 458804 134116 458856
rect 138020 458804 138072 458856
rect 200672 458804 200724 458856
rect 223580 458804 223632 458856
rect 365076 458804 365128 458856
rect 194600 458736 194652 458788
rect 206192 458736 206244 458788
rect 292580 458736 292632 458788
rect 366272 458736 366324 458788
rect 59268 458600 59320 458652
rect 66260 458600 66312 458652
rect 199016 458328 199068 458380
rect 48780 458260 48832 458312
rect 358912 458260 358964 458312
rect 516600 458260 516652 458312
rect 207388 458192 207440 458244
rect 208124 458192 208176 458244
rect 205824 457444 205876 457496
rect 217876 457444 217928 457496
rect 55864 457240 55916 457292
rect 56416 457240 56468 457292
rect 48872 456084 48924 456136
rect 49332 456084 49384 456136
rect 52920 456084 52972 456136
rect 53288 456084 53340 456136
rect 519544 454656 519596 454708
rect 580264 454656 580316 454708
rect 208124 417392 208176 417444
rect 217784 417392 217836 417444
rect 203248 413924 203300 413976
rect 206284 413924 206336 413976
rect 48872 412564 48924 412616
rect 56968 412564 57020 412616
rect 2964 411204 3016 411256
rect 15844 411204 15896 411256
rect 44640 409844 44692 409896
rect 57060 409844 57112 409896
rect 205732 409096 205784 409148
rect 216772 409096 216824 409148
rect 360568 409096 360620 409148
rect 377036 409096 377088 409148
rect 55680 408552 55732 408604
rect 56968 408552 57020 408604
rect 46020 408484 46072 408536
rect 57060 408484 57112 408536
rect 359924 407736 359976 407788
rect 376760 407736 376812 407788
rect 376944 407736 376996 407788
rect 48872 407124 48924 407176
rect 56968 407124 57020 407176
rect 357992 406376 358044 406428
rect 377220 406376 377272 406428
rect 48780 405696 48832 405748
rect 57060 405696 57112 405748
rect 377772 405628 377824 405680
rect 378140 405628 378192 405680
rect 51632 404948 51684 405000
rect 55864 404948 55916 405000
rect 204352 404948 204404 405000
rect 216864 404948 216916 405000
rect 359832 404948 359884 405000
rect 377312 404948 377364 405000
rect 51632 404336 51684 404388
rect 57060 404336 57112 404388
rect 359740 403588 359792 403640
rect 377772 403588 377824 403640
rect 52368 402976 52420 403028
rect 57060 402976 57112 403028
rect 199660 393320 199712 393372
rect 203248 393320 203300 393372
rect 199200 390872 199252 390924
rect 199844 390872 199896 390924
rect 198096 390532 198148 390584
rect 199108 390532 199160 390584
rect 198188 389172 198240 389224
rect 199476 389172 199528 389224
rect 520924 388424 520976 388476
rect 580356 388424 580408 388476
rect 44732 384956 44784 385008
rect 56600 384956 56652 385008
rect 206284 384956 206336 385008
rect 216956 384956 217008 385008
rect 359648 384956 359700 385008
rect 376944 384956 376996 385008
rect 208216 384276 208268 384328
rect 216680 384276 216732 384328
rect 57428 384208 57480 384260
rect 57428 384004 57480 384056
rect 46112 383596 46164 383648
rect 56600 383596 56652 383648
rect 57060 383596 57112 383648
rect 57980 383596 58032 383648
rect 207020 383596 207072 383648
rect 216680 383596 216732 383648
rect 359556 383596 359608 383648
rect 376944 383596 376996 383648
rect 51724 383528 51776 383580
rect 52920 383528 52972 383580
rect 202604 383528 202656 383580
rect 217048 383528 217100 383580
rect 206284 382236 206336 382288
rect 207020 382236 207072 382288
rect 41328 382168 41380 382220
rect 57244 382168 57296 382220
rect 367744 382168 367796 382220
rect 375380 382168 375432 382220
rect 376668 382168 376720 382220
rect 56048 380808 56100 380860
rect 57060 380808 57112 380860
rect 57336 378768 57388 378820
rect 57520 378768 57572 378820
rect 374000 378768 374052 378820
rect 374368 378768 374420 378820
rect 57152 378632 57204 378684
rect 57336 378632 57388 378684
rect 55772 375300 55824 375352
rect 59360 375300 59412 375352
rect 217232 375300 217284 375352
rect 217876 375300 217928 375352
rect 377864 375300 377916 375352
rect 379244 375300 379296 375352
rect 48872 375028 48924 375080
rect 217232 375028 217284 375080
rect 51632 374960 51684 375012
rect 216956 374960 217008 375012
rect 379428 374960 379480 375012
rect 380900 374960 380952 375012
rect 54392 374824 54444 374876
rect 56600 374824 56652 374876
rect 201500 374824 201552 374876
rect 275284 374824 275336 374876
rect 200212 374756 200264 374808
rect 295340 374756 295392 374808
rect 201040 374688 201092 374740
rect 305000 374688 305052 374740
rect 356888 374688 356940 374740
rect 452844 374688 452896 374740
rect 53656 374620 53708 374672
rect 59636 374620 59688 374672
rect 203064 374620 203116 374672
rect 312820 374620 312872 374672
rect 165988 374552 166040 374604
rect 199568 374552 199620 374604
rect 379244 374552 379296 374604
rect 425060 374552 425112 374604
rect 163412 374484 163464 374536
rect 197912 374484 197964 374536
rect 203156 374484 203208 374536
rect 213920 374484 213972 374536
rect 362868 374484 362920 374536
rect 410708 374484 410760 374536
rect 158536 374416 158588 374468
rect 201776 374416 201828 374468
rect 209504 374416 209556 374468
rect 320916 374416 320968 374468
rect 359464 374416 359516 374468
rect 407764 374416 407816 374468
rect 153476 374348 153528 374400
rect 200580 374348 200632 374400
rect 210240 374348 210292 374400
rect 210792 374348 210844 374400
rect 244280 374348 244332 374400
rect 372436 374348 372488 374400
rect 438492 374348 438544 374400
rect 160928 374280 160980 374332
rect 208492 374280 208544 374332
rect 369768 374280 369820 374332
rect 440332 374280 440384 374332
rect 156512 374212 156564 374264
rect 204536 374212 204588 374264
rect 217508 374212 217560 374264
rect 256056 374212 256108 374264
rect 360752 374212 360804 374264
rect 436008 374212 436060 374264
rect 58624 374144 58676 374196
rect 93584 374144 93636 374196
rect 148968 374144 149020 374196
rect 197084 374144 197136 374196
rect 199384 374144 199436 374196
rect 250720 374144 250772 374196
rect 358728 374144 358780 374196
rect 433616 374144 433668 374196
rect 56968 374076 57020 374128
rect 103520 374076 103572 374128
rect 146208 374076 146260 374128
rect 207480 374076 207532 374128
rect 241060 374076 241112 374128
rect 250076 374076 250128 374128
rect 366180 374076 366232 374128
rect 443092 374076 443144 374128
rect 54300 374008 54352 374060
rect 116032 374008 116084 374060
rect 143540 374008 143592 374060
rect 205916 374008 205968 374060
rect 213920 374008 213972 374060
rect 215116 374008 215168 374060
rect 236000 374008 236052 374060
rect 380900 374008 380952 374060
rect 405924 374008 405976 374060
rect 44640 373940 44692 373992
rect 217692 373940 217744 373992
rect 48780 373872 48832 373924
rect 217508 373872 217560 373924
rect 40776 373804 40828 373856
rect 199108 373804 199160 373856
rect 375288 373804 375340 373856
rect 416044 373804 416096 373856
rect 59728 373736 59780 373788
rect 107844 373736 107896 373788
rect 136456 373736 136508 373788
rect 200488 373736 200540 373788
rect 215300 373736 215352 373788
rect 217876 373736 217928 373788
rect 375932 373736 375984 373788
rect 418252 373736 418304 373788
rect 42340 373668 42392 373720
rect 100852 373668 100904 373720
rect 131028 373668 131080 373720
rect 199292 373668 199344 373720
rect 371792 373668 371844 373720
rect 423036 373668 423088 373720
rect 57060 373600 57112 373652
rect 118332 373600 118384 373652
rect 128912 373600 128964 373652
rect 198188 373600 198240 373652
rect 204260 373600 204312 373652
rect 215300 373600 215352 373652
rect 369768 373600 369820 373652
rect 375472 373600 375524 373652
rect 426900 373600 426952 373652
rect 52276 373532 52328 373584
rect 113548 373532 113600 373584
rect 133696 373532 133748 373584
rect 204444 373532 204496 373584
rect 368388 373532 368440 373584
rect 445852 373532 445904 373584
rect 48964 373464 49016 373516
rect 110420 373464 110472 373516
rect 125784 373464 125836 373516
rect 201684 373464 201736 373516
rect 214380 373464 214432 373516
rect 224224 373464 224276 373516
rect 370412 373464 370464 373516
rect 450268 373464 450320 373516
rect 43260 373396 43312 373448
rect 105452 373396 105504 373448
rect 121368 373396 121420 373448
rect 197820 373396 197872 373448
rect 210148 373396 210200 373448
rect 212540 373396 212592 373448
rect 256700 373396 256752 373448
rect 373724 373396 373776 373448
rect 455420 373396 455472 373448
rect 50160 373328 50212 373380
rect 98276 373328 98328 373380
rect 99380 373328 99432 373380
rect 204260 373328 204312 373380
rect 213092 373328 213144 373380
rect 214104 373328 214156 373380
rect 260012 373328 260064 373380
rect 363420 373328 363472 373380
rect 447692 373328 447744 373380
rect 57336 373260 57388 373312
rect 122932 373260 122984 373312
rect 191748 373260 191800 373312
rect 206284 373260 206336 373312
rect 262864 373260 262916 373312
rect 269212 373260 269264 373312
rect 358636 373260 358688 373312
rect 462780 373260 462832 373312
rect 49056 373192 49108 373244
rect 96068 373192 96120 373244
rect 139216 373192 139268 373244
rect 200672 373192 200724 373244
rect 215300 373192 215352 373244
rect 216496 373192 216548 373244
rect 236460 373192 236512 373244
rect 47584 373124 47636 373176
rect 88340 373124 88392 373176
rect 141608 373124 141660 373176
rect 203340 373124 203392 373176
rect 207204 373124 207256 373176
rect 213736 373124 213788 373176
rect 242900 373124 242952 373176
rect 55956 373056 56008 373108
rect 90180 373056 90232 373108
rect 151728 373056 151780 373108
rect 198096 373056 198148 373108
rect 220728 373056 220780 373108
rect 253940 373056 253992 373108
rect 42248 372988 42300 373040
rect 59728 372988 59780 373040
rect 212632 372988 212684 373040
rect 217968 372988 218020 373040
rect 255412 372988 255464 373040
rect 213920 372920 213972 372972
rect 219348 372920 219400 372972
rect 261300 372920 261352 372972
rect 212816 372852 212868 372904
rect 217140 372852 217192 372904
rect 258080 372852 258132 372904
rect 214012 372784 214064 372836
rect 259460 372784 259512 372836
rect 215392 372716 215444 372768
rect 262220 372716 262272 372768
rect 379152 372716 379204 372768
rect 379796 372716 379848 372768
rect 217876 372648 217928 372700
rect 264980 372648 265032 372700
rect 211160 372580 211212 372632
rect 217048 372580 217100 372632
rect 217692 372580 217744 372632
rect 219256 372580 219308 372632
rect 266360 372580 266412 372632
rect 362868 372580 362920 372632
rect 371240 372580 371292 372632
rect 379796 372580 379848 372632
rect 402888 372580 402940 372632
rect 84752 372512 84804 372564
rect 208400 372512 208452 372564
rect 210976 372512 211028 372564
rect 212356 372512 212408 372564
rect 218060 372512 218112 372564
rect 271880 372512 271932 372564
rect 275284 372512 275336 372564
rect 314660 372512 314712 372564
rect 373172 372512 373224 372564
rect 377404 372512 377456 372564
rect 86776 372444 86828 372496
rect 208216 372444 208268 372496
rect 215024 372444 215076 372496
rect 89352 372376 89404 372428
rect 209780 372376 209832 372428
rect 210056 372376 210108 372428
rect 295340 372444 295392 372496
rect 310520 372444 310572 372496
rect 312820 372444 312872 372496
rect 322940 372444 322992 372496
rect 244280 372376 244332 372428
rect 305000 372376 305052 372428
rect 313280 372376 313332 372428
rect 92388 372308 92440 372360
rect 211252 372308 211304 372360
rect 372896 372308 372948 372360
rect 400220 372308 400272 372360
rect 77208 372240 77260 372292
rect 99380 372240 99432 372292
rect 114468 372240 114520 372292
rect 219440 372240 219492 372292
rect 220728 372240 220780 372292
rect 93584 372172 93636 372224
rect 210976 372172 211028 372224
rect 214564 372172 214616 372224
rect 219716 372172 219768 372224
rect 220544 372172 220596 372224
rect 375196 372172 375248 372224
rect 379520 372172 379572 372224
rect 211252 372104 211304 372156
rect 221096 372104 221148 372156
rect 222108 372104 222160 372156
rect 371056 372104 371108 372156
rect 377956 372104 378008 372156
rect 379980 372104 380032 372156
rect 396080 372104 396132 372156
rect 47400 371968 47452 372020
rect 78496 371968 78548 372020
rect 92204 371968 92256 372020
rect 208216 371968 208268 372020
rect 213644 371968 213696 372020
rect 46204 371900 46256 371952
rect 79968 371900 80020 371952
rect 47492 371832 47544 371884
rect 80152 371832 80204 371884
rect 85488 371764 85540 371816
rect 105176 371764 105228 371816
rect 112904 371764 112956 371816
rect 212356 371900 212408 371952
rect 208768 371832 208820 371884
rect 209964 371832 210016 371884
rect 219624 372036 219676 372088
rect 241060 372036 241112 372088
rect 357164 372036 357216 372088
rect 380992 372036 381044 372088
rect 220544 371968 220596 372020
rect 251272 371968 251324 372020
rect 369860 371968 369912 372020
rect 370412 371968 370464 372020
rect 397460 371968 397512 372020
rect 220912 371900 220964 371952
rect 221832 371900 221884 371952
rect 252560 371900 252612 371952
rect 377864 371900 377916 371952
rect 404360 371900 404412 371952
rect 224224 371832 224276 371884
rect 247132 371832 247184 371884
rect 362776 371832 362828 371884
rect 210056 371764 210108 371816
rect 219532 371764 219584 371816
rect 248420 371764 248472 371816
rect 278688 371764 278740 371816
rect 356612 371764 356664 371816
rect 379336 371832 379388 371884
rect 422300 371832 422352 371884
rect 518440 371832 518492 371884
rect 580448 371832 580500 371884
rect 379152 371764 379204 371816
rect 407120 371764 407172 371816
rect 46296 371424 46348 371476
rect 49056 371424 49108 371476
rect 81992 371424 82044 371476
rect 208952 371696 209004 371748
rect 88064 371628 88116 371680
rect 209872 371628 209924 371680
rect 214380 371696 214432 371748
rect 241704 371696 241756 371748
rect 242808 371696 242860 371748
rect 276020 371696 276072 371748
rect 276940 371696 276992 371748
rect 356888 371696 356940 371748
rect 371240 371696 371292 371748
rect 371608 371696 371660 371748
rect 401600 371696 401652 371748
rect 90732 371424 90784 371476
rect 208768 371424 208820 371476
rect 208952 371424 209004 371476
rect 222108 371628 222160 371680
rect 251180 371628 251232 371680
rect 273352 371628 273404 371680
rect 305000 371628 305052 371680
rect 368388 371628 368440 371680
rect 378140 371628 378192 371680
rect 379520 371628 379572 371680
rect 379704 371628 379756 371680
rect 409880 371628 409932 371680
rect 210976 371560 211028 371612
rect 239312 371560 239364 371612
rect 367744 371560 367796 371612
rect 398840 371560 398892 371612
rect 79968 371356 80020 371408
rect 210056 371356 210108 371408
rect 80152 371288 80204 371340
rect 212448 371424 212500 371476
rect 240416 371492 240468 371544
rect 241428 371492 241480 371544
rect 242808 371492 242860 371544
rect 371240 371492 371292 371544
rect 377956 371492 378008 371544
rect 47400 371220 47452 371272
rect 47584 371220 47636 371272
rect 78496 371220 78548 371272
rect 216404 371356 216456 371408
rect 238116 371356 238168 371408
rect 369860 371424 369912 371476
rect 376576 371424 376628 371476
rect 380992 371492 381044 371544
rect 411260 371492 411312 371544
rect 241428 371356 241480 371408
rect 372896 371356 372948 371408
rect 373724 371356 373776 371408
rect 377036 371356 377088 371408
rect 377864 371356 377916 371408
rect 411352 371424 411404 371476
rect 380992 371356 381044 371408
rect 426440 371356 426492 371408
rect 213644 371288 213696 371340
rect 245660 371288 245712 371340
rect 342260 371288 342312 371340
rect 343364 371288 343416 371340
rect 360200 371288 360252 371340
rect 503536 371288 503588 371340
rect 517888 371288 517940 371340
rect 518440 371288 518492 371340
rect 220728 371220 220780 371272
rect 221004 371220 221056 371272
rect 273260 371220 273312 371272
rect 342904 371220 342956 371272
rect 357256 371220 357308 371272
rect 503168 371220 503220 371272
rect 517980 371220 518032 371272
rect 580264 371220 580316 371272
rect 40960 371152 41012 371204
rect 182824 371152 182876 371204
rect 198740 371152 198792 371204
rect 302240 371152 302292 371204
rect 356980 371152 357032 371204
rect 477500 371152 477552 371204
rect 54484 371084 54536 371136
rect 183468 371084 183520 371136
rect 198924 371084 198976 371136
rect 300860 371084 300912 371136
rect 362132 371084 362184 371136
rect 474740 371084 474792 371136
rect 102048 371016 102100 371068
rect 213920 371016 213972 371068
rect 217416 371016 217468 371068
rect 317420 371016 317472 371068
rect 364892 371016 364944 371068
rect 473360 371016 473412 371068
rect 197544 370948 197596 371000
rect 298100 370948 298152 371000
rect 360660 370948 360712 371000
rect 465080 370948 465132 371000
rect 197452 370880 197504 370932
rect 295340 370880 295392 370932
rect 367560 370880 367612 370932
rect 470600 370880 470652 370932
rect 210056 370812 210108 370864
rect 210976 370812 211028 370864
rect 212264 370812 212316 370864
rect 307760 370812 307812 370864
rect 364800 370812 364852 370864
rect 458180 370812 458232 370864
rect 198280 370744 198332 370796
rect 292580 370744 292632 370796
rect 365628 370744 365680 370796
rect 374552 370744 374604 370796
rect 375196 370744 375248 370796
rect 378140 370744 378192 370796
rect 427820 370744 427872 370796
rect 196808 370676 196860 370728
rect 289820 370676 289872 370728
rect 367008 370676 367060 370728
rect 413192 370676 413244 370728
rect 196716 370608 196768 370660
rect 287336 370608 287388 370660
rect 363512 370608 363564 370660
rect 374920 370608 374972 370660
rect 375288 370608 375340 370660
rect 378048 370608 378100 370660
rect 416780 370608 416832 370660
rect 196624 370540 196676 370592
rect 285680 370540 285732 370592
rect 362684 370540 362736 370592
rect 379888 370540 379940 370592
rect 414020 370540 414072 370592
rect 183468 370472 183520 370524
rect 195980 370472 196032 370524
rect 196900 370472 196952 370524
rect 282920 370472 282972 370524
rect 357072 370472 357124 370524
rect 373080 370472 373132 370524
rect 196992 370404 197044 370456
rect 277676 370404 277728 370456
rect 375196 370472 375248 370524
rect 415400 370472 415452 370524
rect 402980 370404 403032 370456
rect 198832 370336 198884 370388
rect 273352 370336 273404 370388
rect 375288 370336 375340 370388
rect 396080 370336 396132 370388
rect 202880 369792 202932 369844
rect 326160 369792 326212 369844
rect 363328 369792 363380 369844
rect 480260 369792 480312 369844
rect 202512 369724 202564 369776
rect 270500 369724 270552 369776
rect 369676 369724 369728 369776
rect 483020 369724 483072 369776
rect 77024 369656 77076 369708
rect 203156 369656 203208 369708
rect 206192 369656 206244 369708
rect 280160 369656 280212 369708
rect 361304 369656 361356 369708
rect 430580 369656 430632 369708
rect 211620 369588 211672 369640
rect 276020 369588 276072 369640
rect 358452 369588 358504 369640
rect 425060 369588 425112 369640
rect 208032 369520 208084 369572
rect 264980 369520 265032 369572
rect 372436 369520 372488 369572
rect 374368 369520 374420 369572
rect 378692 369520 378744 369572
rect 430672 369520 430724 369572
rect 208860 369452 208912 369504
rect 273444 369452 273496 369504
rect 373816 369452 373868 369504
rect 429200 369452 429252 369504
rect 205364 369384 205416 369436
rect 267740 369384 267792 369436
rect 370320 369384 370372 369436
rect 420920 369384 420972 369436
rect 203800 369316 203852 369368
rect 252560 369316 252612 369368
rect 358544 369316 358596 369368
rect 376944 369316 376996 369368
rect 423680 369316 423732 369368
rect 99288 369248 99340 369300
rect 212724 369248 212776 369300
rect 216312 369248 216364 369300
rect 260840 369248 260892 369300
rect 373908 369248 373960 369300
rect 375196 369248 375248 369300
rect 418160 369248 418212 369300
rect 106096 369180 106148 369232
rect 217876 369180 217928 369232
rect 219164 369180 219216 369232
rect 263600 369180 263652 369232
rect 366272 369180 366324 369232
rect 375840 369180 375892 369232
rect 419540 369180 419592 369232
rect 100484 369112 100536 369164
rect 212264 369112 212316 369164
rect 214012 369112 214064 369164
rect 214840 369112 214892 369164
rect 258172 369112 258224 369164
rect 210332 369044 210384 369096
rect 247040 369044 247092 369096
rect 367652 369044 367704 369096
rect 371792 369044 371844 369096
rect 421012 369112 421064 369164
rect 374460 369044 374512 369096
rect 375932 369044 375984 369096
rect 418252 369044 418304 369096
rect 97724 368976 97776 369028
rect 210148 368976 210200 369028
rect 210884 368976 210936 369028
rect 370228 368976 370280 369028
rect 371056 368976 371108 369028
rect 378692 368976 378744 369028
rect 105176 368908 105228 368960
rect 210240 368908 210292 368960
rect 210792 368908 210844 368960
rect 101128 368840 101180 368892
rect 213092 368840 213144 368892
rect 195980 368432 196032 368484
rect 196716 368432 196768 368484
rect 342260 368432 342312 368484
rect 372528 368432 372580 368484
rect 374460 368432 374512 368484
rect 375288 368432 375340 368484
rect 375748 368432 375800 368484
rect 376576 368432 376628 368484
rect 436100 368432 436152 368484
rect 374368 368364 374420 368416
rect 434720 368364 434772 368416
rect 361396 367888 361448 367940
rect 379336 367888 379388 367940
rect 412640 367888 412692 367940
rect 375288 367820 375340 367872
rect 431960 367820 432012 367872
rect 107568 367752 107620 367804
rect 214840 367752 214892 367804
rect 369032 367752 369084 367804
rect 373172 367752 373224 367804
rect 433340 367752 433392 367804
rect 374920 367548 374972 367600
rect 375196 367548 375248 367600
rect 199384 365644 199436 365696
rect 199568 365644 199620 365696
rect 199384 364964 199436 365016
rect 359188 364964 359240 365016
rect 359740 364964 359792 365016
rect 519176 364964 519228 365016
rect 519452 364964 519504 365016
rect 359832 363604 359884 363656
rect 519176 363604 519228 363656
rect 199660 362176 199712 362228
rect 200028 362176 200080 362228
rect 359004 362176 359056 362228
rect 359188 362176 359240 362228
rect 518992 362176 519044 362228
rect 519268 362176 519320 362228
rect 182824 360816 182876 360868
rect 197452 360816 197504 360868
rect 342904 360816 342956 360868
rect 359464 359524 359516 359576
rect 519084 359524 519136 359576
rect 199476 359456 199528 359508
rect 359004 359456 359056 359508
rect 359740 359456 359792 359508
rect 3332 358708 3384 358760
rect 18604 358708 18656 358760
rect 359096 357348 359148 357400
rect 359832 357348 359884 357400
rect 199568 356668 199620 356720
rect 199844 356668 199896 356720
rect 359096 356668 359148 356720
rect 179144 355988 179196 356040
rect 197268 355988 197320 356040
rect 357348 355988 357400 356040
rect 358820 355988 358872 356040
rect 500868 355444 500920 355496
rect 517612 355444 517664 355496
rect 338488 355376 338540 355428
rect 357440 355376 357492 355428
rect 498844 355376 498896 355428
rect 517704 355376 517756 355428
rect 191472 355308 191524 355360
rect 191748 355308 191800 355360
rect 214564 355308 214616 355360
rect 351736 355308 351788 355360
rect 375380 355308 375432 355360
rect 375380 355104 375432 355156
rect 376024 355104 376076 355156
rect 179696 354696 179748 354748
rect 197544 354696 197596 354748
rect 201592 354696 201644 354748
rect 339776 354696 339828 354748
rect 357348 354696 357400 354748
rect 510896 354696 510948 354748
rect 517520 354696 517572 354748
rect 371700 353948 371752 354000
rect 380900 353948 380952 354000
rect 218428 353404 218480 353456
rect 221096 353404 221148 353456
rect 56048 353336 56100 353388
rect 59820 353336 59872 353388
rect 218612 353336 218664 353388
rect 220912 353336 220964 353388
rect 378692 353336 378744 353388
rect 381084 353336 381136 353388
rect 58532 353268 58584 353320
rect 60740 353268 60792 353320
rect 218520 353268 218572 353320
rect 220820 353268 220872 353320
rect 378600 353268 378652 353320
rect 380992 353268 381044 353320
rect 57060 351976 57112 352028
rect 59360 351976 59412 352028
rect 55956 351908 56008 351960
rect 57980 351908 58032 351960
rect 54484 303764 54536 303816
rect 56600 303764 56652 303816
rect 46388 299412 46440 299464
rect 56968 299412 57020 299464
rect 57428 299412 57480 299464
rect 46480 298052 46532 298104
rect 57428 298052 57480 298104
rect 519912 284316 519964 284368
rect 580264 284316 580316 284368
rect 519176 282888 519228 282940
rect 580356 282888 580408 282940
rect 377772 282208 377824 282260
rect 377956 282208 378008 282260
rect 200948 280100 201000 280152
rect 216680 280100 216732 280152
rect 368296 280100 368348 280152
rect 377036 280100 377088 280152
rect 205272 278672 205324 278724
rect 216864 278672 216916 278724
rect 366916 278672 366968 278724
rect 377036 278672 377088 278724
rect 214564 278264 214616 278316
rect 216680 278264 216732 278316
rect 376024 278264 376076 278316
rect 377404 278264 377456 278316
rect 214564 276564 214616 276616
rect 215300 276564 215352 276616
rect 377772 274116 377824 274168
rect 377956 274116 378008 274168
rect 213092 272552 213144 272604
rect 213644 272552 213696 272604
rect 211712 270444 211764 270496
rect 212908 270444 212960 270496
rect 378600 270444 378652 270496
rect 379520 270444 379572 270496
rect 219256 270036 219308 270088
rect 219808 270036 219860 270088
rect 60832 269628 60884 269680
rect 107568 269628 107620 269680
rect 55864 269560 55916 269612
rect 110972 269560 111024 269612
rect 219808 269560 219860 269612
rect 263508 269560 263560 269612
rect 52920 269492 52972 269544
rect 108304 269492 108356 269544
rect 200856 269492 200908 269544
rect 250720 269492 250772 269544
rect 43352 269424 43404 269476
rect 133420 269424 133472 269476
rect 218520 269424 218572 269476
rect 279148 269424 279200 269476
rect 379244 269424 379296 269476
rect 425244 269424 425296 269476
rect 45376 269356 45428 269408
rect 135904 269356 135956 269408
rect 212908 269356 212960 269408
rect 275744 269356 275796 269408
rect 379520 269356 379572 269408
rect 426440 269356 426492 269408
rect 44824 269288 44876 269340
rect 138480 269288 138532 269340
rect 214748 269288 214800 269340
rect 280896 269288 280948 269340
rect 364156 269288 364208 269340
rect 418436 269288 418488 269340
rect 45008 269220 45060 269272
rect 140872 269220 140924 269272
rect 210700 269220 210752 269272
rect 283472 269220 283524 269272
rect 373632 269220 373684 269272
rect 433616 269220 433668 269272
rect 45100 269152 45152 269204
rect 143540 269152 143592 269204
rect 212172 269152 212224 269204
rect 288256 269152 288308 269204
rect 370964 269152 371016 269204
rect 453396 269152 453448 269204
rect 44916 269084 44968 269136
rect 145932 269084 145984 269136
rect 209320 269084 209372 269136
rect 285956 269084 286008 269136
rect 368204 269084 368256 269136
rect 468484 269084 468536 269136
rect 42524 269016 42576 269068
rect 59636 269016 59688 269068
rect 60740 269016 60792 269068
rect 196624 269016 196676 269068
rect 197636 269016 197688 269068
rect 213644 269016 213696 269068
rect 214288 269016 214340 269068
rect 217140 269016 217192 269068
rect 217784 269016 217836 269068
rect 374460 269016 374512 269068
rect 374920 269016 374972 269068
rect 60832 268948 60884 269000
rect 374552 268880 374604 268932
rect 396080 268880 396132 268932
rect 206560 268812 206612 268864
rect 290924 268812 290976 268864
rect 369124 268812 369176 268864
rect 423496 268812 423548 268864
rect 49240 268744 49292 268796
rect 83096 268744 83148 268796
rect 207940 268744 207992 268796
rect 295892 268744 295944 268796
rect 366824 268744 366876 268796
rect 421012 268744 421064 268796
rect 42616 268676 42668 268728
rect 57796 268676 57848 268728
rect 203616 268676 203668 268728
rect 293408 268676 293460 268728
rect 376392 268676 376444 268728
rect 430948 268676 431000 268728
rect 47768 268608 47820 268660
rect 77116 268608 77168 268660
rect 216220 268608 216272 268660
rect 308496 268608 308548 268660
rect 375104 268608 375156 268660
rect 478420 268608 478472 268660
rect 45192 268540 45244 268592
rect 47400 268540 47452 268592
rect 47952 268540 48004 268592
rect 90732 268540 90784 268592
rect 202420 268540 202472 268592
rect 298468 268540 298520 268592
rect 372344 268540 372396 268592
rect 475844 268540 475896 268592
rect 48044 268472 48096 268524
rect 93584 268472 93636 268524
rect 205180 268472 205232 268524
rect 300860 268472 300912 268524
rect 362592 268472 362644 268524
rect 473360 268472 473412 268524
rect 43444 268404 43496 268456
rect 47308 268404 47360 268456
rect 49148 268404 49200 268456
rect 96068 268404 96120 268456
rect 213460 268404 213512 268456
rect 318432 268404 318484 268456
rect 365536 268404 365588 268456
rect 480904 268404 480956 268456
rect 51816 268336 51868 268388
rect 98460 268336 98512 268388
rect 198004 268336 198056 268388
rect 315856 268336 315908 268388
rect 361028 268336 361080 268388
rect 483388 268336 483440 268388
rect 46664 268268 46716 268320
rect 76012 268268 76064 268320
rect 47216 268200 47268 268252
rect 47768 268200 47820 268252
rect 64880 268200 64932 268252
rect 95884 268200 95936 268252
rect 62120 268132 62172 268184
rect 94504 268132 94556 268184
rect 53840 268064 53892 268116
rect 86960 268064 87012 268116
rect 373172 268064 373224 268116
rect 374276 268064 374328 268116
rect 433340 268064 433392 268116
rect 58624 267996 58676 268048
rect 82084 267996 82136 268048
rect 108672 267996 108724 268048
rect 396080 267996 396132 268048
rect 415860 267996 415912 268048
rect 99380 267928 99432 267980
rect 236644 267928 236696 267980
rect 255780 267928 255832 267980
rect 356520 267928 356572 267980
rect 360200 267928 360252 267980
rect 373080 267928 373132 267980
rect 375656 267928 375708 267980
rect 402980 267928 403032 267980
rect 57796 267860 57848 267912
rect 105268 267860 105320 267912
rect 214288 267860 214340 267912
rect 243084 267860 243136 267912
rect 379888 267860 379940 267912
rect 414388 267860 414440 267912
rect 421564 267860 421616 267912
rect 435732 267860 435784 267912
rect 59728 267792 59780 267844
rect 106372 267792 106424 267844
rect 217784 267792 217836 267844
rect 258080 267792 258132 267844
rect 374920 267792 374972 267844
rect 432144 267792 432196 267844
rect 54484 267724 54536 267776
rect 102692 267724 102744 267776
rect 117136 267724 117188 267776
rect 196624 267724 196676 267776
rect 219348 267724 219400 267776
rect 261668 267724 261720 267776
rect 42432 267656 42484 267708
rect 122840 267656 122892 267708
rect 158536 267656 158588 267708
rect 206008 267656 206060 267708
rect 357256 267656 357308 267708
rect 357532 267656 357584 267708
rect 361120 267656 361172 267708
rect 458180 267656 458232 267708
rect 47676 267588 47728 267640
rect 53840 267588 53892 267640
rect 55956 267588 56008 267640
rect 129740 267588 129792 267640
rect 153568 267588 153620 267640
rect 200304 267588 200356 267640
rect 216128 267588 216180 267640
rect 302240 267588 302292 267640
rect 362500 267588 362552 267640
rect 455788 267588 455840 267640
rect 57060 267520 57112 267572
rect 128360 267520 128412 267572
rect 155960 267520 156012 267572
rect 202972 267520 203024 267572
rect 206744 267520 206796 267572
rect 276020 267520 276072 267572
rect 364064 267520 364116 267572
rect 445760 267520 445812 267572
rect 56048 267452 56100 267504
rect 125600 267452 125652 267504
rect 163504 267452 163556 267504
rect 197728 267452 197780 267504
rect 202328 267452 202380 267504
rect 270868 267452 270920 267504
rect 370872 267452 370924 267504
rect 449900 267452 449952 267504
rect 54760 267384 54812 267436
rect 120080 267384 120132 267436
rect 166172 267384 166224 267436
rect 200396 267384 200448 267436
rect 203708 267384 203760 267436
rect 268200 267384 268252 267436
rect 369492 267384 369544 267436
rect 447140 267384 447192 267436
rect 46756 267316 46808 267368
rect 51356 267316 51408 267368
rect 53012 267316 53064 267368
rect 117320 267316 117372 267368
rect 160928 267316 160980 267368
rect 207112 267316 207164 267368
rect 213552 267316 213604 267368
rect 273260 267316 273312 267368
rect 53196 267248 53248 267300
rect 115940 267248 115992 267300
rect 204996 267248 205048 267300
rect 263600 267248 263652 267300
rect 53104 267180 53156 267232
rect 113180 267180 113232 267232
rect 207848 267180 207900 267232
rect 260840 267180 260892 267232
rect 343456 267180 343508 267232
rect 356520 267316 356572 267368
rect 356980 267316 357032 267368
rect 358360 267316 358412 267368
rect 435916 267316 435968 267368
rect 361212 267248 361264 267300
rect 437480 267248 437532 267300
rect 356520 267180 356572 267232
rect 356888 267180 356940 267232
rect 372252 267180 372304 267232
rect 443000 267180 443052 267232
rect 51908 267112 51960 267164
rect 104900 267112 104952 267164
rect 183468 267112 183520 267164
rect 196716 267112 196768 267164
rect 211988 267112 212040 267164
rect 265808 267112 265860 267164
rect 278136 267112 278188 267164
rect 356612 267112 356664 267164
rect 373448 267112 373500 267164
rect 440240 267112 440292 267164
rect 503536 267112 503588 267164
rect 517888 267112 517940 267164
rect 47492 267044 47544 267096
rect 47768 267044 47820 267096
rect 52000 267044 52052 267096
rect 103520 267044 103572 267096
rect 206652 267044 206704 267096
rect 258264 267044 258316 267096
rect 343548 267044 343600 267096
rect 357532 267044 357584 267096
rect 369584 267044 369636 267096
rect 416044 267044 416096 267096
rect 50344 266976 50396 267028
rect 100760 266976 100812 267028
rect 183284 266976 183336 267028
rect 197452 266976 197504 267028
rect 214932 266976 214984 267028
rect 273260 266976 273312 267028
rect 277124 266976 277176 267028
rect 356520 266976 356572 267028
rect 365444 266976 365496 267028
rect 409880 266976 409932 267028
rect 503444 266976 503496 267028
rect 517980 266976 518032 267028
rect 54668 266908 54720 266960
rect 88340 266908 88392 266960
rect 210608 266908 210660 266960
rect 255320 266908 255372 266960
rect 379428 266908 379480 266960
rect 422576 266908 422628 266960
rect 47768 266840 47820 266892
rect 80060 266840 80112 266892
rect 213184 266840 213236 266892
rect 252560 266840 252612 266892
rect 375012 266840 375064 266892
rect 412916 266840 412968 266892
rect 47584 266772 47636 266824
rect 77300 266772 77352 266824
rect 219072 266772 219124 266824
rect 247040 266772 247092 266824
rect 376484 266772 376536 266824
rect 407120 266772 407172 266824
rect 214656 266704 214708 266756
rect 310520 266704 310572 266756
rect 214564 266432 214616 266484
rect 214932 266432 214984 266484
rect 214656 266364 214708 266416
rect 215392 266364 215444 266416
rect 356612 266364 356664 266416
rect 356796 266364 356848 266416
rect 425704 266364 425756 266416
rect 434260 266364 434312 266416
rect 517704 266364 517756 266416
rect 517888 266364 517940 266416
rect 50344 266296 50396 266348
rect 57704 266296 57756 266348
rect 92388 266296 92440 266348
rect 262220 266296 262272 266348
rect 379796 266296 379848 266348
rect 403164 266296 403216 266348
rect 63500 266228 63552 266280
rect 92480 266228 92532 266280
rect 218612 266228 218664 266280
rect 219164 266228 219216 266280
rect 252560 266228 252612 266280
rect 378692 266228 378744 266280
rect 411260 266228 411312 266280
rect 54116 266160 54168 266212
rect 84200 266160 84252 266212
rect 216772 266160 216824 266212
rect 218428 266160 218480 266212
rect 251272 266160 251324 266212
rect 379704 266160 379756 266212
rect 409880 266160 409932 266212
rect 58716 266092 58768 266144
rect 89720 266092 89772 266144
rect 213644 266092 213696 266144
rect 245660 266092 245712 266144
rect 371608 266092 371660 266144
rect 372344 266092 372396 266144
rect 401692 266092 401744 266144
rect 53932 266024 53984 266076
rect 85580 266024 85632 266076
rect 219072 266024 219124 266076
rect 219716 266024 219768 266076
rect 251180 266024 251232 266076
rect 379152 266024 379204 266076
rect 407120 266024 407172 266076
rect 85396 265956 85448 266008
rect 220728 265956 220780 266008
rect 249800 265956 249852 266008
rect 373632 265956 373684 266008
rect 400220 265956 400272 266008
rect 54576 265888 54628 265940
rect 56048 265888 56100 265940
rect 88340 265888 88392 265940
rect 213092 265888 213144 265940
rect 213644 265888 213696 265940
rect 219256 265888 219308 265940
rect 219532 265888 219584 265940
rect 248512 265888 248564 265940
rect 376576 265888 376628 265940
rect 377864 265888 377916 265940
rect 404360 265888 404412 265940
rect 50252 265820 50304 265872
rect 52000 265820 52052 265872
rect 78588 265820 78640 265872
rect 111800 265820 111852 265872
rect 57704 265752 57756 265804
rect 91100 265752 91152 265804
rect 244280 265820 244332 265872
rect 370412 265820 370464 265872
rect 372528 265820 372580 265872
rect 398196 265820 398248 265872
rect 52552 265684 52604 265736
rect 100760 265684 100812 265736
rect 215024 265684 215076 265736
rect 216312 265684 216364 265736
rect 52736 265616 52788 265668
rect 113272 265616 113324 265668
rect 214380 265616 214432 265668
rect 216220 265616 216272 265668
rect 247040 265752 247092 265804
rect 367744 265752 367796 265804
rect 370964 265752 371016 265804
rect 398840 265752 398892 265804
rect 217876 265684 217928 265736
rect 219716 265684 219768 265736
rect 265164 265684 265216 265736
rect 373724 265684 373776 265736
rect 376576 265684 376628 265736
rect 376668 265684 376720 265736
rect 378600 265684 378652 265736
rect 408500 265684 408552 265736
rect 214840 265548 214892 265600
rect 218520 265548 218572 265600
rect 267096 265616 267148 265668
rect 371700 265616 371752 265668
rect 373172 265616 373224 265668
rect 405740 265616 405792 265668
rect 377956 265480 378008 265532
rect 411352 265480 411404 265532
rect 375288 265344 375340 265396
rect 375104 265276 375156 265328
rect 379796 265276 379848 265328
rect 375196 265208 375248 265260
rect 379980 265208 380032 265260
rect 377036 265140 377088 265192
rect 377956 265140 378008 265192
rect 213000 265072 213052 265124
rect 215760 265072 215812 265124
rect 230388 265072 230440 265124
rect 375748 265072 375800 265124
rect 379152 265072 379204 265124
rect 212264 265004 212316 265056
rect 215668 265004 215720 265056
rect 233148 265004 233200 265056
rect 377956 265004 378008 265056
rect 379704 265004 379756 265056
rect 210884 264936 210936 264988
rect 214748 264936 214800 264988
rect 231768 264936 231820 264988
rect 374552 264936 374604 264988
rect 375288 264936 375340 264988
rect 378692 264936 378744 264988
rect 379244 264936 379296 264988
rect 391940 264936 391992 264988
rect 48136 264868 48188 264920
rect 54116 264868 54168 264920
rect 54484 264868 54536 264920
rect 212356 264868 212408 264920
rect 272156 264868 272208 264920
rect 378048 264868 378100 264920
rect 416780 264868 416832 264920
rect 45468 264800 45520 264852
rect 58716 264800 58768 264852
rect 219900 264800 219952 264852
rect 253940 264800 253992 264852
rect 379336 264800 379388 264852
rect 412916 264800 412968 264852
rect 43996 264732 44048 264784
rect 57244 264732 57296 264784
rect 57704 264732 57756 264784
rect 230388 264732 230440 264784
rect 259552 264732 259604 264784
rect 369768 264732 369820 264784
rect 378968 264732 379020 264784
rect 388168 264732 388220 264784
rect 420920 264732 420972 264784
rect 43812 264664 43864 264716
rect 52552 264664 52604 264716
rect 53104 264664 53156 264716
rect 233148 264664 233200 264716
rect 259460 264664 259512 264716
rect 389180 264664 389232 264716
rect 419540 264664 419592 264716
rect 46848 264596 46900 264648
rect 53932 264596 53984 264648
rect 54576 264596 54628 264648
rect 231768 264596 231820 264648
rect 256700 264596 256752 264648
rect 390560 264596 390612 264648
rect 418252 264596 418304 264648
rect 46572 264528 46624 264580
rect 147680 264528 147732 264580
rect 391940 264528 391992 264580
rect 418160 264528 418212 264580
rect 43904 264392 43956 264444
rect 47952 264392 48004 264444
rect 63500 264392 63552 264444
rect 45284 264324 45336 264376
rect 47492 264324 47544 264376
rect 78588 264324 78640 264376
rect 210792 264324 210844 264376
rect 215024 264324 215076 264376
rect 244372 264324 244424 264376
rect 43720 264256 43772 264308
rect 49148 264256 49200 264308
rect 82084 264256 82136 264308
rect 208124 264256 208176 264308
rect 214932 264256 214984 264308
rect 269764 264256 269816 264308
rect 43628 264188 43680 264240
rect 47860 264188 47912 264240
rect 96620 264188 96672 264240
rect 209504 264188 209556 264240
rect 213460 264188 213512 264240
rect 271236 264188 271288 264240
rect 377128 263576 377180 263628
rect 378048 263576 378100 263628
rect 378692 263576 378744 263628
rect 379336 263576 379388 263628
rect 376392 263508 376444 263560
rect 436100 263508 436152 263560
rect 378048 263440 378100 263492
rect 437480 263440 437532 263492
rect 375840 263100 375892 263152
rect 376392 263100 376444 263152
rect 357440 252560 357492 252612
rect 356888 252492 356940 252544
rect 213184 251132 213236 251184
rect 215300 251132 215352 251184
rect 215852 251132 215904 251184
rect 263600 251132 263652 251184
rect 340236 251132 340288 251184
rect 357440 251200 357492 251252
rect 368388 251132 368440 251184
rect 371792 251132 371844 251184
rect 373448 251132 373500 251184
rect 373816 251132 373868 251184
rect 430580 251132 430632 251184
rect 217140 251064 217192 251116
rect 217968 251064 218020 251116
rect 236644 251064 236696 251116
rect 372252 251064 372304 251116
rect 372436 251064 372488 251116
rect 421564 251064 421616 251116
rect 517612 251064 517664 251116
rect 517888 251064 517940 251116
rect 197360 250928 197412 250980
rect 197544 250928 197596 250980
rect 371148 250724 371200 250776
rect 374460 250724 374512 250776
rect 425704 250724 425756 250776
rect 371056 250656 371108 250708
rect 373540 250656 373592 250708
rect 430672 250656 430724 250708
rect 180248 250588 180300 250640
rect 197636 250588 197688 250640
rect 371792 250588 371844 250640
rect 429200 250588 429252 250640
rect 500408 250588 500460 250640
rect 517888 250588 517940 250640
rect 82820 250520 82872 250572
rect 100852 250520 100904 250572
rect 209596 250520 209648 250572
rect 67548 250452 67600 250504
rect 98000 250452 98052 250504
rect 179328 250452 179380 250504
rect 197544 250452 197596 250504
rect 338488 250520 338540 250572
rect 356888 250520 356940 250572
rect 362868 250520 362920 250572
rect 372436 250520 372488 250572
rect 438860 250520 438912 250572
rect 499028 250520 499080 250572
rect 517796 250520 517848 250572
rect 219624 250452 219676 250504
rect 267740 250452 267792 250504
rect 279976 250452 280028 250504
rect 357624 250452 357676 250504
rect 379704 250452 379756 250504
rect 396080 250452 396132 250504
rect 510896 249840 510948 249892
rect 517520 249840 517572 249892
rect 190920 249772 190972 249824
rect 213184 249772 213236 249824
rect 351000 249772 351052 249824
rect 369124 249772 369176 249824
rect 376024 249772 376076 249824
rect 50436 249704 50488 249756
rect 52736 249704 52788 249756
rect 58440 249704 58492 249756
rect 60924 249704 60976 249756
rect 58532 249636 58584 249688
rect 60832 249636 60884 249688
rect 55956 249364 56008 249416
rect 61016 249364 61068 249416
rect 54668 249160 54720 249212
rect 60740 249160 60792 249212
rect 52736 249092 52788 249144
rect 67548 249092 67600 249144
rect 53012 249024 53064 249076
rect 82820 249024 82872 249076
rect 42708 248344 42760 248396
rect 52920 248344 52972 248396
rect 52736 243652 52788 243704
rect 53012 243652 53064 243704
rect 52828 243584 52880 243636
rect 52828 243380 52880 243432
rect 3056 202784 3108 202836
rect 40684 202784 40736 202836
rect 520188 182180 520240 182232
rect 580264 182180 580316 182232
rect 519268 182112 519320 182164
rect 519452 182112 519504 182164
rect 580356 182112 580408 182164
rect 207756 175176 207808 175228
rect 216680 175176 216732 175228
rect 363972 175176 364024 175228
rect 376852 175176 376904 175228
rect 369124 173816 369176 173868
rect 376852 173816 376904 173868
rect 203524 173748 203576 173800
rect 217048 173748 217100 173800
rect 372160 173748 372212 173800
rect 376760 173748 376812 173800
rect 198004 173136 198056 173188
rect 213184 173136 213236 173188
rect 216680 173136 216732 173188
rect 358728 173136 358780 173188
rect 369124 173136 369176 173188
rect 374460 165520 374512 165572
rect 375564 165520 375616 165572
rect 375564 164432 375616 164484
rect 434352 164432 434404 164484
rect 50528 164364 50580 164416
rect 96068 164364 96120 164416
rect 363788 164364 363840 164416
rect 425980 164364 426032 164416
rect 59084 164296 59136 164348
rect 140872 164296 140924 164348
rect 205088 164296 205140 164348
rect 258448 164296 258500 164348
rect 366732 164296 366784 164348
rect 451004 164296 451056 164348
rect 41052 164228 41104 164280
rect 163320 164228 163372 164280
rect 202236 164228 202288 164280
rect 318432 164228 318484 164280
rect 362408 164228 362460 164280
rect 480904 164228 480956 164280
rect 375840 164160 375892 164212
rect 376392 164160 376444 164212
rect 374552 164092 374604 164144
rect 393320 164092 393372 164144
rect 394516 164092 394568 164144
rect 49424 164024 49476 164076
rect 98460 164024 98512 164076
rect 365168 164024 365220 164076
rect 423496 164024 423548 164076
rect 52092 163956 52144 164008
rect 101036 163956 101088 164008
rect 362316 163956 362368 164008
rect 421012 163956 421064 164008
rect 50804 163888 50856 163940
rect 103520 163888 103572 163940
rect 356704 163888 356756 163940
rect 416044 163888 416096 163940
rect 52184 163820 52236 163872
rect 105912 163820 105964 163872
rect 366640 163820 366692 163872
rect 428188 163820 428240 163872
rect 50712 163752 50764 163804
rect 108212 163752 108264 163804
rect 116216 163752 116268 163804
rect 117044 163752 117096 163804
rect 196624 163752 196676 163804
rect 369308 163752 369360 163804
rect 430948 163752 431000 163804
rect 60004 163684 60056 163736
rect 145932 163684 145984 163736
rect 213368 163684 213420 163736
rect 261024 163684 261076 163736
rect 369400 163684 369452 163736
rect 470600 163684 470652 163736
rect 59176 163616 59228 163668
rect 148508 163616 148560 163668
rect 209136 163616 209188 163668
rect 298468 163616 298520 163668
rect 372068 163616 372120 163668
rect 473452 163616 473504 163668
rect 510528 163616 510580 163668
rect 517520 163616 517572 163668
rect 59912 163548 59964 163600
rect 150900 163548 150952 163600
rect 211896 163548 211948 163600
rect 305920 163548 305972 163600
rect 373356 163548 373408 163600
rect 475844 163548 475896 163600
rect 58900 163480 58952 163532
rect 153384 163480 153436 163532
rect 206376 163480 206428 163532
rect 300860 163480 300912 163532
rect 368112 163480 368164 163532
rect 478420 163480 478472 163532
rect 196716 163412 196768 163464
rect 197360 163412 197412 163464
rect 377128 163140 377180 163192
rect 396724 163140 396776 163192
rect 394516 163072 394568 163124
rect 415308 163072 415360 163124
rect 374920 163004 374972 163056
rect 431960 163004 432012 163056
rect 378416 162936 378468 162988
rect 438032 162936 438084 162988
rect 52920 162868 52972 162920
rect 54392 162868 54444 162920
rect 73804 162868 73856 162920
rect 218244 162868 218296 162920
rect 218520 162868 218572 162920
rect 267556 162868 267608 162920
rect 376392 162868 376444 162920
rect 436928 162868 436980 162920
rect 55128 162800 55180 162852
rect 133420 162800 133472 162852
rect 209044 162800 209096 162852
rect 320916 162800 320968 162852
rect 356704 162800 356756 162852
rect 356980 162800 357032 162852
rect 415308 162800 415360 162852
rect 418160 162800 418212 162852
rect 517612 162800 517664 162852
rect 517980 162800 518032 162852
rect 56232 162732 56284 162784
rect 130844 162732 130896 162784
rect 204904 162732 204956 162784
rect 308588 162732 308640 162784
rect 365260 162732 365312 162784
rect 455788 162732 455840 162784
rect 54852 162664 54904 162716
rect 128360 162664 128412 162716
rect 207664 162664 207716 162716
rect 303436 162664 303488 162716
rect 370688 162664 370740 162716
rect 458364 162664 458416 162716
rect 56140 162596 56192 162648
rect 125876 162596 125928 162648
rect 218888 162596 218940 162648
rect 293316 162596 293368 162648
rect 363880 162596 363932 162648
rect 448244 162596 448296 162648
rect 55036 162528 55088 162580
rect 122840 162528 122892 162580
rect 211804 162528 211856 162580
rect 283748 162528 283800 162580
rect 371976 162528 372028 162580
rect 445852 162528 445904 162580
rect 53380 162460 53432 162512
rect 120724 162460 120776 162512
rect 215944 162460 215996 162512
rect 285956 162460 286008 162512
rect 369216 162460 369268 162512
rect 440884 162460 440936 162512
rect 53288 162392 53340 162444
rect 115940 162392 115992 162444
rect 210516 162392 210568 162444
rect 278412 162392 278464 162444
rect 368020 162392 368072 162444
rect 438492 162392 438544 162444
rect 56416 162324 56468 162376
rect 118332 162324 118384 162376
rect 206468 162324 206520 162376
rect 268292 162324 268344 162376
rect 374828 162324 374880 162376
rect 443460 162324 443512 162376
rect 54944 162256 54996 162308
rect 113548 162256 113600 162308
rect 183468 162256 183520 162308
rect 197360 162256 197412 162308
rect 218980 162256 219032 162308
rect 280804 162256 280856 162308
rect 343456 162256 343508 162308
rect 356704 162256 356756 162308
rect 366548 162256 366600 162308
rect 433524 162256 433576 162308
rect 503260 162256 503312 162308
rect 517612 162256 517664 162308
rect 53564 162188 53616 162240
rect 110972 162188 111024 162240
rect 216036 162188 216088 162240
rect 273444 162188 273496 162240
rect 370596 162188 370648 162240
rect 435916 162188 435968 162240
rect 48228 162120 48280 162172
rect 93676 162120 93728 162172
rect 183192 162120 183244 162172
rect 197452 162120 197504 162172
rect 210424 162120 210476 162172
rect 265440 162120 265492 162172
rect 343364 162120 343416 162172
rect 357532 162120 357584 162172
rect 358084 162120 358136 162172
rect 413652 162120 413704 162172
rect 503628 162120 503680 162172
rect 517520 162120 517572 162172
rect 49332 162052 49384 162104
rect 90732 162052 90784 162104
rect 202144 162052 202196 162104
rect 255964 162052 256016 162104
rect 358268 162052 358320 162104
rect 408316 162052 408368 162104
rect 56508 161984 56560 162036
rect 88340 161984 88392 162036
rect 213276 161984 213328 162036
rect 263692 161984 263744 162036
rect 378784 161984 378836 162036
rect 418436 161984 418488 162036
rect 218796 161916 218848 161968
rect 247868 161916 247920 161968
rect 376300 161916 376352 161968
rect 410616 161916 410668 161968
rect 360936 161848 360988 161900
rect 453212 161848 453264 161900
rect 421564 161576 421616 161628
rect 439044 161576 439096 161628
rect 87604 161440 87656 161492
rect 96896 161440 96948 161492
rect 55956 161372 56008 161424
rect 117320 161372 117372 161424
rect 219532 161372 219584 161424
rect 267740 161372 267792 161424
rect 372252 161372 372304 161424
rect 435364 161508 435416 161560
rect 434720 161440 434772 161492
rect 434628 161372 434680 161424
rect 54668 161304 54720 161356
rect 114744 161304 114796 161356
rect 216036 161304 216088 161356
rect 263600 161304 263652 161356
rect 379520 161304 379572 161356
rect 426440 161304 426492 161356
rect 59176 161236 59228 161288
rect 106372 161236 106424 161288
rect 219808 161236 219860 161288
rect 266360 161236 266412 161288
rect 379336 161236 379388 161288
rect 422300 161236 422352 161288
rect 59728 161168 59780 161220
rect 106280 161168 106332 161220
rect 219624 161168 219676 161220
rect 264980 161168 265032 161220
rect 59084 161100 59136 161152
rect 53012 161032 53064 161084
rect 56508 161032 56560 161084
rect 219348 161100 219400 161152
rect 260840 161100 260892 161152
rect 58532 160964 58584 161016
rect 59176 160964 59228 161016
rect 95240 161032 95292 161084
rect 217784 161032 217836 161084
rect 258080 161032 258132 161084
rect 98000 160964 98052 161016
rect 47400 160896 47452 160948
rect 53472 160896 53524 160948
rect 109040 160896 109092 160948
rect 47308 160828 47360 160880
rect 52092 160828 52144 160880
rect 110420 160828 110472 160880
rect 211528 160828 211580 160880
rect 213368 160828 213420 160880
rect 52368 160760 52420 160812
rect 59084 160760 59136 160812
rect 59360 160760 59412 160812
rect 118700 160760 118752 160812
rect 262220 160760 262272 160812
rect 373448 160760 373500 160812
rect 376300 160760 376352 160812
rect 429292 160760 429344 160812
rect 47492 160692 47544 160744
rect 52184 160692 52236 160744
rect 111800 160692 111852 160744
rect 214656 160692 214708 160744
rect 216128 160692 216180 160744
rect 213368 160624 213420 160676
rect 273260 160692 273312 160744
rect 373540 160692 373592 160744
rect 374828 160692 374880 160744
rect 430580 160692 430632 160744
rect 59728 160284 59780 160336
rect 60004 160284 60056 160336
rect 53564 160080 53616 160132
rect 54668 160080 54720 160132
rect 58440 160080 58492 160132
rect 59360 160080 59412 160132
rect 218428 160080 218480 160132
rect 219348 160080 219400 160132
rect 379520 160080 379572 160132
rect 379888 160080 379940 160132
rect 215760 160012 215812 160064
rect 259460 160012 259512 160064
rect 376668 160012 376720 160064
rect 420920 160012 420972 160064
rect 215668 159944 215720 159996
rect 259552 159944 259604 159996
rect 375380 159944 375432 159996
rect 419540 159944 419592 159996
rect 378048 159876 378100 159928
rect 418160 159876 418212 159928
rect 214748 159332 214800 159384
rect 218888 159332 218940 159384
rect 256700 159332 256752 159384
rect 215760 159196 215812 159248
rect 216404 159196 216456 159248
rect 215208 158720 215260 158772
rect 215668 158720 215720 158772
rect 377128 156612 377180 156664
rect 378048 156612 378100 156664
rect 53012 148996 53064 149048
rect 53196 148996 53248 149048
rect 114560 148996 114612 149048
rect 213552 148996 213604 149048
rect 276112 148996 276164 149048
rect 374276 148996 374328 149048
rect 434720 148996 434772 149048
rect 214840 148928 214892 148980
rect 274732 148928 274784 148980
rect 372344 148928 372396 148980
rect 401600 148928 401652 148980
rect 212172 148860 212224 148912
rect 241520 148860 241572 148912
rect 372160 148860 372212 148912
rect 373632 148860 373684 148912
rect 400220 148860 400272 148912
rect 213276 148792 213328 148844
rect 240140 148792 240192 148844
rect 49056 148588 49108 148640
rect 54944 148588 54996 148640
rect 81440 148588 81492 148640
rect 47768 148520 47820 148572
rect 53380 148520 53432 148572
rect 80060 148520 80112 148572
rect 46480 148452 46532 148504
rect 51908 148452 51960 148504
rect 78680 148452 78732 148504
rect 212908 148452 212960 148504
rect 213552 148452 213604 148504
rect 372528 148452 372580 148504
rect 374736 148452 374788 148504
rect 397460 148452 397512 148504
rect 56232 148384 56284 148436
rect 116216 148384 116268 148436
rect 376576 148384 376628 148436
rect 398840 148384 398892 148436
rect 53288 148316 53340 148368
rect 114652 148316 114704 148368
rect 215852 148316 215904 148368
rect 238760 148316 238812 148368
rect 371792 148316 371844 148368
rect 379980 148316 380032 148368
rect 429200 148316 429252 148368
rect 374276 148180 374328 148232
rect 375012 148180 375064 148232
rect 57796 147568 57848 147620
rect 104900 147568 104952 147620
rect 212080 147568 212132 147620
rect 215852 147568 215904 147620
rect 370964 147568 371016 147620
rect 376024 147568 376076 147620
rect 376576 147568 376628 147620
rect 378968 147568 379020 147620
rect 379428 147568 379480 147620
rect 426532 147568 426584 147620
rect 58624 147500 58676 147552
rect 103520 147500 103572 147552
rect 56140 147160 56192 147212
rect 58624 147160 58676 147212
rect 59912 146888 59964 146940
rect 107660 146888 107712 146940
rect 54208 146208 54260 146260
rect 58808 146208 58860 146260
rect 99380 146208 99432 146260
rect 179052 146208 179104 146260
rect 197544 146208 197596 146260
rect 217140 146208 217192 146260
rect 255412 146208 255464 146260
rect 276020 146208 276072 146260
rect 356612 146208 356664 146260
rect 358728 146208 358780 146260
rect 510620 146208 510672 146260
rect 56968 146140 57020 146192
rect 57244 146140 57296 146192
rect 59820 146140 59872 146192
rect 93860 146140 93912 146192
rect 179696 146140 179748 146192
rect 197636 146140 197688 146192
rect 219900 146140 219952 146192
rect 253940 146140 253992 146192
rect 338488 146140 338540 146192
rect 356888 146140 356940 146192
rect 374552 146140 374604 146192
rect 375656 146140 375708 146192
rect 377220 146140 377272 146192
rect 377956 146140 378008 146192
rect 378600 146140 378652 146192
rect 378968 146140 379020 146192
rect 379612 146140 379664 146192
rect 379796 146140 379848 146192
rect 414020 146140 414072 146192
rect 498660 146140 498712 146192
rect 517796 146140 517848 146192
rect 518072 146140 518124 146192
rect 91192 146072 91244 146124
rect 218796 146072 218848 146124
rect 219164 146072 219216 146124
rect 252560 146072 252612 146124
rect 340236 146072 340288 146124
rect 357440 146072 357492 146124
rect 374460 146072 374512 146124
rect 375104 146072 375156 146124
rect 53196 146004 53248 146056
rect 53840 146004 53892 146056
rect 86960 146004 87012 146056
rect 216772 146004 216824 146056
rect 56048 145936 56100 145988
rect 88432 145936 88484 145988
rect 54576 145868 54628 145920
rect 54852 145868 54904 145920
rect 85580 145868 85632 145920
rect 58900 145800 58952 145852
rect 89812 145800 89864 145852
rect 47584 145732 47636 145784
rect 52368 145732 52420 145784
rect 77300 145732 77352 145784
rect 251180 146004 251232 146056
rect 396724 146072 396776 146124
rect 416780 146072 416832 146124
rect 499856 146072 499908 146124
rect 517888 146072 517940 146124
rect 518440 146072 518492 146124
rect 409972 146004 410024 146056
rect 219072 145936 219124 145988
rect 251272 145936 251324 145988
rect 374368 145936 374420 145988
rect 378692 145936 378744 145988
rect 379244 145936 379296 145988
rect 411352 145936 411404 145988
rect 217876 145868 217928 145920
rect 249800 145868 249852 145920
rect 375748 145868 375800 145920
rect 407212 145868 407264 145920
rect 217876 145732 217928 145784
rect 218612 145732 218664 145784
rect 219256 145732 219308 145784
rect 224316 145800 224368 145852
rect 247132 145800 247184 145852
rect 375104 145800 375156 145852
rect 378968 145800 379020 145852
rect 408500 145800 408552 145852
rect 248420 145732 248472 145784
rect 402980 145732 403032 145784
rect 49240 145664 49292 145716
rect 54668 145664 54720 145716
rect 82820 145664 82872 145716
rect 216220 145664 216272 145716
rect 224132 145664 224184 145716
rect 224224 145664 224276 145716
rect 244280 145664 244332 145716
rect 375656 145664 375708 145716
rect 403072 145664 403124 145716
rect 56324 145596 56376 145648
rect 84292 145596 84344 145648
rect 216312 145596 216364 145648
rect 244372 145596 244424 145648
rect 280068 145596 280120 145648
rect 356612 145596 356664 145648
rect 357624 145596 357676 145648
rect 376576 145596 376628 145648
rect 404360 145596 404412 145648
rect 518440 145596 518492 145648
rect 580264 145596 580316 145648
rect 58808 145528 58860 145580
rect 91100 145528 91152 145580
rect 191748 145528 191800 145580
rect 198004 145528 198056 145580
rect 204904 145528 204956 145580
rect 214748 145528 214800 145580
rect 245660 145528 245712 145580
rect 351644 145528 351696 145580
rect 358728 145528 358780 145580
rect 375196 145528 375248 145580
rect 405740 145528 405792 145580
rect 518072 145528 518124 145580
rect 580356 145528 580408 145580
rect 58716 145460 58768 145512
rect 84200 145460 84252 145512
rect 214472 145460 214524 145512
rect 242900 145460 242952 145512
rect 375748 145460 375800 145512
rect 376484 145460 376536 145512
rect 378600 145460 378652 145512
rect 396080 145460 396132 145512
rect 47216 145392 47268 145444
rect 55036 145392 55088 145444
rect 76012 145392 76064 145444
rect 215576 145392 215628 145444
rect 218520 145392 218572 145444
rect 236092 145392 236144 145444
rect 378692 145392 378744 145444
rect 396172 145392 396224 145444
rect 46664 145324 46716 145376
rect 54760 145324 54812 145376
rect 75920 145324 75972 145376
rect 215116 145324 215168 145376
rect 219164 145324 219216 145376
rect 236000 145324 236052 145376
rect 378784 145324 378836 145376
rect 393320 145324 393372 145376
rect 49148 145256 49200 145308
rect 59912 145256 59964 145308
rect 377036 145256 377088 145308
rect 411260 145256 411312 145308
rect 215024 145188 215076 145240
rect 224224 145188 224276 145240
rect 54484 144848 54536 144900
rect 55956 144848 56008 144900
rect 56324 144848 56376 144900
rect 213644 144848 213696 144900
rect 214748 144848 214800 144900
rect 373172 144848 373224 144900
rect 375196 144848 375248 144900
rect 377956 144848 378008 144900
rect 421564 144848 421616 144900
rect 53104 144780 53156 144832
rect 55864 144780 55916 144832
rect 56416 144780 56468 144832
rect 213460 144780 213512 144832
rect 214656 144780 214708 144832
rect 375104 144780 375156 144832
rect 378600 144780 378652 144832
rect 52000 144712 52052 144764
rect 58716 144712 58768 144764
rect 212356 144712 212408 144764
rect 215852 144712 215904 144764
rect 373724 144712 373776 144764
rect 376208 144712 376260 144764
rect 376576 144712 376628 144764
rect 47952 144644 48004 144696
rect 58624 144644 58676 144696
rect 210700 144644 210752 144696
rect 214564 144644 214616 144696
rect 50344 144576 50396 144628
rect 58808 144576 58860 144628
rect 56140 144508 56192 144560
rect 56416 144508 56468 144560
rect 56232 144440 56284 144492
rect 56232 144236 56284 144288
rect 520188 79976 520240 80028
rect 580448 79976 580500 80028
rect 364984 70320 365036 70372
rect 376944 70320 376996 70372
rect 374644 68960 374696 69012
rect 377312 68960 377364 69012
rect 358728 68280 358780 68332
rect 376944 68280 376996 68332
rect 358084 68144 358136 68196
rect 358728 68144 358780 68196
rect 204904 67600 204956 67652
rect 216680 67600 216732 67652
rect 378692 59780 378744 59832
rect 397092 59780 397144 59832
rect 218520 59712 218572 59764
rect 237104 59712 237156 59764
rect 378600 59712 378652 59764
rect 396080 59712 396132 59764
rect 55036 59644 55088 59696
rect 77116 59644 77168 59696
rect 217140 59644 217192 59696
rect 255872 59644 255924 59696
rect 378048 59644 378100 59696
rect 416964 59644 417016 59696
rect 54668 59576 54720 59628
rect 83096 59576 83148 59628
rect 218428 59576 218480 59628
rect 261760 59576 261812 59628
rect 378784 59576 378836 59628
rect 418160 59576 418212 59628
rect 54208 59508 54260 59560
rect 99472 59508 99524 59560
rect 216404 59508 216456 59560
rect 260656 59508 260708 59560
rect 379336 59508 379388 59560
rect 422852 59508 422904 59560
rect 49608 59440 49660 59492
rect 113548 59440 113600 59492
rect 215208 59440 215260 59492
rect 259460 59440 259512 59492
rect 375932 59440 375984 59492
rect 423956 59440 424008 59492
rect 50896 59372 50948 59424
rect 120908 59372 120960 59424
rect 216036 59372 216088 59424
rect 263876 59372 263928 59424
rect 358176 59372 358228 59424
rect 418436 59372 418488 59424
rect 55956 59304 56008 59356
rect 84200 59304 84252 59356
rect 217968 59304 218020 59356
rect 358084 59304 358136 59356
rect 59820 59236 59872 59288
rect 94504 59236 94556 59288
rect 218888 59236 218940 59288
rect 256976 59236 257028 59288
rect 374552 59236 374604 59288
rect 403072 59236 403124 59288
rect 59084 59168 59136 59220
rect 95884 59168 95936 59220
rect 217784 59168 217836 59220
rect 258080 59168 258132 59220
rect 376668 59168 376720 59220
rect 421748 59168 421800 59220
rect 56508 59100 56560 59152
rect 98092 59100 98144 59152
rect 219624 59100 219676 59152
rect 265256 59100 265308 59152
rect 375288 59100 375340 59152
rect 420644 59100 420696 59152
rect 55864 59032 55916 59084
rect 100760 59032 100812 59084
rect 216128 59032 216180 59084
rect 262772 59032 262824 59084
rect 373264 59032 373316 59084
rect 425980 59032 426032 59084
rect 58532 58964 58584 59016
rect 102784 58964 102836 59016
rect 206928 58964 206980 59016
rect 295892 58964 295944 59016
rect 362224 58964 362276 59016
rect 423496 58964 423548 59016
rect 54392 58896 54444 58948
rect 101772 58896 101824 58948
rect 211620 58896 211672 58948
rect 303436 58896 303488 58948
rect 366364 58896 366416 58948
rect 453396 58896 453448 58948
rect 56232 58828 56284 58880
rect 116952 58828 117004 58880
rect 201408 58828 201460 58880
rect 298468 58828 298520 58880
rect 360844 58828 360896 58880
rect 463516 58828 463568 58880
rect 53012 58760 53064 58812
rect 113272 58760 113324 58812
rect 198648 58760 198700 58812
rect 315856 58760 315908 58812
rect 366456 58760 366508 58812
rect 480904 58760 480956 58812
rect 50068 58692 50120 58744
rect 148508 58692 148560 58744
rect 206836 58692 206888 58744
rect 323308 58692 323360 58744
rect 361488 58692 361540 58744
rect 485964 58692 486016 58744
rect 52828 58624 52880 58676
rect 150900 58624 150952 58676
rect 219256 58624 219308 58676
rect 428188 58624 428240 58676
rect 374460 58556 374512 58608
rect 404176 58556 404228 58608
rect 57888 57876 57940 57928
rect 204904 57876 204956 57928
rect 208308 57876 208360 57928
rect 325884 57876 325936 57928
rect 343180 57876 343232 57928
rect 357532 57876 357584 57928
rect 364248 57876 364300 57928
rect 478420 57876 478472 57928
rect 503260 57876 503312 57928
rect 517612 57876 517664 57928
rect 51448 57808 51500 57860
rect 145564 57808 145616 57860
rect 183284 57808 183336 57860
rect 197452 57808 197504 57860
rect 211068 57808 211120 57860
rect 318340 57808 318392 57860
rect 343456 57808 343508 57860
rect 356704 57808 356756 57860
rect 378508 57808 378560 57860
rect 470876 57808 470928 57860
rect 503536 57808 503588 57860
rect 517520 57808 517572 57860
rect 41236 57740 41288 57792
rect 133420 57740 133472 57792
rect 183468 57740 183520 57792
rect 197360 57740 197412 57792
rect 205548 57740 205600 57792
rect 310980 57740 311032 57792
rect 363604 57740 363656 57792
rect 443460 57740 443512 57792
rect 41144 57672 41196 57724
rect 123484 57672 123536 57724
rect 218980 57672 219032 57724
rect 320916 57672 320968 57724
rect 367928 57672 367980 57724
rect 448244 57672 448296 57724
rect 53748 57604 53800 57656
rect 130844 57604 130896 57656
rect 213736 57604 213788 57656
rect 313372 57604 313424 57656
rect 367836 57604 367888 57656
rect 440884 57604 440936 57656
rect 57244 57536 57296 57588
rect 57888 57536 57940 57588
rect 55128 57468 55180 57520
rect 128360 57536 128412 57588
rect 209688 57536 209740 57588
rect 305828 57536 305880 57588
rect 363696 57536 363748 57588
rect 433616 57536 433668 57588
rect 58992 57468 59044 57520
rect 125876 57468 125928 57520
rect 218336 57468 218388 57520
rect 300860 57468 300912 57520
rect 370504 57468 370556 57520
rect 438492 57468 438544 57520
rect 52092 57400 52144 57452
rect 111156 57400 111208 57452
rect 279056 57400 279108 57452
rect 356612 57400 356664 57452
rect 371884 57400 371936 57452
rect 435916 57400 435968 57452
rect 51540 57332 51592 57384
rect 88340 57332 88392 57384
rect 216496 57332 216548 57384
rect 293316 57332 293368 57384
rect 376116 57332 376168 57384
rect 430948 57332 431000 57384
rect 58348 57264 58400 57316
rect 58992 57264 59044 57316
rect 59268 57264 59320 57316
rect 90732 57264 90784 57316
rect 216588 57264 216640 57316
rect 287612 57264 287664 57316
rect 365076 57264 365128 57316
rect 416044 57264 416096 57316
rect 52368 57196 52420 57248
rect 78220 57196 78272 57248
rect 218704 57196 218756 57248
rect 265348 57196 265400 57248
rect 379704 57196 379756 57248
rect 415492 57196 415544 57248
rect 54760 57128 54812 57180
rect 76012 57128 76064 57180
rect 213828 57128 213880 57180
rect 283656 57128 283708 57180
rect 54944 56516 54996 56568
rect 81808 56516 81860 56568
rect 214472 56516 214524 56568
rect 242900 56516 242952 56568
rect 376024 56516 376076 56568
rect 399484 56516 399536 56568
rect 53472 56448 53524 56500
rect 109224 56448 109276 56500
rect 215944 56448 215996 56500
rect 239220 56448 239272 56500
rect 372252 56448 372304 56500
rect 435732 56448 435784 56500
rect 59912 56380 59964 56432
rect 108028 56380 108080 56432
rect 219164 56380 219216 56432
rect 236000 56380 236052 56432
rect 378416 56380 378468 56432
rect 438216 56380 438268 56432
rect 57796 56312 57848 56364
rect 104992 56312 105044 56364
rect 214932 56312 214984 56364
rect 269764 56312 269816 56364
rect 374920 56312 374972 56364
rect 432236 56312 432288 56364
rect 59176 56244 59228 56296
rect 106740 56244 106792 56296
rect 218244 56244 218296 56296
rect 267004 56244 267056 56296
rect 379428 56244 379480 56296
rect 427636 56244 427688 56296
rect 56416 56176 56468 56228
rect 103796 56176 103848 56228
rect 219808 56176 219860 56228
rect 266360 56176 266412 56228
rect 379888 56176 379940 56228
rect 426440 56176 426492 56228
rect 60004 56108 60056 56160
rect 106372 56108 106424 56160
rect 218796 56108 218848 56160
rect 253388 56108 253440 56160
rect 379796 56108 379848 56160
rect 414572 56108 414624 56160
rect 58808 56040 58860 56092
rect 92112 56040 92164 56092
rect 219072 56040 219124 56092
rect 251180 56040 251232 56092
rect 378876 56040 378928 56092
rect 412640 56040 412692 56092
rect 56324 55972 56376 56024
rect 88708 55972 88760 56024
rect 214748 55972 214800 56024
rect 246396 55972 246448 56024
rect 379152 55972 379204 56024
rect 411260 55972 411312 56024
rect 54852 55904 54904 55956
rect 86500 55904 86552 55956
rect 218612 55904 218664 55956
rect 248604 55904 248656 55956
rect 378968 55904 379020 55956
rect 408684 55904 408736 55956
rect 58716 55836 58768 55888
rect 85396 55836 85448 55888
rect 213368 55836 213420 55888
rect 273628 55836 273680 55888
rect 372344 55836 372396 55888
rect 401692 55836 401744 55888
rect 53564 55768 53616 55820
rect 115756 55768 115808 55820
rect 219992 55768 220044 55820
rect 408316 55768 408368 55820
rect 51908 55700 51960 55752
rect 79508 55700 79560 55752
rect 215852 55700 215904 55752
rect 272156 55700 272208 55752
rect 44088 55156 44140 55208
rect 115940 55156 115992 55208
rect 213552 55156 213604 55208
rect 274640 55156 274692 55208
rect 376392 55156 376444 55208
rect 436100 55156 436152 55208
rect 53288 55088 53340 55140
rect 113180 55088 113232 55140
rect 214840 55088 214892 55140
rect 273352 55088 273404 55140
rect 375012 55088 375064 55140
rect 433340 55088 433392 55140
rect 52184 55020 52236 55072
rect 111800 55020 111852 55072
rect 214656 55020 214708 55072
rect 270500 55020 270552 55072
rect 375564 55020 375616 55072
rect 433432 55020 433484 55072
rect 58624 54952 58676 55004
rect 92480 54952 92532 55004
rect 219532 54952 219584 55004
rect 267740 54952 267792 55004
rect 374828 54952 374880 55004
rect 430580 54952 430632 55004
rect 56968 54884 57020 54936
rect 91192 54884 91244 54936
rect 219900 54884 219952 54936
rect 253940 54884 253992 54936
rect 376300 54884 376352 54936
rect 429200 54884 429252 54936
rect 53196 54816 53248 54868
rect 86960 54816 87012 54868
rect 217876 54816 217928 54868
rect 251364 54816 251416 54868
rect 379980 54816 380032 54868
rect 427820 54816 427872 54868
rect 58900 54748 58952 54800
rect 89720 54748 89772 54800
rect 216220 54748 216272 54800
rect 247040 54748 247092 54800
rect 377036 54748 377088 54800
rect 411352 54748 411404 54800
rect 53380 54680 53432 54732
rect 80060 54680 80112 54732
rect 212172 54680 212224 54732
rect 241520 54680 241572 54732
rect 377220 54680 377272 54732
rect 409880 54680 409932 54732
rect 215024 54612 215076 54664
rect 244280 54612 244332 54664
rect 375104 54612 375156 54664
rect 405832 54612 405884 54664
rect 216312 54544 216364 54596
rect 244372 54544 244424 54596
rect 376576 54544 376628 54596
rect 407212 54544 407264 54596
rect 213276 54476 213328 54528
rect 240140 54476 240192 54528
rect 376208 54476 376260 54528
rect 404360 54476 404412 54528
rect 214564 54408 214616 54460
rect 237380 54408 237432 54460
rect 372160 54408 372212 54460
rect 400220 54408 400272 54460
rect 374736 54340 374788 54392
rect 397460 54340 397512 54392
rect 2780 20340 2832 20392
rect 4804 20340 4856 20392
rect 572 3408 624 3460
rect 57244 3408 57296 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 639606 3464 684247
rect 3424 639600 3476 639606
rect 3424 639542 3476 639548
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 561134 3464 579935
rect 3424 561128 3476 561134
rect 3424 561070 3476 561076
rect 3424 559564 3476 559570
rect 3424 559506 3476 559512
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 58585 3464 559506
rect 3528 555490 3556 632023
rect 18604 630760 18656 630766
rect 18604 630702 18656 630708
rect 4804 556844 4856 556850
rect 4804 556786 4856 556792
rect 3516 555484 3568 555490
rect 3516 555426 3568 555432
rect 3516 553444 3568 553450
rect 3516 553386 3568 553392
rect 3528 97617 3556 553386
rect 3608 540116 3660 540122
rect 3608 540058 3660 540064
rect 3620 514865 3648 540058
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3608 476808 3660 476814
rect 3608 476750 3660 476756
rect 3620 462641 3648 476750
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 4816 20398 4844 556786
rect 15844 468512 15896 468518
rect 15844 468454 15896 468460
rect 15856 411262 15884 468454
rect 15844 411256 15896 411262
rect 15844 411198 15896 411204
rect 18616 358766 18644 630702
rect 40052 549234 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 57888 700324 57940 700330
rect 57888 700266 57940 700272
rect 40682 632088 40738 632097
rect 40682 632023 40738 632032
rect 40040 549228 40092 549234
rect 40040 549170 40092 549176
rect 40592 462868 40644 462874
rect 40592 462810 40644 462816
rect 40604 373289 40632 462810
rect 40590 373280 40646 373289
rect 40590 373215 40646 373224
rect 18604 358760 18656 358766
rect 18604 358702 18656 358708
rect 40696 202842 40724 632023
rect 54852 625320 54904 625326
rect 54852 625262 54904 625268
rect 54864 559774 54892 625262
rect 55128 625252 55180 625258
rect 55128 625194 55180 625200
rect 54944 622600 54996 622606
rect 54944 622542 54996 622548
rect 54852 559768 54904 559774
rect 54852 559710 54904 559716
rect 54956 543250 54984 622542
rect 55036 622464 55088 622470
rect 55036 622406 55088 622412
rect 55048 543590 55076 622406
rect 55140 543658 55168 625194
rect 56508 625184 56560 625190
rect 56508 625126 56560 625132
rect 56324 622668 56376 622674
rect 56324 622610 56376 622616
rect 55128 543652 55180 543658
rect 55128 543594 55180 543600
rect 55036 543584 55088 543590
rect 55036 543526 55088 543532
rect 56336 543318 56364 622610
rect 56416 622532 56468 622538
rect 56416 622474 56468 622480
rect 56324 543312 56376 543318
rect 56324 543254 56376 543260
rect 54944 543244 54996 543250
rect 54944 543186 54996 543192
rect 56428 543182 56456 622474
rect 56520 543386 56548 625126
rect 57796 623892 57848 623898
rect 57796 623834 57848 623840
rect 57702 620664 57758 620673
rect 57702 620599 57758 620608
rect 57518 614408 57574 614417
rect 57518 614343 57574 614352
rect 57426 589928 57482 589937
rect 57426 589863 57482 589872
rect 57334 586392 57390 586401
rect 57334 586327 57390 586336
rect 57058 577688 57114 577697
rect 57058 577623 57114 577632
rect 57072 559910 57100 577623
rect 57150 574968 57206 574977
rect 57150 574903 57206 574912
rect 57164 560250 57192 574903
rect 57348 572354 57376 586327
rect 57336 572348 57388 572354
rect 57336 572290 57388 572296
rect 57334 571568 57390 571577
rect 57334 571503 57390 571512
rect 57242 565448 57298 565457
rect 57242 565383 57298 565392
rect 57152 560244 57204 560250
rect 57152 560186 57204 560192
rect 57060 559904 57112 559910
rect 57060 559846 57112 559852
rect 57256 545834 57284 565383
rect 57348 557054 57376 571503
rect 57440 558890 57468 589863
rect 57532 583778 57560 614343
rect 57610 593464 57666 593473
rect 57610 593399 57666 593408
rect 57520 583772 57572 583778
rect 57520 583714 57572 583720
rect 57518 583672 57574 583681
rect 57518 583607 57574 583616
rect 57428 558884 57480 558890
rect 57428 558826 57480 558832
rect 57336 557048 57388 557054
rect 57336 556990 57388 556996
rect 57532 551478 57560 583607
rect 57520 551472 57572 551478
rect 57520 551414 57572 551420
rect 57624 547398 57652 593399
rect 57716 552770 57744 620599
rect 57704 552764 57756 552770
rect 57704 552706 57756 552712
rect 57612 547392 57664 547398
rect 57612 547334 57664 547340
rect 57244 545828 57296 545834
rect 57244 545770 57296 545776
rect 57808 543522 57836 623834
rect 57900 599593 57928 700266
rect 104912 638246 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 137928 683188 137980 683194
rect 137928 683130 137980 683136
rect 104900 638240 104952 638246
rect 104900 638182 104952 638188
rect 100576 625728 100628 625734
rect 100576 625670 100628 625676
rect 124312 625728 124364 625734
rect 124312 625670 124364 625676
rect 137836 625728 137888 625734
rect 137836 625670 137888 625676
rect 94780 625592 94832 625598
rect 94780 625534 94832 625540
rect 83188 625524 83240 625530
rect 83188 625466 83240 625472
rect 77392 625184 77444 625190
rect 77392 625126 77444 625132
rect 59360 623960 59412 623966
rect 59360 623902 59412 623908
rect 59266 617808 59322 617817
rect 59266 617743 59322 617752
rect 59082 611688 59138 611697
rect 59082 611623 59138 611632
rect 58898 608288 58954 608297
rect 58898 608223 58954 608232
rect 57886 599584 57942 599593
rect 57886 599519 57942 599528
rect 57886 596048 57942 596057
rect 57886 595983 57942 595992
rect 57900 561202 57928 595983
rect 58624 583772 58676 583778
rect 58624 583714 58676 583720
rect 58530 568848 58586 568857
rect 58530 568783 58586 568792
rect 57888 561196 57940 561202
rect 57888 561138 57940 561144
rect 57796 543516 57848 543522
rect 57796 543458 57848 543464
rect 56508 543380 56560 543386
rect 56508 543322 56560 543328
rect 56416 543176 56468 543182
rect 56416 543118 56468 543124
rect 57900 509969 57928 561138
rect 58544 554130 58572 568783
rect 58532 554124 58584 554130
rect 58532 554066 58584 554072
rect 58636 543046 58664 583714
rect 58806 581088 58862 581097
rect 58806 581023 58862 581032
rect 58716 572348 58768 572354
rect 58716 572290 58768 572296
rect 58728 543454 58756 572290
rect 58716 543448 58768 543454
rect 58716 543390 58768 543396
rect 58820 543114 58848 581023
rect 58912 558210 58940 608223
rect 58990 602168 59046 602177
rect 58990 602103 59046 602112
rect 58900 558204 58952 558210
rect 58900 558146 58952 558152
rect 59004 551410 59032 602103
rect 59096 559842 59124 611623
rect 59174 605568 59230 605577
rect 59174 605503 59230 605512
rect 59084 559836 59136 559842
rect 59084 559778 59136 559784
rect 58992 551404 59044 551410
rect 58992 551346 59044 551352
rect 59188 548554 59216 605503
rect 59280 555626 59308 617743
rect 59268 555620 59320 555626
rect 59268 555562 59320 555568
rect 59176 548548 59228 548554
rect 59176 548490 59228 548496
rect 59372 547874 59400 623902
rect 69020 623824 69072 623830
rect 69020 623766 69072 623772
rect 69032 623084 69060 623766
rect 77404 623084 77432 625126
rect 80612 623892 80664 623898
rect 80612 623834 80664 623840
rect 80624 623084 80652 623834
rect 83200 623084 83228 625466
rect 88984 625320 89036 625326
rect 88984 625262 89036 625268
rect 86408 623892 86460 623898
rect 86408 623834 86460 623840
rect 86420 623084 86448 623834
rect 88996 623084 89024 625262
rect 92204 625252 92256 625258
rect 92204 625194 92256 625200
rect 92216 623084 92244 625194
rect 94792 623084 94820 625534
rect 98000 623960 98052 623966
rect 98000 623902 98052 623908
rect 98012 623084 98040 623902
rect 100588 623084 100616 625670
rect 112168 625660 112220 625666
rect 112168 625602 112220 625608
rect 122840 625660 122892 625666
rect 122840 625602 122892 625608
rect 109592 625456 109644 625462
rect 109592 625398 109644 625404
rect 103796 625388 103848 625394
rect 103796 625330 103848 625336
rect 103808 623084 103836 625330
rect 106370 625288 106426 625297
rect 106370 625223 106426 625232
rect 106384 623084 106412 625223
rect 109604 623084 109632 625398
rect 112180 623084 112208 625602
rect 122288 625592 122340 625598
rect 122288 625534 122340 625540
rect 120908 625456 120960 625462
rect 120908 625398 120960 625404
rect 115388 625252 115440 625258
rect 115388 625194 115440 625200
rect 115400 623084 115428 625194
rect 74644 622674 74842 622690
rect 74632 622668 74842 622674
rect 74684 622662 74842 622668
rect 74632 622610 74684 622616
rect 65524 622600 65576 622606
rect 65576 622548 65826 622554
rect 65524 622542 65826 622548
rect 65536 622526 65826 622542
rect 71240 622538 71622 622554
rect 71228 622532 71622 622538
rect 71280 622526 71622 622532
rect 71228 622474 71280 622480
rect 62948 622464 63000 622470
rect 59464 622390 60030 622418
rect 63000 622412 63250 622418
rect 62948 622406 63250 622412
rect 62960 622390 63250 622406
rect 117990 622402 118280 622418
rect 117990 622396 118292 622402
rect 117990 622390 118240 622396
rect 59464 552906 59492 622390
rect 120566 622390 120764 622418
rect 118240 622338 118292 622344
rect 59542 562788 59598 562797
rect 59542 562723 59598 562732
rect 59452 552900 59504 552906
rect 59452 552842 59504 552848
rect 59556 550050 59584 562723
rect 62120 560244 62172 560250
rect 62120 560186 62172 560192
rect 60030 560102 60320 560130
rect 60292 558754 60320 560102
rect 60740 558884 60792 558890
rect 60740 558826 60792 558832
rect 60280 558748 60332 558754
rect 60280 558690 60332 558696
rect 60752 557534 60780 558826
rect 62132 557534 62160 560186
rect 62606 560102 62896 560130
rect 62764 558748 62816 558754
rect 62764 558690 62816 558696
rect 60752 557506 60964 557534
rect 62132 557506 62436 557534
rect 59544 550044 59596 550050
rect 59544 549986 59596 549992
rect 59372 547846 60320 547874
rect 58808 543108 58860 543114
rect 58808 543050 58860 543056
rect 58624 543040 58676 543046
rect 58624 542982 58676 542988
rect 60292 539963 60320 547846
rect 60936 539963 60964 557506
rect 61660 543720 61712 543726
rect 61660 543662 61712 543668
rect 61672 539963 61700 543662
rect 62408 539963 62436 557506
rect 62776 547262 62804 558690
rect 62868 558346 62896 560102
rect 65076 560102 65182 560130
rect 68402 560102 68784 560130
rect 70978 560102 71360 560130
rect 63500 559632 63552 559638
rect 63500 559574 63552 559580
rect 62856 558340 62908 558346
rect 62856 558282 62908 558288
rect 62764 547256 62816 547262
rect 62764 547198 62816 547204
rect 63132 547188 63184 547194
rect 63132 547130 63184 547136
rect 63144 539963 63172 547130
rect 63512 543930 63540 559574
rect 65076 557598 65104 560102
rect 67732 559904 67784 559910
rect 67732 559846 67784 559852
rect 67640 559700 67692 559706
rect 67640 559642 67692 559648
rect 64144 557592 64196 557598
rect 64144 557534 64196 557540
rect 65064 557592 65116 557598
rect 65064 557534 65116 557540
rect 63776 556912 63828 556918
rect 63776 556854 63828 556860
rect 63500 543924 63552 543930
rect 63500 543866 63552 543872
rect 63788 539963 63816 556854
rect 64156 543726 64184 557534
rect 64880 555552 64932 555558
rect 64880 555494 64932 555500
rect 64512 543924 64564 543930
rect 64892 543912 64920 555494
rect 66720 554056 66772 554062
rect 66720 553998 66772 554004
rect 65984 551336 66036 551342
rect 65984 551278 66036 551284
rect 64892 543884 65288 543912
rect 64512 543866 64564 543872
rect 64144 543720 64196 543726
rect 64144 543662 64196 543668
rect 64524 539963 64552 543866
rect 65260 539963 65288 543884
rect 65996 539963 66024 551278
rect 66732 539963 66760 553998
rect 67652 543912 67680 559642
rect 67744 557534 67772 559846
rect 68756 558482 68784 560102
rect 68744 558476 68796 558482
rect 68744 558418 68796 558424
rect 71044 558476 71096 558482
rect 71044 558418 71096 558424
rect 67744 557506 68876 557534
rect 67652 543884 68140 543912
rect 67364 543652 67416 543658
rect 67364 543594 67416 543600
rect 67376 539963 67404 543594
rect 68112 539963 68140 543884
rect 68848 539963 68876 557506
rect 69020 552696 69072 552702
rect 69020 552638 69072 552644
rect 69032 543912 69060 552638
rect 69112 550180 69164 550186
rect 69112 550122 69164 550128
rect 69124 544066 69152 550122
rect 70952 549976 71004 549982
rect 70952 549918 71004 549924
rect 69112 544060 69164 544066
rect 69112 544002 69164 544008
rect 70308 544060 70360 544066
rect 70308 544002 70360 544008
rect 69032 543884 69612 543912
rect 69584 539963 69612 543884
rect 70320 539963 70348 544002
rect 70964 539963 70992 549918
rect 71056 544406 71084 558418
rect 71332 558278 71360 560102
rect 73816 560102 74198 560130
rect 76774 560102 77064 560130
rect 71320 558272 71372 558278
rect 71320 558214 71372 558220
rect 73816 557938 73844 560102
rect 77036 558414 77064 560102
rect 79888 560102 79994 560130
rect 82570 560102 82768 560130
rect 85790 560102 86080 560130
rect 88366 560102 88656 560130
rect 78680 559768 78732 559774
rect 78680 559710 78732 559716
rect 77024 558408 77076 558414
rect 77024 558350 77076 558356
rect 74540 558204 74592 558210
rect 74540 558146 74592 558152
rect 71780 557932 71832 557938
rect 71780 557874 71832 557880
rect 73804 557932 73856 557938
rect 73804 557874 73856 557880
rect 71792 557534 71820 557874
rect 71792 557506 72464 557534
rect 71688 545760 71740 545766
rect 71688 545702 71740 545708
rect 71044 544400 71096 544406
rect 71044 544342 71096 544348
rect 71700 539963 71728 545702
rect 72436 539963 72464 557506
rect 73252 554192 73304 554198
rect 73252 554134 73304 554140
rect 73264 540138 73292 554134
rect 73804 543176 73856 543182
rect 73804 543118 73856 543124
rect 73188 540110 73292 540138
rect 73188 539920 73216 540110
rect 73816 539963 73844 543118
rect 74552 539963 74580 558146
rect 75920 552900 75972 552906
rect 75920 552842 75972 552848
rect 75276 552832 75328 552838
rect 75276 552774 75328 552780
rect 75288 539963 75316 552774
rect 75932 543946 75960 552842
rect 77392 552764 77444 552770
rect 77392 552706 77444 552712
rect 76748 548616 76800 548622
rect 76748 548558 76800 548564
rect 75932 543918 76052 543946
rect 76024 539963 76052 543918
rect 76760 539963 76788 548558
rect 77404 539963 77432 552706
rect 78692 543930 78720 559710
rect 79888 558210 79916 560102
rect 82740 558482 82768 560102
rect 82912 559836 82964 559842
rect 82912 559778 82964 559784
rect 82728 558476 82780 558482
rect 82728 558418 82780 558424
rect 80704 558340 80756 558346
rect 80704 558282 80756 558288
rect 79876 558204 79928 558210
rect 79876 558146 79928 558152
rect 78864 556980 78916 556986
rect 78864 556922 78916 556928
rect 78680 543924 78732 543930
rect 78680 543866 78732 543872
rect 78128 543176 78180 543182
rect 78128 543118 78180 543124
rect 78140 539963 78168 543118
rect 78876 539963 78904 556922
rect 80060 552764 80112 552770
rect 80060 552706 80112 552712
rect 80072 543946 80100 552706
rect 80716 550118 80744 558282
rect 82924 557534 82952 559778
rect 85580 559768 85632 559774
rect 85580 559710 85632 559716
rect 82924 557506 83228 557534
rect 81716 557048 81768 557054
rect 81716 556990 81768 556996
rect 80980 551540 81032 551546
rect 80980 551482 81032 551488
rect 80704 550112 80756 550118
rect 80704 550054 80756 550060
rect 79600 543924 79652 543930
rect 80072 543918 80376 543946
rect 79600 543866 79652 543872
rect 79612 539963 79640 543866
rect 80348 539963 80376 543918
rect 80992 539963 81020 551482
rect 81728 539963 81756 556990
rect 82452 545896 82504 545902
rect 82452 545838 82504 545844
rect 82464 539963 82492 545838
rect 83200 539963 83228 557506
rect 84568 547324 84620 547330
rect 84568 547266 84620 547272
rect 83924 543380 83976 543386
rect 83924 543322 83976 543328
rect 83936 539963 83964 543322
rect 84580 539963 84608 547266
rect 85592 543946 85620 559710
rect 85672 558408 85724 558414
rect 85672 558350 85724 558356
rect 85684 557534 85712 558350
rect 86052 558346 86080 560102
rect 87052 559836 87104 559842
rect 87052 559778 87104 559784
rect 86958 559600 87014 559609
rect 86958 559535 87014 559544
rect 86040 558340 86092 558346
rect 86040 558282 86092 558288
rect 85684 557506 86816 557534
rect 85592 543918 86080 543946
rect 85304 543380 85356 543386
rect 85304 543322 85356 543328
rect 85316 539963 85344 543322
rect 86052 539963 86080 543918
rect 86788 539963 86816 557506
rect 86972 543946 87000 559535
rect 87064 557534 87092 559778
rect 87064 557506 88196 557534
rect 86972 543918 87460 543946
rect 87432 539963 87460 543918
rect 88168 539963 88196 557506
rect 88628 552906 88656 560102
rect 91112 560102 91586 560130
rect 94162 560102 94544 560130
rect 88984 558476 89036 558482
rect 88984 558418 89036 558424
rect 88616 552900 88668 552906
rect 88616 552842 88668 552848
rect 88432 548684 88484 548690
rect 88432 548626 88484 548632
rect 88444 543930 88472 548626
rect 88432 543924 88484 543930
rect 88432 543866 88484 543872
rect 88996 543726 89024 558418
rect 89812 551472 89864 551478
rect 89812 551414 89864 551420
rect 89824 543930 89852 551414
rect 89628 543924 89680 543930
rect 89628 543866 89680 543872
rect 89812 543924 89864 543930
rect 89812 543866 89864 543872
rect 91008 543924 91060 543930
rect 91008 543866 91060 543872
rect 88984 543720 89036 543726
rect 88984 543662 89036 543668
rect 88892 543584 88944 543590
rect 88892 543526 88944 543532
rect 88904 539963 88932 543526
rect 89640 539963 89668 543866
rect 90364 543720 90416 543726
rect 90364 543662 90416 543668
rect 90376 539963 90404 543662
rect 91020 539963 91048 543866
rect 91112 543590 91140 560102
rect 93860 559904 93912 559910
rect 93860 559846 93912 559852
rect 92572 555620 92624 555626
rect 92572 555562 92624 555568
rect 91744 547392 91796 547398
rect 91744 547334 91796 547340
rect 91100 543584 91152 543590
rect 91100 543526 91152 543532
rect 91756 539963 91784 547334
rect 92584 540138 92612 555562
rect 93872 547874 93900 559846
rect 94516 558414 94544 560102
rect 97000 560102 97382 560130
rect 99958 560102 100248 560130
rect 96804 559972 96856 559978
rect 96804 559914 96856 559920
rect 94504 558408 94556 558414
rect 94504 558350 94556 558356
rect 93952 558272 94004 558278
rect 93952 558214 94004 558220
rect 93964 551478 93992 558214
rect 93952 551472 94004 551478
rect 93952 551414 94004 551420
rect 96816 547874 96844 559914
rect 97000 552838 97028 560102
rect 98092 560040 98144 560046
rect 98092 559982 98144 559988
rect 98104 557534 98132 559982
rect 100220 558278 100248 560102
rect 102888 560102 103178 560130
rect 104912 560102 105754 560130
rect 106280 560108 106332 560114
rect 102888 558822 102916 560102
rect 100760 558816 100812 558822
rect 100760 558758 100812 558764
rect 102876 558816 102928 558822
rect 102876 558758 102928 558764
rect 100208 558272 100260 558278
rect 100208 558214 100260 558220
rect 98104 557506 98224 557534
rect 96988 552832 97040 552838
rect 96988 552774 97040 552780
rect 93872 547846 93992 547874
rect 96816 547846 97488 547874
rect 93216 543516 93268 543522
rect 93216 543458 93268 543464
rect 92508 540110 92612 540138
rect 92508 539920 92536 540110
rect 93228 539963 93256 543458
rect 93964 539963 93992 547846
rect 94596 544468 94648 544474
rect 94596 544410 94648 544416
rect 94608 539963 94636 544410
rect 96804 543584 96856 543590
rect 96804 543526 96856 543532
rect 95332 543448 95384 543454
rect 95332 543390 95384 543396
rect 96068 543448 96120 543454
rect 96068 543390 96120 543396
rect 95344 539963 95372 543390
rect 96080 539963 96108 543390
rect 96816 539963 96844 543526
rect 97460 539963 97488 547846
rect 98196 539963 98224 557506
rect 100392 555620 100444 555626
rect 100392 555562 100444 555568
rect 99656 543312 99708 543318
rect 99656 543254 99708 543260
rect 98920 543244 98972 543250
rect 98920 543186 98972 543192
rect 98932 539963 98960 543186
rect 99668 539963 99696 543254
rect 100404 539963 100432 555562
rect 100772 543930 100800 558758
rect 104164 558408 104216 558414
rect 104164 558350 104216 558356
rect 103520 552900 103572 552906
rect 103520 552842 103572 552848
rect 102508 551404 102560 551410
rect 102508 551346 102560 551352
rect 101036 550044 101088 550050
rect 101036 549986 101088 549992
rect 100760 543924 100812 543930
rect 100760 543866 100812 543872
rect 101048 539963 101076 549986
rect 101772 543924 101824 543930
rect 101772 543866 101824 543872
rect 101784 539963 101812 543866
rect 102520 539963 102548 551346
rect 103244 545828 103296 545834
rect 103244 545770 103296 545776
rect 103256 539963 103284 545770
rect 103532 543946 103560 552842
rect 104176 544066 104204 558350
rect 104912 548690 104940 560102
rect 106280 560050 106332 560056
rect 108592 560102 108974 560130
rect 110524 560102 111550 560130
rect 114664 560102 114770 560130
rect 117346 560102 117452 560130
rect 104900 548684 104952 548690
rect 104900 548626 104952 548632
rect 105360 547256 105412 547262
rect 105360 547198 105412 547204
rect 104164 544060 104216 544066
rect 104164 544002 104216 544008
rect 103532 543918 104664 543946
rect 103980 543244 104032 543250
rect 103980 543186 104032 543192
rect 103992 539963 104020 543186
rect 104636 539963 104664 543918
rect 105372 539963 105400 547198
rect 106292 543930 106320 560050
rect 108304 558340 108356 558346
rect 108304 558282 108356 558288
rect 106924 552900 106976 552906
rect 106924 552842 106976 552848
rect 106280 543924 106332 543930
rect 106280 543866 106332 543872
rect 106096 543720 106148 543726
rect 106096 543662 106148 543668
rect 106108 539963 106136 543662
rect 106936 543454 106964 552842
rect 108212 548548 108264 548554
rect 108212 548490 108264 548496
rect 107568 543924 107620 543930
rect 107568 543866 107620 543872
rect 106924 543448 106976 543454
rect 106924 543390 106976 543396
rect 106832 543312 106884 543318
rect 106832 543254 106884 543260
rect 106844 539963 106872 543254
rect 107580 539963 107608 543866
rect 108224 539963 108252 548490
rect 108316 543726 108344 558282
rect 108592 554198 108620 560102
rect 108580 554192 108632 554198
rect 108580 554134 108632 554140
rect 110420 554124 110472 554130
rect 110420 554066 110472 554072
rect 109684 550112 109736 550118
rect 109684 550054 109736 550060
rect 108948 544400 109000 544406
rect 108948 544342 109000 544348
rect 108304 543720 108356 543726
rect 108304 543662 108356 543668
rect 108960 539963 108988 544342
rect 109696 539963 109724 550054
rect 110432 543946 110460 554066
rect 110524 547194 110552 560102
rect 111892 558408 111944 558414
rect 111892 558350 111944 558356
rect 111904 547874 111932 558350
rect 112444 558340 112496 558346
rect 112444 558282 112496 558288
rect 112456 548622 112484 558282
rect 114560 558204 114612 558210
rect 114560 558146 114612 558152
rect 112444 548616 112496 548622
rect 112444 548558 112496 548564
rect 111904 547846 112576 547874
rect 110512 547188 110564 547194
rect 110512 547130 110564 547136
rect 110432 543918 111104 543946
rect 110420 543584 110472 543590
rect 110420 543526 110472 543532
rect 110432 539963 110460 543526
rect 111076 539963 111104 543918
rect 111800 543720 111852 543726
rect 111800 543662 111852 543668
rect 111812 539963 111840 543662
rect 112548 539963 112576 547846
rect 113272 544060 113324 544066
rect 113272 544002 113324 544008
rect 113284 539963 113312 544002
rect 114572 543930 114600 558146
rect 114664 552702 114692 560102
rect 116584 558816 116636 558822
rect 116584 558758 116636 558764
rect 115204 558272 115256 558278
rect 115204 558214 115256 558220
rect 114652 552696 114704 552702
rect 114652 552638 114704 552644
rect 114652 551472 114704 551478
rect 114652 551414 114704 551420
rect 114560 543924 114612 543930
rect 114560 543866 114612 543872
rect 114008 543448 114060 543454
rect 114008 543390 114060 543396
rect 114020 539963 114048 543390
rect 114664 539963 114692 551414
rect 115216 543726 115244 558214
rect 116596 545902 116624 558758
rect 117424 558346 117452 560102
rect 120184 560102 120566 560130
rect 120184 558822 120212 560102
rect 120172 558816 120224 558822
rect 120172 558758 120224 558764
rect 120736 558754 120764 622390
rect 120814 598360 120870 598369
rect 120814 598295 120870 598304
rect 119344 558748 119396 558754
rect 119344 558690 119396 558696
rect 120724 558748 120776 558754
rect 120724 558690 120776 558696
rect 117412 558340 117464 558346
rect 117412 558282 117464 558288
rect 118700 558340 118752 558346
rect 118700 558282 118752 558288
rect 116584 545896 116636 545902
rect 116584 545838 116636 545844
rect 115388 543924 115440 543930
rect 115388 543866 115440 543872
rect 115204 543720 115256 543726
rect 115204 543662 115256 543668
rect 115400 539963 115428 543866
rect 116124 543720 116176 543726
rect 116124 543662 116176 543668
rect 116136 539963 116164 543662
rect 118240 543516 118292 543522
rect 118240 543458 118292 543464
rect 116860 543108 116912 543114
rect 116860 543050 116912 543056
rect 116872 539963 116900 543050
rect 117596 543040 117648 543046
rect 117596 542982 117648 542988
rect 117608 539963 117636 542982
rect 118252 539963 118280 543458
rect 118712 543402 118740 558282
rect 119356 543590 119384 558690
rect 120828 552770 120856 598295
rect 120920 560046 120948 625398
rect 121644 625388 121696 625394
rect 121644 625330 121696 625336
rect 121552 622396 121604 622402
rect 121552 622338 121604 622344
rect 120998 576872 121054 576881
rect 120998 576807 121054 576816
rect 120908 560040 120960 560046
rect 120908 559982 120960 559988
rect 120816 552764 120868 552770
rect 120816 552706 120868 552712
rect 121012 550186 121040 576807
rect 121458 571024 121514 571033
rect 121458 570959 121514 570968
rect 121090 564904 121146 564913
rect 121090 564839 121146 564848
rect 121000 550180 121052 550186
rect 121000 550122 121052 550128
rect 120264 549908 120316 549914
rect 120264 549850 120316 549856
rect 120276 543946 120304 549850
rect 121104 544066 121132 564839
rect 121182 562184 121238 562193
rect 121182 562119 121238 562128
rect 121196 554062 121224 562119
rect 121472 556986 121500 570959
rect 121564 559842 121592 622338
rect 121552 559836 121604 559842
rect 121552 559778 121604 559784
rect 121460 556980 121512 556986
rect 121460 556922 121512 556928
rect 121184 554056 121236 554062
rect 121184 553998 121236 554004
rect 121460 552832 121512 552838
rect 121460 552774 121512 552780
rect 121092 544060 121144 544066
rect 121092 544002 121144 544008
rect 121472 543946 121500 552774
rect 121552 551472 121604 551478
rect 121552 551414 121604 551420
rect 121564 544066 121592 551414
rect 121656 547874 121684 625330
rect 121734 613864 121790 613873
rect 121734 613799 121790 613808
rect 121748 559774 121776 613799
rect 121826 611144 121882 611153
rect 121826 611079 121882 611088
rect 121736 559768 121788 559774
rect 121736 559710 121788 559716
rect 121840 559706 121868 611079
rect 121918 601624 121974 601633
rect 121918 601559 121974 601568
rect 121828 559700 121880 559706
rect 121828 559642 121880 559648
rect 121932 549982 121960 601559
rect 122194 586664 122250 586673
rect 122194 586599 122250 586608
rect 122102 583264 122158 583273
rect 122102 583199 122158 583208
rect 122010 580544 122066 580553
rect 122010 580479 122066 580488
rect 121920 549976 121972 549982
rect 121920 549918 121972 549924
rect 121656 547846 121960 547874
rect 121552 544060 121604 544066
rect 121552 544002 121604 544008
rect 120276 543918 121132 543946
rect 121472 543918 121868 543946
rect 119344 543584 119396 543590
rect 119344 543526 119396 543532
rect 120448 543584 120500 543590
rect 120448 543526 120500 543532
rect 118712 543374 119752 543402
rect 118976 543040 119028 543046
rect 118976 542982 119028 542988
rect 118988 539963 119016 542982
rect 119724 539963 119752 543374
rect 120460 539963 120488 543526
rect 121104 539963 121132 543918
rect 121840 539963 121868 543918
rect 121932 543182 121960 547846
rect 122024 547330 122052 580479
rect 122116 551546 122144 583199
rect 122208 555558 122236 586599
rect 122196 555552 122248 555558
rect 122196 555494 122248 555500
rect 122104 551540 122156 551546
rect 122104 551482 122156 551488
rect 122012 547324 122064 547330
rect 122012 547266 122064 547272
rect 122300 543386 122328 625534
rect 122852 559978 122880 625602
rect 124220 625320 124272 625326
rect 124220 625262 124272 625268
rect 123022 619984 123078 619993
rect 123022 619919 123078 619928
rect 122930 568304 122986 568313
rect 122930 568239 122986 568248
rect 122840 559972 122892 559978
rect 122840 559914 122892 559920
rect 122840 557048 122892 557054
rect 122840 556990 122892 556996
rect 122656 547188 122708 547194
rect 122656 547130 122708 547136
rect 122564 544060 122616 544066
rect 122564 544002 122616 544008
rect 122288 543380 122340 543386
rect 122288 543322 122340 543328
rect 121920 543176 121972 543182
rect 121920 543118 121972 543124
rect 122576 539963 122604 544002
rect 122668 543590 122696 547130
rect 122852 543946 122880 556990
rect 122944 556918 122972 568239
rect 123036 559638 123064 619919
rect 123114 617264 123170 617273
rect 123114 617199 123170 617208
rect 123024 559632 123076 559638
rect 123024 559574 123076 559580
rect 123128 558414 123156 617199
rect 123574 607744 123630 607753
rect 123574 607679 123630 607688
rect 123206 605024 123262 605033
rect 123206 604959 123262 604968
rect 123116 558408 123168 558414
rect 123116 558350 123168 558356
rect 122932 556912 122984 556918
rect 122932 556854 122984 556860
rect 123220 551342 123248 604959
rect 123390 595504 123446 595513
rect 123390 595439 123446 595448
rect 123298 592784 123354 592793
rect 123298 592719 123354 592728
rect 123208 551336 123260 551342
rect 123208 551278 123260 551284
rect 123312 544474 123340 592719
rect 123404 552906 123432 595439
rect 123482 574424 123538 574433
rect 123482 574359 123538 574368
rect 123496 555626 123524 574359
rect 123484 555620 123536 555626
rect 123484 555562 123536 555568
rect 123392 552900 123444 552906
rect 123392 552842 123444 552848
rect 123588 545766 123616 607679
rect 124126 589384 124182 589393
rect 124126 589319 124128 589328
rect 124180 589319 124182 589328
rect 124128 589290 124180 589296
rect 124036 547324 124088 547330
rect 124036 547266 124088 547272
rect 123576 545760 123628 545766
rect 123576 545702 123628 545708
rect 123300 544468 123352 544474
rect 123300 544410 123352 544416
rect 122852 543918 123340 543946
rect 122656 543584 122708 543590
rect 122656 543526 122708 543532
rect 123312 539963 123340 543918
rect 124048 539963 124076 547266
rect 124232 543930 124260 625262
rect 124324 559910 124352 625670
rect 135168 625660 135220 625666
rect 135168 625602 135220 625608
rect 124404 625524 124456 625530
rect 124404 625466 124456 625472
rect 124312 559904 124364 559910
rect 124312 559846 124364 559852
rect 124312 554192 124364 554198
rect 124312 554134 124364 554140
rect 124220 543924 124272 543930
rect 124220 543866 124272 543872
rect 124324 543130 124352 554134
rect 124416 543318 124444 625466
rect 124680 625252 124732 625258
rect 124680 625194 124732 625200
rect 124588 623892 124640 623898
rect 124588 623834 124640 623840
rect 124496 623824 124548 623830
rect 124496 623766 124548 623772
rect 124508 543454 124536 623766
rect 124600 557534 124628 623834
rect 124692 560114 124720 625194
rect 133880 625184 133932 625190
rect 133880 625126 133932 625132
rect 133144 623892 133196 623898
rect 133144 623834 133196 623840
rect 126244 622804 126296 622810
rect 126244 622746 126296 622752
rect 125600 576904 125652 576910
rect 125600 576846 125652 576852
rect 124680 560108 124732 560114
rect 124680 560050 124732 560056
rect 124600 557506 124812 557534
rect 124496 543448 124548 543454
rect 124496 543390 124548 543396
rect 124404 543312 124456 543318
rect 124404 543254 124456 543260
rect 124784 543250 124812 557506
rect 125612 543930 125640 576846
rect 126152 555620 126204 555626
rect 126152 555562 126204 555568
rect 125416 543924 125468 543930
rect 125416 543866 125468 543872
rect 125600 543924 125652 543930
rect 125600 543866 125652 543872
rect 124772 543244 124824 543250
rect 124772 543186 124824 543192
rect 124324 543102 124720 543130
rect 124692 539963 124720 543102
rect 125428 539963 125456 543866
rect 126164 539963 126192 555562
rect 126256 543522 126284 622746
rect 132500 607232 132552 607238
rect 132500 607174 132552 607180
rect 131764 589348 131816 589354
rect 131764 589290 131816 589296
rect 131776 560250 131804 589290
rect 131764 560244 131816 560250
rect 131764 560186 131816 560192
rect 129740 558408 129792 558414
rect 129740 558350 129792 558356
rect 129752 557534 129780 558350
rect 129752 557506 130516 557534
rect 129004 552900 129056 552906
rect 129004 552842 129056 552848
rect 127624 545760 127676 545766
rect 127624 545702 127676 545708
rect 126888 543924 126940 543930
rect 126888 543866 126940 543872
rect 126244 543516 126296 543522
rect 126244 543458 126296 543464
rect 126900 539963 126928 543866
rect 127636 539963 127664 545702
rect 128268 543312 128320 543318
rect 128268 543254 128320 543260
rect 128280 539963 128308 543254
rect 129016 539963 129044 552842
rect 129740 544468 129792 544474
rect 129740 544410 129792 544416
rect 129752 539963 129780 544410
rect 130488 539963 130516 557506
rect 131212 549976 131264 549982
rect 131212 549918 131264 549924
rect 131224 539963 131252 549918
rect 132512 543946 132540 607174
rect 132592 558204 132644 558210
rect 132592 558146 132644 558152
rect 132604 557534 132632 558146
rect 132604 557506 132816 557534
rect 132512 543918 132632 543946
rect 131856 543584 131908 543590
rect 131856 543526 131908 543532
rect 131868 539963 131896 543526
rect 132604 539963 132632 543918
rect 132788 543402 132816 557506
rect 133156 543590 133184 623834
rect 133892 543946 133920 625126
rect 135076 622668 135128 622674
rect 135076 622610 135128 622616
rect 134892 622600 134944 622606
rect 134892 622542 134944 622548
rect 134524 594856 134576 594862
rect 134524 594798 134576 594804
rect 134536 561202 134564 594798
rect 134616 589348 134668 589354
rect 134616 589290 134668 589296
rect 134524 561196 134576 561202
rect 134524 561138 134576 561144
rect 133972 558272 134024 558278
rect 133972 558214 134024 558220
rect 133984 544082 134012 558214
rect 134628 557534 134656 589290
rect 134628 557506 134840 557534
rect 133984 544054 134748 544082
rect 133892 543918 134104 543946
rect 133144 543584 133196 543590
rect 133144 543526 133196 543532
rect 132788 543374 133368 543402
rect 133340 539963 133368 543374
rect 134076 539963 134104 543918
rect 134720 539963 134748 544054
rect 134812 543046 134840 557506
rect 134904 543454 134932 622542
rect 134984 622532 135036 622538
rect 134984 622474 135036 622480
rect 134996 543590 135024 622474
rect 134984 543584 135036 543590
rect 134984 543526 135036 543532
rect 134892 543448 134944 543454
rect 134892 543390 134944 543396
rect 135088 543182 135116 622610
rect 135076 543176 135128 543182
rect 135076 543118 135128 543124
rect 135180 543114 135208 625602
rect 136456 625592 136508 625598
rect 136456 625534 136508 625540
rect 135260 625252 135312 625258
rect 135260 625194 135312 625200
rect 135272 557534 135300 625194
rect 136364 622736 136416 622742
rect 136364 622678 136416 622684
rect 135272 557506 136220 557534
rect 135444 543720 135496 543726
rect 135444 543662 135496 543668
rect 135168 543108 135220 543114
rect 135168 543050 135220 543056
rect 134800 543040 134852 543046
rect 134800 542982 134852 542988
rect 135456 539963 135484 543662
rect 136192 539963 136220 557506
rect 136376 543522 136404 622678
rect 136364 543516 136416 543522
rect 136364 543458 136416 543464
rect 136468 543386 136496 625534
rect 137744 625388 137796 625394
rect 137744 625330 137796 625336
rect 136640 623824 136692 623830
rect 136640 623766 136692 623772
rect 136548 622464 136600 622470
rect 136548 622406 136600 622412
rect 136560 596034 136588 622406
rect 136652 596174 136680 623766
rect 137374 620664 137430 620673
rect 137374 620599 137430 620608
rect 136730 608288 136786 608297
rect 136730 608223 136786 608232
rect 136744 607238 136772 608223
rect 136732 607232 136784 607238
rect 136732 607174 136784 607180
rect 136652 596146 136772 596174
rect 136638 596048 136694 596057
rect 136560 596006 136638 596034
rect 136560 594862 136588 596006
rect 136638 595983 136694 595992
rect 136548 594856 136600 594862
rect 136548 594798 136600 594804
rect 136744 586514 136772 596146
rect 136914 589928 136970 589937
rect 136914 589863 136970 589872
rect 136928 589354 136956 589863
rect 136916 589348 136968 589354
rect 136916 589290 136968 589296
rect 136652 586486 136772 586514
rect 136652 543930 136680 586486
rect 136730 577688 136786 577697
rect 136730 577623 136786 577632
rect 136744 576910 136772 577623
rect 136732 576904 136784 576910
rect 136732 576846 136784 576852
rect 137282 574968 137338 574977
rect 137282 574903 137338 574912
rect 137190 568848 137246 568857
rect 137190 568783 137246 568792
rect 137204 551342 137232 568783
rect 137192 551336 137244 551342
rect 137192 551278 137244 551284
rect 136916 548548 136968 548554
rect 136916 548490 136968 548496
rect 136640 543924 136692 543930
rect 136640 543866 136692 543872
rect 136456 543380 136508 543386
rect 136456 543322 136508 543328
rect 136928 539963 136956 548490
rect 137296 547194 137324 574903
rect 137284 547188 137336 547194
rect 137284 547130 137336 547136
rect 137388 543726 137416 620599
rect 137650 611688 137706 611697
rect 137650 611623 137706 611632
rect 137466 583808 137522 583817
rect 137466 583743 137522 583752
rect 137480 556986 137508 583743
rect 137558 571568 137614 571577
rect 137558 571503 137614 571512
rect 137468 556980 137520 556986
rect 137468 556922 137520 556928
rect 137572 543862 137600 571503
rect 137664 560182 137692 611623
rect 137652 560176 137704 560182
rect 137652 560118 137704 560124
rect 137756 559706 137784 625330
rect 137744 559700 137796 559706
rect 137744 559642 137796 559648
rect 137652 543924 137704 543930
rect 137652 543866 137704 543872
rect 137560 543856 137612 543862
rect 137560 543798 137612 543804
rect 137376 543720 137428 543726
rect 137376 543662 137428 543668
rect 137664 539963 137692 543866
rect 137848 543658 137876 625670
rect 137940 599593 137968 683130
rect 169772 641034 169800 702406
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 169760 641028 169812 641034
rect 169760 640970 169812 640976
rect 299492 636886 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 305644 700392 305696 700398
rect 305644 700334 305696 700340
rect 299480 636880 299532 636886
rect 299480 636822 299532 636828
rect 291200 634840 291252 634846
rect 291200 634782 291252 634788
rect 280988 633684 281040 633690
rect 280988 633626 281040 633632
rect 218704 630692 218756 630698
rect 218704 630634 218756 630640
rect 217784 629944 217836 629950
rect 217784 629886 217836 629892
rect 214012 625796 214064 625802
rect 214012 625738 214064 625744
rect 186504 625728 186556 625734
rect 186504 625670 186556 625676
rect 206468 625728 206520 625734
rect 206468 625670 206520 625676
rect 160284 625660 160336 625666
rect 160284 625602 160336 625608
rect 139216 625524 139268 625530
rect 139216 625466 139268 625472
rect 139124 625456 139176 625462
rect 139124 625398 139176 625404
rect 139030 617808 139086 617817
rect 139030 617743 139086 617752
rect 138570 614408 138626 614417
rect 138570 614343 138626 614352
rect 137926 599584 137982 599593
rect 137926 599519 137982 599528
rect 137926 593464 137982 593473
rect 137926 593399 137982 593408
rect 137940 544542 137968 593399
rect 138478 562728 138534 562737
rect 138478 562663 138534 562672
rect 138492 556918 138520 562663
rect 138480 556912 138532 556918
rect 138480 556854 138532 556860
rect 138296 545964 138348 545970
rect 138296 545906 138348 545912
rect 137928 544536 137980 544542
rect 137928 544478 137980 544484
rect 137836 543652 137888 543658
rect 137836 543594 137888 543600
rect 138308 539963 138336 545906
rect 138584 543250 138612 614343
rect 138938 605568 138994 605577
rect 138938 605503 138994 605512
rect 138846 602168 138902 602177
rect 138846 602103 138902 602112
rect 138754 587208 138810 587217
rect 138754 587143 138810 587152
rect 138662 581088 138718 581097
rect 138662 581023 138718 581032
rect 138676 555558 138704 581023
rect 138664 555552 138716 555558
rect 138664 555494 138716 555500
rect 138768 548622 138796 587143
rect 138860 554062 138888 602103
rect 138848 554056 138900 554062
rect 138848 553998 138900 554004
rect 138952 552702 138980 605503
rect 139044 559842 139072 617743
rect 139032 559836 139084 559842
rect 139032 559778 139084 559784
rect 139136 559094 139164 625398
rect 139228 559638 139256 625466
rect 139860 625184 139912 625190
rect 139860 625126 139912 625132
rect 157524 625184 157576 625190
rect 157524 625126 157576 625132
rect 139306 565448 139362 565457
rect 139306 565383 139362 565392
rect 139320 559774 139348 565383
rect 139308 559768 139360 559774
rect 139308 559710 139360 559716
rect 139216 559632 139268 559638
rect 139216 559574 139268 559580
rect 139124 559088 139176 559094
rect 139124 559030 139176 559036
rect 138940 552696 138992 552702
rect 138940 552638 138992 552644
rect 138756 548616 138808 548622
rect 138756 548558 138808 548564
rect 139872 546514 139900 625126
rect 140136 625116 140188 625122
rect 140136 625058 140188 625064
rect 140148 623098 140176 625058
rect 151268 623892 151320 623898
rect 151268 623834 151320 623840
rect 140070 623070 140176 623098
rect 151280 623098 151308 623834
rect 157536 623098 157564 625126
rect 151280 623070 151662 623098
rect 157458 623070 157564 623098
rect 160296 623098 160324 625602
rect 162860 625592 162912 625598
rect 162860 625534 162912 625540
rect 162872 623098 162900 625534
rect 166172 625524 166224 625530
rect 166172 625466 166224 625472
rect 166184 623098 166212 625466
rect 174452 625456 174504 625462
rect 174452 625398 174504 625404
rect 171876 625320 171928 625326
rect 171876 625262 171928 625268
rect 168748 623824 168800 623830
rect 168748 623766 168800 623772
rect 168760 623098 168788 623766
rect 171888 623098 171916 625262
rect 174464 623098 174492 625398
rect 180340 625388 180392 625394
rect 180340 625330 180392 625336
rect 180352 623098 180380 625330
rect 183652 625252 183704 625258
rect 183652 625194 183704 625200
rect 183664 623098 183692 625194
rect 160296 623070 160678 623098
rect 162872 623070 163254 623098
rect 166184 623070 166474 623098
rect 168760 623070 169050 623098
rect 171888 623070 172270 623098
rect 174464 623070 174846 623098
rect 180352 623070 180642 623098
rect 183664 623070 183862 623098
rect 186516 622962 186544 625670
rect 190000 625388 190052 625394
rect 190000 625330 190052 625336
rect 204536 625388 204588 625394
rect 204536 625330 204588 625336
rect 190012 623098 190040 625330
rect 192576 625252 192628 625258
rect 192576 625194 192628 625200
rect 204444 625252 204496 625258
rect 204444 625194 204496 625200
rect 192588 623098 192616 625194
rect 195704 625184 195756 625190
rect 195704 625126 195756 625132
rect 201684 625184 201736 625190
rect 201684 625126 201736 625132
rect 195716 623098 195744 625126
rect 189658 623070 190040 623098
rect 192234 623070 192616 623098
rect 195454 623070 195744 623098
rect 186438 622934 186544 622962
rect 177868 622810 178066 622826
rect 177856 622804 178066 622810
rect 177908 622798 178066 622804
rect 177856 622746 177908 622752
rect 145564 622736 145616 622742
rect 145616 622684 145866 622690
rect 145564 622678 145866 622684
rect 145576 622662 145866 622678
rect 149086 622674 149192 622690
rect 149086 622668 149204 622674
rect 149086 622662 149152 622668
rect 149152 622610 149204 622616
rect 154580 622600 154632 622606
rect 143000 622538 143290 622554
rect 154632 622548 154882 622554
rect 154580 622542 154882 622548
rect 142988 622532 143290 622538
rect 143040 622526 143290 622532
rect 154592 622526 154882 622542
rect 142988 622474 143040 622480
rect 198030 622402 198320 622418
rect 198030 622396 198332 622402
rect 198030 622390 198280 622396
rect 200606 622390 200712 622418
rect 198280 622338 198332 622344
rect 159836 560238 160034 560266
rect 194612 560238 194810 560266
rect 140780 560176 140832 560182
rect 140070 560102 140360 560130
rect 140780 560118 140832 560124
rect 140332 558482 140360 560102
rect 140320 558476 140372 558482
rect 140320 558418 140372 558424
rect 140792 557534 140820 560118
rect 142646 560102 142936 560130
rect 142160 559088 142212 559094
rect 142160 559030 142212 559036
rect 140792 557506 141280 557534
rect 140504 547392 140556 547398
rect 140504 547334 140556 547340
rect 139860 546508 139912 546514
rect 139860 546450 139912 546456
rect 139032 545896 139084 545902
rect 139032 545838 139084 545844
rect 138572 543244 138624 543250
rect 138572 543186 138624 543192
rect 139044 539963 139072 545838
rect 139768 543856 139820 543862
rect 139768 543798 139820 543804
rect 139780 539963 139808 543798
rect 140516 539963 140544 547334
rect 141252 539963 141280 557506
rect 141884 546508 141936 546514
rect 141884 546450 141936 546456
rect 141896 539963 141924 546450
rect 142172 543930 142200 559030
rect 142908 558550 142936 560102
rect 144932 560102 145222 560130
rect 147784 560102 148442 560130
rect 151018 560102 151400 560130
rect 142896 558544 142948 558550
rect 142896 558486 142948 558492
rect 144932 558346 144960 560102
rect 147680 558680 147732 558686
rect 147680 558622 147732 558628
rect 144920 558340 144972 558346
rect 144920 558282 144972 558288
rect 143540 555688 143592 555694
rect 143540 555630 143592 555636
rect 142620 550044 142672 550050
rect 142620 549986 142672 549992
rect 142160 543924 142212 543930
rect 142160 543866 142212 543872
rect 142632 539963 142660 549986
rect 143552 543946 143580 555630
rect 144736 551404 144788 551410
rect 144736 551346 144788 551352
rect 143356 543924 143408 543930
rect 143552 543918 144132 543946
rect 143356 543866 143408 543872
rect 143368 539963 143396 543866
rect 144104 539963 144132 543918
rect 144748 539963 144776 551346
rect 147692 543930 147720 558622
rect 147784 544406 147812 560102
rect 150624 559836 150676 559842
rect 150624 559778 150676 559784
rect 149060 556980 149112 556986
rect 149060 556922 149112 556928
rect 147864 547188 147916 547194
rect 147864 547130 147916 547136
rect 147772 544400 147824 544406
rect 147772 544342 147824 544348
rect 147680 543924 147732 543930
rect 147680 543866 147732 543872
rect 145472 543652 145524 543658
rect 145472 543594 145524 543600
rect 145484 539963 145512 543594
rect 146944 543584 146996 543590
rect 146944 543526 146996 543532
rect 146208 543040 146260 543046
rect 146208 542982 146260 542988
rect 146220 539963 146248 542982
rect 146956 539963 146984 543526
rect 147876 540138 147904 547130
rect 148324 543924 148376 543930
rect 148324 543866 148376 543872
rect 147708 540110 147904 540138
rect 147708 539920 147736 540110
rect 148336 539963 148364 543866
rect 149072 539963 149100 556922
rect 149796 544536 149848 544542
rect 149796 544478 149848 544484
rect 149808 539963 149836 544478
rect 150636 540138 150664 559778
rect 151372 558618 151400 560102
rect 153856 560102 154238 560130
rect 156432 560102 156814 560130
rect 151820 559700 151872 559706
rect 151820 559642 151872 559648
rect 151360 558612 151412 558618
rect 151360 558554 151412 558560
rect 151832 557534 151860 559642
rect 153856 558414 153884 560102
rect 156144 559836 156196 559842
rect 156144 559778 156196 559784
rect 154580 559700 154632 559706
rect 154580 559642 154632 559648
rect 153844 558408 153896 558414
rect 153844 558350 153896 558356
rect 151832 557506 151952 557534
rect 151268 543108 151320 543114
rect 151268 543050 151320 543056
rect 150560 540110 150664 540138
rect 150560 539920 150588 540110
rect 151280 539963 151308 543050
rect 151924 539963 151952 557506
rect 153384 548616 153436 548622
rect 153384 548558 153436 548564
rect 152648 544536 152700 544542
rect 152648 544478 152700 544484
rect 152660 539963 152688 544478
rect 153396 539963 153424 548558
rect 154592 543930 154620 559642
rect 154672 558408 154724 558414
rect 154672 558350 154724 558356
rect 154684 557534 154712 558350
rect 156156 557534 156184 559778
rect 154684 557506 154896 557534
rect 156156 557506 156276 557534
rect 154580 543924 154632 543930
rect 154580 543866 154632 543872
rect 154120 543108 154172 543114
rect 154120 543050 154172 543056
rect 154132 539963 154160 543050
rect 154868 539963 154896 557506
rect 155500 543924 155552 543930
rect 155500 543866 155552 543872
rect 155512 539963 155540 543866
rect 156248 539963 156276 557506
rect 156432 551410 156460 560102
rect 157984 559904 158036 559910
rect 157984 559846 158036 559852
rect 156420 551404 156472 551410
rect 156420 551346 156472 551352
rect 157892 548616 157944 548622
rect 157892 548558 157944 548564
rect 156972 543516 157024 543522
rect 156972 543458 157024 543464
rect 156984 539963 157012 543458
rect 157708 543448 157760 543454
rect 157708 543390 157760 543396
rect 157720 539963 157748 543390
rect 157904 543130 157932 548558
rect 157996 543318 158024 559846
rect 159364 558476 159416 558482
rect 159364 558418 159416 558424
rect 158720 558340 158772 558346
rect 158720 558282 158772 558288
rect 158732 543930 158760 558282
rect 159088 556912 159140 556918
rect 159088 556854 159140 556860
rect 158720 543924 158772 543930
rect 158720 543866 158772 543872
rect 157984 543312 158036 543318
rect 157984 543254 158036 543260
rect 157904 543102 158392 543130
rect 158364 539963 158392 543102
rect 159100 539963 159128 556854
rect 159376 543726 159404 558418
rect 159836 556918 159864 560238
rect 162320 560102 162610 560130
rect 165632 560102 165830 560130
rect 168406 560102 168512 560130
rect 160100 559768 160152 559774
rect 160100 559710 160152 559716
rect 159824 556912 159876 556918
rect 159824 556854 159876 556860
rect 160112 543930 160140 559710
rect 161664 559632 161716 559638
rect 161664 559574 161716 559580
rect 161572 558816 161624 558822
rect 161572 558758 161624 558764
rect 160744 558544 160796 558550
rect 160744 558486 160796 558492
rect 160560 554056 160612 554062
rect 160560 553998 160612 554004
rect 159824 543924 159876 543930
rect 159824 543866 159876 543872
rect 160100 543924 160152 543930
rect 160100 543866 160152 543872
rect 159364 543720 159416 543726
rect 159364 543662 159416 543668
rect 159836 539963 159864 543866
rect 160572 539963 160600 553998
rect 160756 543318 160784 558486
rect 161584 543930 161612 558758
rect 161676 557534 161704 559574
rect 162320 558686 162348 560102
rect 164332 559972 164384 559978
rect 164332 559914 164384 559920
rect 162308 558680 162360 558686
rect 162308 558622 162360 558628
rect 161676 557506 161980 557534
rect 161296 543924 161348 543930
rect 161296 543866 161348 543872
rect 161572 543924 161624 543930
rect 161572 543866 161624 543872
rect 160744 543312 160796 543318
rect 160744 543254 160796 543260
rect 161308 539963 161336 543866
rect 161952 539963 161980 557506
rect 164344 543930 164372 559914
rect 164884 558612 164936 558618
rect 164884 558554 164936 558560
rect 162676 543924 162728 543930
rect 162676 543866 162728 543872
rect 164332 543924 164384 543930
rect 164332 543866 164384 543872
rect 162688 539963 162716 543866
rect 163412 543720 163464 543726
rect 163412 543662 163464 543668
rect 163424 539963 163452 543662
rect 164896 543658 164924 558554
rect 165528 543924 165580 543930
rect 165528 543866 165580 543872
rect 164884 543652 164936 543658
rect 164884 543594 164936 543600
rect 164148 543448 164200 543454
rect 164148 543390 164200 543396
rect 164160 539963 164188 543390
rect 164884 543380 164936 543386
rect 164884 543322 164936 543328
rect 164896 539963 164924 543322
rect 165540 539963 165568 543866
rect 165632 543726 165660 560102
rect 168484 558822 168512 560102
rect 171336 560102 171626 560130
rect 174004 560102 174202 560130
rect 177040 560102 177422 560130
rect 179616 560102 179998 560130
rect 182928 560102 183218 560130
rect 185504 560102 185794 560130
rect 188632 560102 189014 560130
rect 190564 560102 191590 560130
rect 168472 558816 168524 558822
rect 168472 558758 168524 558764
rect 171336 558414 171364 560102
rect 173900 558816 173952 558822
rect 173900 558758 173952 558764
rect 171324 558408 171376 558414
rect 171324 558350 171376 558356
rect 173440 556912 173492 556918
rect 173440 556854 173492 556860
rect 171324 554260 171376 554266
rect 171324 554202 171376 554208
rect 166264 552696 166316 552702
rect 166264 552638 166316 552644
rect 165620 543720 165672 543726
rect 165620 543662 165672 543668
rect 166276 539963 166304 552638
rect 169116 551336 169168 551342
rect 169116 551278 169168 551284
rect 168380 544604 168432 544610
rect 168380 544546 168432 544552
rect 167000 544400 167052 544406
rect 167000 544342 167052 544348
rect 167012 539963 167040 544342
rect 167736 543312 167788 543318
rect 167736 543254 167788 543260
rect 167748 539963 167776 543254
rect 168392 539963 168420 544546
rect 169128 539963 169156 551278
rect 169852 543720 169904 543726
rect 169852 543662 169904 543668
rect 169864 539963 169892 543662
rect 170588 543312 170640 543318
rect 170588 543254 170640 543260
rect 170600 539963 170628 543254
rect 171336 539963 171364 554202
rect 172704 543652 172756 543658
rect 172704 543594 172756 543600
rect 171968 543176 172020 543182
rect 171968 543118 172020 543124
rect 171980 539963 172008 543118
rect 172716 539963 172744 543594
rect 173452 539963 173480 556854
rect 173912 543266 173940 558758
rect 174004 543454 174032 560102
rect 177040 558210 177068 560102
rect 179616 558822 179644 560102
rect 182364 560040 182416 560046
rect 182364 559982 182416 559988
rect 182272 559768 182324 559774
rect 182272 559710 182324 559716
rect 179696 559632 179748 559638
rect 179696 559574 179748 559580
rect 179604 558816 179656 558822
rect 179604 558758 179656 558764
rect 177028 558204 177080 558210
rect 177028 558146 177080 558152
rect 177304 558204 177356 558210
rect 177304 558146 177356 558152
rect 174912 555552 174964 555558
rect 174912 555494 174964 555500
rect 173992 543448 174044 543454
rect 173992 543390 174044 543396
rect 173912 543238 174216 543266
rect 174188 539963 174216 543238
rect 174924 539963 174952 555494
rect 176660 551540 176712 551546
rect 176660 551482 176712 551488
rect 176672 543946 176700 551482
rect 177316 549982 177344 558146
rect 179708 557534 179736 559574
rect 179708 557506 179920 557534
rect 178040 557116 178092 557122
rect 178040 557058 178092 557064
rect 177764 550112 177816 550118
rect 177764 550054 177816 550060
rect 177304 549976 177356 549982
rect 177304 549918 177356 549924
rect 176672 543918 177068 543946
rect 175556 543244 175608 543250
rect 175556 543186 175608 543192
rect 175568 539963 175596 543186
rect 176292 543176 176344 543182
rect 176292 543118 176344 543124
rect 176304 539963 176332 543118
rect 177040 539963 177068 543918
rect 177776 539963 177804 550054
rect 178052 543946 178080 557058
rect 179512 556912 179564 556918
rect 179512 556854 179564 556860
rect 179144 552696 179196 552702
rect 179144 552638 179196 552644
rect 178052 543918 178540 543946
rect 178512 539963 178540 543918
rect 179156 539963 179184 552638
rect 179524 543998 179552 556854
rect 179512 543992 179564 543998
rect 179512 543934 179564 543940
rect 179892 539963 179920 557506
rect 181352 555552 181404 555558
rect 181352 555494 181404 555500
rect 180616 543992 180668 543998
rect 180616 543934 180668 543940
rect 180628 539963 180656 543934
rect 181364 539963 181392 555494
rect 182284 543946 182312 559710
rect 182376 557534 182404 559982
rect 182928 558346 182956 560102
rect 182916 558340 182968 558346
rect 182916 558282 182968 558288
rect 185504 557938 185532 560102
rect 188344 558476 188396 558482
rect 188344 558418 188396 558424
rect 187884 558408 187936 558414
rect 187884 558350 187936 558356
rect 184204 557932 184256 557938
rect 184204 557874 184256 557880
rect 185492 557932 185544 557938
rect 185492 557874 185544 557880
rect 182376 557506 183508 557534
rect 182284 543918 182772 543946
rect 181996 543244 182048 543250
rect 181996 543186 182048 543192
rect 182008 539963 182036 543186
rect 182744 539963 182772 543918
rect 183480 539963 183508 557506
rect 184216 547194 184244 557874
rect 186320 554056 186372 554062
rect 186320 553998 186372 554004
rect 185584 547256 185636 547262
rect 185584 547198 185636 547204
rect 184204 547188 184256 547194
rect 184204 547130 184256 547136
rect 184940 546032 184992 546038
rect 184940 545974 184992 545980
rect 184204 544400 184256 544406
rect 184204 544342 184256 544348
rect 184216 539963 184244 544342
rect 184952 539963 184980 545974
rect 185596 539963 185624 547198
rect 186332 543930 186360 553998
rect 186412 551336 186464 551342
rect 186412 551278 186464 551284
rect 186320 543924 186372 543930
rect 186320 543866 186372 543872
rect 186424 540138 186452 551278
rect 187792 547188 187844 547194
rect 187792 547130 187844 547136
rect 187056 543924 187108 543930
rect 187056 543866 187108 543872
rect 186348 540110 186452 540138
rect 186348 539920 186376 540110
rect 187068 539963 187096 543866
rect 187804 539963 187832 547130
rect 187896 543946 187924 558350
rect 188356 547398 188384 558418
rect 188632 558210 188660 560102
rect 190460 558340 190512 558346
rect 190460 558282 190512 558288
rect 188620 558204 188672 558210
rect 188620 558146 188672 558152
rect 189080 549976 189132 549982
rect 189080 549918 189132 549924
rect 188344 547392 188396 547398
rect 188344 547334 188396 547340
rect 189092 543946 189120 549918
rect 189908 548684 189960 548690
rect 189908 548626 189960 548632
rect 187896 543918 188568 543946
rect 189092 543918 189212 543946
rect 188540 539963 188568 543918
rect 189184 539963 189212 543918
rect 189920 539963 189948 548626
rect 190472 547874 190500 558282
rect 190564 549914 190592 560102
rect 191840 558204 191892 558210
rect 191840 558146 191892 558152
rect 190552 549908 190604 549914
rect 190552 549850 190604 549856
rect 190472 547846 191420 547874
rect 190644 547392 190696 547398
rect 190644 547334 190696 547340
rect 190656 539963 190684 547334
rect 191392 539963 191420 547846
rect 191852 543930 191880 558146
rect 194612 557534 194640 560238
rect 197386 560102 197492 560130
rect 197464 558278 197492 560102
rect 200224 560102 200606 560130
rect 199384 558544 199436 558550
rect 199384 558486 199436 558492
rect 197452 558272 197504 558278
rect 197452 558214 197504 558220
rect 194612 557506 194732 557534
rect 194600 556980 194652 556986
rect 194600 556922 194652 556928
rect 193220 555756 193272 555762
rect 193220 555698 193272 555704
rect 192116 551608 192168 551614
rect 192116 551550 192168 551556
rect 191840 543924 191892 543930
rect 191840 543866 191892 543872
rect 192128 539963 192156 551550
rect 193232 543930 193260 555698
rect 193496 550180 193548 550186
rect 193496 550122 193548 550128
rect 192760 543924 192812 543930
rect 192760 543866 192812 543872
rect 193220 543924 193272 543930
rect 193220 543866 193272 543872
rect 192772 539963 192800 543866
rect 193508 539963 193536 550122
rect 194612 543946 194640 556922
rect 194704 545766 194732 557506
rect 198004 554124 198056 554130
rect 198004 554066 198056 554072
rect 195980 552764 196032 552770
rect 195980 552706 196032 552712
rect 194692 545760 194744 545766
rect 194692 545702 194744 545708
rect 195992 543946 196020 552706
rect 197084 549908 197136 549914
rect 197084 549850 197136 549856
rect 194232 543924 194284 543930
rect 194612 543918 195008 543946
rect 195992 543918 196388 543946
rect 194232 543866 194284 543872
rect 194244 539963 194272 543866
rect 194980 539963 195008 543918
rect 195612 543380 195664 543386
rect 195612 543322 195664 543328
rect 195624 539963 195652 543322
rect 196360 539963 196388 543918
rect 197096 539963 197124 549850
rect 197820 545760 197872 545766
rect 197820 545702 197872 545708
rect 197832 539963 197860 545702
rect 198016 543250 198044 554066
rect 199200 548752 199252 548758
rect 199200 548694 199252 548700
rect 198556 545828 198608 545834
rect 198556 545770 198608 545776
rect 198004 543244 198056 543250
rect 198004 543186 198056 543192
rect 198568 539963 198596 545770
rect 199212 539963 199240 548694
rect 199396 543318 199424 558486
rect 200224 558482 200252 560102
rect 200212 558476 200264 558482
rect 200212 558418 200264 558424
rect 199476 558272 199528 558278
rect 199476 558214 199528 558220
rect 199384 543312 199436 543318
rect 199384 543254 199436 543260
rect 199488 543114 199516 558214
rect 200212 551404 200264 551410
rect 200212 551346 200264 551352
rect 200224 543946 200252 551346
rect 200684 544610 200712 622390
rect 201500 622396 201552 622402
rect 201500 622338 201552 622344
rect 200762 610600 200818 610609
rect 200762 610535 200818 610544
rect 200776 555626 200804 610535
rect 200854 598360 200910 598369
rect 200854 598295 200910 598304
rect 200764 555620 200816 555626
rect 200764 555562 200816 555568
rect 200868 545970 200896 598295
rect 200946 574152 201002 574161
rect 200946 574087 201002 574096
rect 200960 548622 200988 574087
rect 201038 568304 201094 568313
rect 201038 568239 201094 568248
rect 201052 552838 201080 568239
rect 201130 562184 201186 562193
rect 201130 562119 201186 562128
rect 201144 554198 201172 562119
rect 201132 554192 201184 554198
rect 201132 554134 201184 554140
rect 201040 552832 201092 552838
rect 201040 552774 201092 552780
rect 200948 548616 201000 548622
rect 200948 548558 201000 548564
rect 200856 545964 200908 545970
rect 200856 545906 200908 545912
rect 200672 544604 200724 544610
rect 200672 544546 200724 544552
rect 200224 543918 200712 543946
rect 199936 543448 199988 543454
rect 199936 543390 199988 543396
rect 199476 543108 199528 543114
rect 199476 543050 199528 543056
rect 199948 539963 199976 543390
rect 200684 539963 200712 543918
rect 201408 543720 201460 543726
rect 201408 543662 201460 543668
rect 201420 539963 201448 543662
rect 201512 543046 201540 622338
rect 201590 619984 201646 619993
rect 201590 619919 201646 619928
rect 201604 551478 201632 619919
rect 201696 559978 201724 625126
rect 204260 623824 204312 623830
rect 204260 623766 204312 623772
rect 202970 617264 203026 617273
rect 202970 617199 203026 617208
rect 201866 613864 201922 613873
rect 201866 613799 201922 613808
rect 201774 605024 201830 605033
rect 201774 604959 201830 604968
rect 201684 559972 201736 559978
rect 201684 559914 201736 559920
rect 201592 551472 201644 551478
rect 201592 551414 201644 551420
rect 201788 547330 201816 604959
rect 201880 555694 201908 613799
rect 202878 607744 202934 607753
rect 202878 607679 202934 607688
rect 201958 592784 202014 592793
rect 201958 592719 202014 592728
rect 201868 555688 201920 555694
rect 201868 555630 201920 555636
rect 201776 547324 201828 547330
rect 201776 547266 201828 547272
rect 201972 544542 202000 592719
rect 202234 586664 202290 586673
rect 202234 586599 202290 586608
rect 202050 583264 202106 583273
rect 202050 583199 202106 583208
rect 202064 545902 202092 583199
rect 202142 580544 202198 580553
rect 202142 580479 202198 580488
rect 202156 550050 202184 580479
rect 202248 557054 202276 586599
rect 202326 571024 202382 571033
rect 202326 570959 202382 570968
rect 202236 557048 202288 557054
rect 202236 556990 202288 556996
rect 202144 550044 202196 550050
rect 202144 549986 202196 549992
rect 202340 548554 202368 570959
rect 202328 548548 202380 548554
rect 202328 548490 202380 548496
rect 202052 545896 202104 545902
rect 202052 545838 202104 545844
rect 201960 544536 202012 544542
rect 201960 544478 202012 544484
rect 202892 544474 202920 607679
rect 202984 558550 203012 617199
rect 203062 601624 203118 601633
rect 203062 601559 203118 601568
rect 202972 558544 203024 558550
rect 202972 558486 203024 558492
rect 203076 552906 203104 601559
rect 203154 595504 203210 595513
rect 203154 595439 203210 595448
rect 203168 558278 203196 595439
rect 204166 589384 204222 589393
rect 204166 589319 204168 589328
rect 204220 589319 204222 589328
rect 204168 589290 204220 589296
rect 203246 577144 203302 577153
rect 203246 577079 203302 577088
rect 203260 559910 203288 577079
rect 203338 564904 203394 564913
rect 203338 564839 203394 564848
rect 203248 559904 203300 559910
rect 203248 559846 203300 559852
rect 203156 558272 203208 558278
rect 203156 558214 203208 558220
rect 203352 554266 203380 564839
rect 203340 554260 203392 554266
rect 203340 554202 203392 554208
rect 203064 552900 203116 552906
rect 203064 552842 203116 552848
rect 202880 544468 202932 544474
rect 202880 544410 202932 544416
rect 202144 543244 202196 543250
rect 202144 543186 202196 543192
rect 201500 543040 201552 543046
rect 201500 542982 201552 542988
rect 202156 539963 202184 543186
rect 203524 543108 203576 543114
rect 203524 543050 203576 543056
rect 202788 543040 202840 543046
rect 202788 542982 202840 542988
rect 202800 539963 202828 542982
rect 203536 539963 203564 543050
rect 204272 539963 204300 623766
rect 204352 622736 204404 622742
rect 204352 622678 204404 622684
rect 204364 543946 204392 622678
rect 204456 559706 204484 625194
rect 204548 559842 204576 625330
rect 206284 623892 206336 623898
rect 206284 623834 206336 623840
rect 204904 607232 204956 607238
rect 204904 607174 204956 607180
rect 204536 559836 204588 559842
rect 204536 559778 204588 559784
rect 204444 559700 204496 559706
rect 204444 559642 204496 559648
rect 204916 547398 204944 607174
rect 205640 548616 205692 548622
rect 205640 548558 205692 548564
rect 204904 547392 204956 547398
rect 204904 547334 204956 547340
rect 204364 543918 205036 543946
rect 205008 539963 205036 543918
rect 205652 539963 205680 548558
rect 206296 543726 206324 623834
rect 206376 622600 206428 622606
rect 206376 622542 206428 622548
rect 206388 547874 206416 622542
rect 206480 548690 206508 625670
rect 212540 625660 212592 625666
rect 212540 625602 212592 625608
rect 209780 625388 209832 625394
rect 209780 625330 209832 625336
rect 208400 622668 208452 622674
rect 208400 622610 208452 622616
rect 207020 593428 207072 593434
rect 207020 593370 207072 593376
rect 206560 574116 206612 574122
rect 206560 574058 206612 574064
rect 206572 557122 206600 574058
rect 207032 557534 207060 593370
rect 207032 557506 207888 557534
rect 206560 557116 206612 557122
rect 206560 557058 206612 557064
rect 206468 548684 206520 548690
rect 206468 548626 206520 548632
rect 206388 547846 206508 547874
rect 206376 545964 206428 545970
rect 206376 545906 206428 545912
rect 206284 543720 206336 543726
rect 206284 543662 206336 543668
rect 206388 539963 206416 545906
rect 206480 543386 206508 547846
rect 207112 543720 207164 543726
rect 207112 543662 207164 543668
rect 206468 543380 206520 543386
rect 206468 543322 206520 543328
rect 207124 539963 207152 543662
rect 207860 539963 207888 557506
rect 208412 543930 208440 622610
rect 208492 616888 208544 616894
rect 208492 616830 208544 616836
rect 208504 557534 208532 616830
rect 209044 562352 209096 562358
rect 209044 562294 209096 562300
rect 208504 557506 208624 557534
rect 208400 543924 208452 543930
rect 208400 543866 208452 543872
rect 208596 539963 208624 557506
rect 209056 543726 209084 562294
rect 209792 543946 209820 625330
rect 210424 623960 210476 623966
rect 210424 623902 210476 623908
rect 210332 550044 210384 550050
rect 210332 549986 210384 549992
rect 209228 543924 209280 543930
rect 209792 543918 210004 543946
rect 209228 543866 209280 543872
rect 209044 543720 209096 543726
rect 209044 543662 209096 543668
rect 209240 539963 209268 543866
rect 209976 539963 210004 543918
rect 210344 543266 210372 549986
rect 210436 543454 210464 623902
rect 211804 622532 211856 622538
rect 211804 622474 211856 622480
rect 210516 589416 210568 589422
rect 210516 589358 210568 589364
rect 210528 551546 210556 589358
rect 211160 586900 211212 586906
rect 211160 586842 211212 586848
rect 210608 571396 210660 571402
rect 210608 571338 210660 571344
rect 210516 551540 210568 551546
rect 210516 551482 210568 551488
rect 210620 545766 210648 571338
rect 211068 547392 211120 547398
rect 211068 547334 211120 547340
rect 210608 545760 210660 545766
rect 210608 545702 210660 545708
rect 210424 543448 210476 543454
rect 210424 543390 210476 543396
rect 210344 543238 210740 543266
rect 210712 539963 210740 543238
rect 211080 543046 211108 547334
rect 211172 543946 211200 586842
rect 211620 551472 211672 551478
rect 211620 551414 211672 551420
rect 211172 543918 211476 543946
rect 211068 543040 211120 543046
rect 211068 542982 211120 542988
rect 211448 539963 211476 543918
rect 211632 542994 211660 551414
rect 211816 543114 211844 622474
rect 212552 543930 212580 625602
rect 213920 625320 213972 625326
rect 213920 625262 213972 625268
rect 213184 619676 213236 619682
rect 213184 619618 213236 619624
rect 212632 558476 212684 558482
rect 212632 558418 212684 558424
rect 212644 557534 212672 558418
rect 212644 557506 212856 557534
rect 212540 543924 212592 543930
rect 212540 543866 212592 543872
rect 211804 543108 211856 543114
rect 211804 543050 211856 543056
rect 211632 542966 212212 542994
rect 212184 539963 212212 542966
rect 212828 539963 212856 557506
rect 213196 550186 213224 619618
rect 213184 550180 213236 550186
rect 213184 550122 213236 550128
rect 213932 543946 213960 625262
rect 214024 557534 214052 625738
rect 215300 624096 215352 624102
rect 215300 624038 215352 624044
rect 214564 622804 214616 622810
rect 214564 622746 214616 622752
rect 214024 557506 214512 557534
rect 213552 543924 213604 543930
rect 213932 543918 214328 543946
rect 213552 543866 213604 543872
rect 213564 539963 213592 543866
rect 214300 539963 214328 543918
rect 214484 542994 214512 557506
rect 214576 543182 214604 622746
rect 215312 563054 215340 624038
rect 217324 622396 217376 622402
rect 217324 622338 217376 622344
rect 216678 620664 216734 620673
rect 216678 620599 216734 620608
rect 216692 619682 216720 620599
rect 216680 619676 216732 619682
rect 216680 619618 216732 619624
rect 216678 617808 216734 617817
rect 216678 617743 216734 617752
rect 216692 616894 216720 617743
rect 216680 616888 216732 616894
rect 216680 616830 216732 616836
rect 215942 611688 215998 611697
rect 215942 611623 215998 611632
rect 215312 563026 215800 563054
rect 214564 543176 214616 543182
rect 214564 543118 214616 543124
rect 214484 542966 215064 542994
rect 215036 539963 215064 542966
rect 215772 539963 215800 563026
rect 215956 548758 215984 611623
rect 216678 608288 216734 608297
rect 216678 608223 216734 608232
rect 216692 607238 216720 608223
rect 216680 607232 216732 607238
rect 216680 607174 216732 607180
rect 217230 602168 217286 602177
rect 217230 602103 217286 602112
rect 216678 593464 216734 593473
rect 216678 593399 216680 593408
rect 216732 593399 216734 593408
rect 216680 593370 216732 593376
rect 216678 589928 216734 589937
rect 216678 589863 216734 589872
rect 216692 589422 216720 589863
rect 216680 589416 216732 589422
rect 216680 589358 216732 589364
rect 216772 589348 216824 589354
rect 216772 589290 216824 589296
rect 216678 587208 216734 587217
rect 216678 587143 216734 587152
rect 216692 586906 216720 587143
rect 216680 586900 216732 586906
rect 216680 586842 216732 586848
rect 216034 577688 216090 577697
rect 216034 577623 216090 577632
rect 215944 548752 215996 548758
rect 215944 548694 215996 548700
rect 216048 546038 216076 577623
rect 216678 574968 216734 574977
rect 216678 574903 216734 574912
rect 216692 574122 216720 574903
rect 216680 574116 216732 574122
rect 216680 574058 216732 574064
rect 216678 571568 216734 571577
rect 216678 571503 216734 571512
rect 216692 571402 216720 571503
rect 216680 571396 216732 571402
rect 216680 571338 216732 571344
rect 216784 560250 216812 589290
rect 217138 562728 217194 562737
rect 217138 562663 217194 562672
rect 216772 560244 216824 560250
rect 216772 560186 216824 560192
rect 216128 559700 216180 559706
rect 216128 559642 216180 559648
rect 216036 546032 216088 546038
rect 216036 545974 216088 545980
rect 216140 543250 216168 559642
rect 216128 543244 216180 543250
rect 216128 543186 216180 543192
rect 216404 543176 216456 543182
rect 216404 543118 216456 543124
rect 216416 539963 216444 543118
rect 217152 539963 217180 562663
rect 217244 543726 217272 602103
rect 217336 551614 217364 622338
rect 217690 614408 217746 614417
rect 217690 614343 217746 614352
rect 217414 583808 217470 583817
rect 217414 583743 217470 583752
rect 217428 562358 217456 583743
rect 217704 581738 217732 614343
rect 217796 599593 217824 629886
rect 217876 625592 217928 625598
rect 217876 625534 217928 625540
rect 217782 599584 217838 599593
rect 217782 599519 217838 599528
rect 217692 581732 217744 581738
rect 217692 581674 217744 581680
rect 217690 581088 217746 581097
rect 217690 581023 217746 581032
rect 217598 565448 217654 565457
rect 217598 565383 217654 565392
rect 217416 562352 217468 562358
rect 217416 562294 217468 562300
rect 217324 551608 217376 551614
rect 217324 551550 217376 551556
rect 217232 543720 217284 543726
rect 217232 543662 217284 543668
rect 217612 543658 217640 565383
rect 217704 560318 217732 581023
rect 217692 560312 217744 560318
rect 217692 560254 217744 560260
rect 217888 559366 217916 625534
rect 217968 622872 218020 622878
rect 217968 622814 218020 622820
rect 217876 559360 217928 559366
rect 217876 559302 217928 559308
rect 217876 545896 217928 545902
rect 217876 545838 217928 545844
rect 217600 543652 217652 543658
rect 217600 543594 217652 543600
rect 217888 539963 217916 545838
rect 217980 543250 218008 622814
rect 218716 622470 218744 630634
rect 280712 630012 280764 630018
rect 280712 629954 280764 629960
rect 225420 625796 225472 625802
rect 225420 625738 225472 625744
rect 218888 625524 218940 625530
rect 218888 625466 218940 625472
rect 218796 625456 218848 625462
rect 218796 625398 218848 625404
rect 218704 622464 218756 622470
rect 218704 622406 218756 622412
rect 218716 596193 218744 622406
rect 218702 596184 218758 596193
rect 218702 596119 218758 596128
rect 218704 581732 218756 581738
rect 218704 581674 218756 581680
rect 218612 543720 218664 543726
rect 218612 543662 218664 543668
rect 217968 543244 218020 543250
rect 217968 543186 218020 543192
rect 218624 539963 218652 543662
rect 218716 543046 218744 581674
rect 218808 555762 218836 625398
rect 218900 560046 218928 625466
rect 219348 625252 219400 625258
rect 219348 625194 219400 625200
rect 219254 605568 219310 605577
rect 219254 605503 219310 605512
rect 219162 568848 219218 568857
rect 219162 568783 219218 568792
rect 218888 560040 218940 560046
rect 218888 559982 218940 559988
rect 218796 555756 218848 555762
rect 218796 555698 218848 555704
rect 219176 544542 219204 568783
rect 219268 557530 219296 605503
rect 219360 559094 219388 625194
rect 219624 624028 219676 624034
rect 219624 623970 219676 623976
rect 219636 615494 219664 623970
rect 225432 623098 225460 625738
rect 231308 625728 231360 625734
rect 231308 625670 231360 625676
rect 231320 623098 231348 625670
rect 271880 625660 271932 625666
rect 271880 625602 271932 625608
rect 242900 625592 242952 625598
rect 242900 625534 242952 625540
rect 234620 624096 234672 624102
rect 234620 624038 234672 624044
rect 234632 623098 234660 624038
rect 237564 623960 237616 623966
rect 237564 623902 237616 623908
rect 225432 623070 225814 623098
rect 231320 623070 231610 623098
rect 234632 623070 234830 623098
rect 237576 622962 237604 623902
rect 242912 623098 242940 625534
rect 251916 625524 251968 625530
rect 251916 625466 251968 625472
rect 246028 624028 246080 624034
rect 246028 623970 246080 623976
rect 246040 623098 246068 623970
rect 251928 623098 251956 625466
rect 263600 625456 263652 625462
rect 263600 625398 263652 625404
rect 260196 625388 260248 625394
rect 260196 625330 260248 625336
rect 254492 623892 254544 623898
rect 254492 623834 254544 623840
rect 254504 623098 254532 623834
rect 260208 623098 260236 625330
rect 263612 623098 263640 625398
rect 269212 625320 269264 625326
rect 269212 625262 269264 625268
rect 269224 623098 269252 625262
rect 271892 623098 271920 625602
rect 275100 625252 275152 625258
rect 275100 625194 275152 625200
rect 275112 623098 275140 625194
rect 277676 623824 277728 623830
rect 277676 623766 277728 623772
rect 277688 623098 277716 623766
rect 242912 623070 243202 623098
rect 246040 623070 246422 623098
rect 251928 623070 252218 623098
rect 254504 623070 254794 623098
rect 260208 623070 260590 623098
rect 263612 623070 263810 623098
rect 269224 623070 269606 623098
rect 271892 623070 272182 623098
rect 275112 623070 275402 623098
rect 277688 623070 277978 623098
rect 237406 622934 237604 622962
rect 228732 622872 228784 622878
rect 228784 622820 229034 622826
rect 228732 622814 229034 622820
rect 228744 622798 229034 622814
rect 257632 622810 258014 622826
rect 257620 622804 258014 622810
rect 257672 622798 258014 622804
rect 257620 622746 257672 622752
rect 222844 622736 222896 622742
rect 222896 622684 223238 622690
rect 222844 622678 223238 622684
rect 222856 622662 223238 622678
rect 240336 622674 240626 622690
rect 240324 622668 240626 622674
rect 240376 622662 240626 622668
rect 240324 622610 240376 622616
rect 248696 622600 248748 622606
rect 248748 622548 248998 622554
rect 248696 622542 248998 622548
rect 248708 622526 248998 622542
rect 266280 622538 266386 622554
rect 280724 622538 280752 629954
rect 266268 622532 266386 622538
rect 266320 622526 266386 622532
rect 280712 622532 280764 622538
rect 266268 622474 266320 622480
rect 280712 622474 280764 622480
rect 219728 622402 220018 622418
rect 219716 622396 220018 622402
rect 219768 622390 220018 622396
rect 280554 622390 280844 622418
rect 219716 622338 219768 622344
rect 280712 622328 280764 622334
rect 280712 622270 280764 622276
rect 219636 615466 219756 615494
rect 219728 563054 219756 615466
rect 219728 563026 219848 563054
rect 219348 559088 219400 559094
rect 219348 559030 219400 559036
rect 219256 557524 219308 557530
rect 219256 557466 219308 557472
rect 219532 553648 219584 553654
rect 219532 553590 219584 553596
rect 219164 544536 219216 544542
rect 219164 544478 219216 544484
rect 219544 543726 219572 553590
rect 219820 553394 219848 563026
rect 220176 560312 220228 560318
rect 220176 560254 220228 560260
rect 219912 560102 220018 560130
rect 219912 553654 219940 560102
rect 219900 553648 219952 553654
rect 219900 553590 219952 553596
rect 220188 553394 220216 560254
rect 222594 560102 222976 560130
rect 222200 559360 222252 559366
rect 222200 559302 222252 559308
rect 219728 553366 219848 553394
rect 220096 553366 220216 553394
rect 219728 543946 219756 553366
rect 219728 543918 220032 543946
rect 219532 543720 219584 543726
rect 219532 543662 219584 543668
rect 219256 543652 219308 543658
rect 219256 543594 219308 543600
rect 218704 543040 218756 543046
rect 218704 542982 218756 542988
rect 219268 539963 219296 543594
rect 220004 539963 220032 543918
rect 220096 543114 220124 553366
rect 220728 544468 220780 544474
rect 220728 544410 220780 544416
rect 220084 543108 220136 543114
rect 220084 543050 220136 543056
rect 220740 539963 220768 544410
rect 222212 543930 222240 559302
rect 222292 558544 222344 558550
rect 222292 558486 222344 558492
rect 222200 543924 222252 543930
rect 222200 543866 222252 543872
rect 221464 543720 221516 543726
rect 221464 543662 221516 543668
rect 221476 539963 221504 543662
rect 222304 540138 222332 558486
rect 222948 557598 222976 560102
rect 225064 560102 225170 560130
rect 228008 560102 228390 560130
rect 230492 560102 230966 560130
rect 233896 560102 234186 560130
rect 236012 560102 236762 560130
rect 238772 560102 239982 560130
rect 241532 560102 242558 560130
rect 245672 560102 245778 560130
rect 247052 560102 248354 560130
rect 251192 560102 251574 560130
rect 253952 560102 254150 560130
rect 257080 560102 257370 560130
rect 259656 560102 259946 560130
rect 262784 560102 263166 560130
rect 265360 560102 265742 560130
rect 268672 560102 268962 560130
rect 271248 560102 271538 560130
rect 274652 560102 274758 560130
rect 276952 560102 277334 560130
rect 280264 560102 280554 560130
rect 223580 559088 223632 559094
rect 223580 559030 223632 559036
rect 222936 557592 222988 557598
rect 222936 557534 222988 557540
rect 222844 543924 222896 543930
rect 222844 543866 222896 543872
rect 222228 540110 222332 540138
rect 222228 539920 222256 540110
rect 222856 539963 222884 543866
rect 223592 539963 223620 559030
rect 224408 557592 224460 557598
rect 224408 557534 224460 557540
rect 223672 557524 223724 557530
rect 223672 557466 223724 557472
rect 223684 543946 223712 557466
rect 223684 543918 224356 543946
rect 224328 539963 224356 543918
rect 224420 543726 224448 557534
rect 225064 550118 225092 560102
rect 228008 558822 228036 560102
rect 225144 558816 225196 558822
rect 225144 558758 225196 558764
rect 227996 558816 228048 558822
rect 227996 558758 228048 558764
rect 225052 550112 225104 550118
rect 225052 550054 225104 550060
rect 224408 543720 224460 543726
rect 224408 543662 224460 543668
rect 225156 540138 225184 558758
rect 227720 558272 227772 558278
rect 227720 558214 227772 558220
rect 226432 552968 226484 552974
rect 226432 552910 226484 552916
rect 225788 543720 225840 543726
rect 225788 543662 225840 543668
rect 225080 540110 225184 540138
rect 225080 539920 225108 540110
rect 225800 539963 225828 543662
rect 226444 539963 226472 552910
rect 227168 544536 227220 544542
rect 227168 544478 227220 544484
rect 227180 539963 227208 544478
rect 227732 543946 227760 558214
rect 230492 557534 230520 560102
rect 231952 558612 232004 558618
rect 231952 558554 232004 558560
rect 231964 557534 231992 558554
rect 233896 558414 233924 560102
rect 233884 558408 233936 558414
rect 233884 558350 233936 558356
rect 230492 557506 230796 557534
rect 231964 557506 232268 557534
rect 228640 555688 228692 555694
rect 228640 555630 228692 555636
rect 227732 543918 227944 543946
rect 227916 539963 227944 543918
rect 228652 539963 228680 555630
rect 229284 554192 229336 554198
rect 229284 554134 229336 554140
rect 229296 539963 229324 554134
rect 230020 543244 230072 543250
rect 230020 543186 230072 543192
rect 230032 539963 230060 543186
rect 230768 539963 230796 557506
rect 231492 543244 231544 543250
rect 231492 543186 231544 543192
rect 231504 539963 231532 543186
rect 232240 539963 232268 557506
rect 236012 547398 236040 560102
rect 236000 547392 236052 547398
rect 236000 547334 236052 547340
rect 235080 547324 235132 547330
rect 235080 547266 235132 547272
rect 234344 545760 234396 545766
rect 234344 545702 234396 545708
rect 232872 543108 232924 543114
rect 232872 543050 232924 543056
rect 232884 539963 232912 543050
rect 233608 543040 233660 543046
rect 233608 542982 233660 542988
rect 233620 539963 233648 542982
rect 234356 539963 234384 545702
rect 235092 539963 235120 547266
rect 237932 543788 237984 543794
rect 237932 543730 237984 543736
rect 237196 542428 237248 542434
rect 237196 542370 237248 542376
rect 236460 541884 236512 541890
rect 236460 541826 236512 541832
rect 235816 541816 235868 541822
rect 235816 541758 235868 541764
rect 235828 539963 235856 541758
rect 236472 539963 236500 541826
rect 237208 539963 237236 542370
rect 237944 539963 237972 543730
rect 238772 543250 238800 560102
rect 241532 545970 241560 560102
rect 245672 558278 245700 560102
rect 245660 558272 245712 558278
rect 245660 558214 245712 558220
rect 242900 555620 242952 555626
rect 242900 555562 242952 555568
rect 241520 545964 241572 545970
rect 241520 545906 241572 545912
rect 242256 545148 242308 545154
rect 242256 545090 242308 545096
rect 238760 543244 238812 543250
rect 238760 543186 238812 543192
rect 238666 543144 238722 543153
rect 238666 543079 238722 543088
rect 239404 543108 239456 543114
rect 238680 539963 238708 543079
rect 239404 543050 239456 543056
rect 239416 539963 239444 543050
rect 240784 543040 240836 543046
rect 240784 542982 240836 542988
rect 240048 541340 240100 541346
rect 240048 541282 240100 541288
rect 240060 539963 240088 541282
rect 240796 539963 240824 542982
rect 241518 542736 241574 542745
rect 241518 542671 241574 542680
rect 241532 539963 241560 542671
rect 242268 539963 242296 545090
rect 242912 539963 242940 555562
rect 246488 550180 246540 550186
rect 246488 550122 246540 550128
rect 245108 550112 245160 550118
rect 245108 550054 245160 550060
rect 243636 541544 243688 541550
rect 243636 541486 243688 541492
rect 243648 539963 243676 541486
rect 244372 541476 244424 541482
rect 244372 541418 244424 541424
rect 244384 539963 244412 541418
rect 245120 539963 245148 550054
rect 245842 543008 245898 543017
rect 245842 542943 245898 542952
rect 245856 539963 245884 542943
rect 246500 539963 246528 550122
rect 247052 544474 247080 560102
rect 251192 558482 251220 560102
rect 253952 558550 253980 560102
rect 255964 560040 256016 560046
rect 255964 559982 256016 559988
rect 253940 558544 253992 558550
rect 253940 558486 253992 558492
rect 251180 558476 251232 558482
rect 251180 558418 251232 558424
rect 249800 558272 249852 558278
rect 249800 558214 249852 558220
rect 249812 557534 249840 558214
rect 249812 557506 250852 557534
rect 247960 552832 248012 552838
rect 247960 552774 248012 552780
rect 247040 544468 247092 544474
rect 247040 544410 247092 544416
rect 247224 541068 247276 541074
rect 247224 541010 247276 541016
rect 247236 539963 247264 541010
rect 247972 539963 248000 552774
rect 250076 545964 250128 545970
rect 250076 545906 250128 545912
rect 248694 542872 248750 542881
rect 248694 542807 248750 542816
rect 248708 539963 248736 542807
rect 249432 541136 249484 541142
rect 249432 541078 249484 541084
rect 249444 539963 249472 541078
rect 250088 539963 250116 545906
rect 250824 539963 250852 557506
rect 255320 552900 255372 552906
rect 255320 552842 255372 552848
rect 253664 551540 253716 551546
rect 253664 551482 253716 551488
rect 251548 548548 251600 548554
rect 251548 548490 251600 548496
rect 251560 539963 251588 548490
rect 252284 543856 252336 543862
rect 252284 543798 252336 543804
rect 252296 539963 252324 543798
rect 252928 543312 252980 543318
rect 252928 543254 252980 543260
rect 252940 539963 252968 543254
rect 253676 539963 253704 551482
rect 255332 543930 255360 552842
rect 255320 543924 255372 543930
rect 255320 543866 255372 543872
rect 255976 543182 256004 559982
rect 257080 558346 257108 560102
rect 258080 559836 258132 559842
rect 258080 559778 258132 559784
rect 257068 558340 257120 558346
rect 257068 558282 257120 558288
rect 258092 557534 258120 559778
rect 259656 558618 259684 560102
rect 260840 559904 260892 559910
rect 260840 559846 260892 559852
rect 260104 558816 260156 558822
rect 260104 558758 260156 558764
rect 259644 558612 259696 558618
rect 259644 558554 259696 558560
rect 258092 557506 258764 557534
rect 256516 543924 256568 543930
rect 256516 543866 256568 543872
rect 255964 543176 256016 543182
rect 255964 543118 256016 543124
rect 255134 542464 255190 542473
rect 255134 542399 255190 542408
rect 254400 541272 254452 541278
rect 254400 541214 254452 541220
rect 254412 539963 254440 541214
rect 255148 539963 255176 542399
rect 255872 541408 255924 541414
rect 255872 541350 255924 541356
rect 255884 539963 255912 541350
rect 256528 539963 256556 543866
rect 257252 543380 257304 543386
rect 257252 543322 257304 543328
rect 257264 539963 257292 543322
rect 257988 543176 258040 543182
rect 257988 543118 258040 543124
rect 258000 539963 258028 543118
rect 258736 539963 258764 557506
rect 259460 551608 259512 551614
rect 259460 551550 259512 551556
rect 259472 539963 259500 551550
rect 260116 545902 260144 558758
rect 260852 557534 260880 559846
rect 262784 558822 262812 560102
rect 262772 558816 262824 558822
rect 262772 558758 262824 558764
rect 265360 557938 265388 560102
rect 264244 557932 264296 557938
rect 264244 557874 264296 557880
rect 265348 557932 265400 557938
rect 265348 557874 265400 557880
rect 262864 557660 262916 557666
rect 262864 557602 262916 557608
rect 260852 557506 261616 557534
rect 260196 547460 260248 547466
rect 260196 547402 260248 547408
rect 260104 545896 260156 545902
rect 260104 545838 260156 545844
rect 260208 540138 260236 547402
rect 260840 541612 260892 541618
rect 260840 541554 260892 541560
rect 260132 540110 260236 540138
rect 260132 539920 260160 540110
rect 260852 539963 260880 541554
rect 261588 539963 261616 557506
rect 262876 549982 262904 557602
rect 262864 549976 262916 549982
rect 262864 549918 262916 549924
rect 264256 548622 264284 557874
rect 268672 557666 268700 560102
rect 269120 558340 269172 558346
rect 269120 558282 269172 558288
rect 268660 557660 268712 557666
rect 268660 557602 268712 557608
rect 267740 557592 267792 557598
rect 267740 557534 267792 557540
rect 269132 557534 269160 558282
rect 267752 557506 268056 557534
rect 269132 557506 269528 557534
rect 266544 554260 266596 554266
rect 266544 554202 266596 554208
rect 264244 548616 264296 548622
rect 264244 548558 264296 548564
rect 263692 547392 263744 547398
rect 263692 547334 263744 547340
rect 263048 541680 263100 541686
rect 263048 541622 263100 541628
rect 262312 540184 262364 540190
rect 262312 540126 262364 540132
rect 262324 539963 262352 540126
rect 263060 539963 263088 541622
rect 263704 539963 263732 547334
rect 264426 541104 264482 541113
rect 264426 541039 264482 541048
rect 264440 539963 264468 541039
rect 265900 540388 265952 540394
rect 265900 540330 265952 540336
rect 265164 540320 265216 540326
rect 265164 540262 265216 540268
rect 265176 539963 265204 540262
rect 265912 539963 265940 540330
rect 266556 539963 266584 554202
rect 267280 544536 267332 544542
rect 267280 544478 267332 544484
rect 267292 539963 267320 544478
rect 268028 539963 268056 557506
rect 268752 541748 268804 541754
rect 268752 541690 268804 541696
rect 268764 539963 268792 541690
rect 269500 539963 269528 557506
rect 271248 552702 271276 560102
rect 273260 559972 273312 559978
rect 273260 559914 273312 559920
rect 271236 552696 271288 552702
rect 271236 552638 271288 552644
rect 270132 544604 270184 544610
rect 270132 544546 270184 544552
rect 270144 539963 270172 544546
rect 271604 544468 271656 544474
rect 271604 544410 271656 544416
rect 270868 542700 270920 542706
rect 270868 542642 270920 542648
rect 270880 539963 270908 542642
rect 271616 539963 271644 544410
rect 273272 543930 273300 559914
rect 274652 547262 274680 560102
rect 276952 558210 276980 560102
rect 280264 558822 280292 560102
rect 278044 558816 278096 558822
rect 278044 558758 278096 558764
rect 280252 558816 280304 558822
rect 280252 558758 280304 558764
rect 276940 558204 276992 558210
rect 276940 558146 276992 558152
rect 274640 547256 274692 547262
rect 274640 547198 274692 547204
rect 275192 545896 275244 545902
rect 275192 545838 275244 545844
rect 273260 543924 273312 543930
rect 273260 543866 273312 543872
rect 274456 543924 274508 543930
rect 274456 543866 274508 543872
rect 273720 542632 273772 542638
rect 273720 542574 273772 542580
rect 272340 541000 272392 541006
rect 272340 540942 272392 540948
rect 272352 539963 272380 540942
rect 273076 540252 273128 540258
rect 273076 540194 273128 540200
rect 273088 539963 273116 540194
rect 273732 539963 273760 542574
rect 274468 539963 274496 543866
rect 275204 539963 275232 545838
rect 278056 545834 278084 558758
rect 279516 552696 279568 552702
rect 279516 552638 279568 552644
rect 278044 545828 278096 545834
rect 278044 545770 278096 545776
rect 276572 543244 276624 543250
rect 276572 543186 276624 543192
rect 275928 542768 275980 542774
rect 275928 542710 275980 542716
rect 275940 539963 275968 542710
rect 276584 539963 276612 543186
rect 278044 542904 278096 542910
rect 278044 542846 278096 542852
rect 277308 542836 277360 542842
rect 277308 542778 277360 542784
rect 277320 539963 277348 542778
rect 278056 539963 278084 542846
rect 278780 540456 278832 540462
rect 278780 540398 278832 540404
rect 278792 539963 278820 540398
rect 279528 539963 279556 552638
rect 280724 547874 280752 622270
rect 280816 552974 280844 622390
rect 280894 594960 280950 594969
rect 280894 594895 280950 594904
rect 280804 552968 280856 552974
rect 280804 552910 280856 552916
rect 280908 551478 280936 594895
rect 280896 551472 280948 551478
rect 280896 551414 280948 551420
rect 280724 547846 280936 547874
rect 280160 542972 280212 542978
rect 280160 542914 280212 542920
rect 280172 539963 280200 542914
rect 280908 539963 280936 547846
rect 281000 543182 281028 633626
rect 281080 633616 281132 633622
rect 281080 633558 281132 633564
rect 280988 543176 281040 543182
rect 280988 543118 281040 543124
rect 281092 543114 281120 633558
rect 289820 633548 289872 633554
rect 289820 633490 289872 633496
rect 288440 633480 288492 633486
rect 288440 633422 288492 633428
rect 284944 631372 284996 631378
rect 284944 631314 284996 631320
rect 281630 619984 281686 619993
rect 281630 619919 281686 619928
rect 281170 592784 281226 592793
rect 281170 592719 281226 592728
rect 281184 550050 281212 592719
rect 281538 568304 281594 568313
rect 281538 568239 281594 568248
rect 281262 564904 281318 564913
rect 281262 564839 281318 564848
rect 281276 554198 281304 564839
rect 281552 562290 281580 568239
rect 281540 562284 281592 562290
rect 281540 562226 281592 562232
rect 281538 562184 281594 562193
rect 281538 562119 281594 562128
rect 281552 559774 281580 562119
rect 281540 559768 281592 559774
rect 281540 559710 281592 559716
rect 281644 556918 281672 619919
rect 281722 617264 281778 617273
rect 281722 617199 281778 617208
rect 281632 556912 281684 556918
rect 281632 556854 281684 556860
rect 281736 555694 281764 617199
rect 283010 613864 283066 613873
rect 283010 613799 283066 613808
rect 281998 611144 282054 611153
rect 281998 611079 282054 611088
rect 281814 586664 281870 586673
rect 281814 586599 281870 586608
rect 281724 555688 281776 555694
rect 281724 555630 281776 555636
rect 281828 555558 281856 586599
rect 281906 577144 281962 577153
rect 281906 577079 281962 577088
rect 281816 555552 281868 555558
rect 281816 555494 281868 555500
rect 281264 554192 281316 554198
rect 281264 554134 281316 554140
rect 281920 551342 281948 577079
rect 281908 551336 281960 551342
rect 281908 551278 281960 551284
rect 281172 550044 281224 550050
rect 281172 549986 281224 549992
rect 282012 544406 282040 611079
rect 282918 574424 282974 574433
rect 282918 574359 282974 574368
rect 282092 562284 282144 562290
rect 282092 562226 282144 562232
rect 282104 559638 282132 562226
rect 282932 560046 282960 574359
rect 282920 560040 282972 560046
rect 282920 559982 282972 559988
rect 283024 559706 283052 613799
rect 283654 607744 283710 607753
rect 283654 607679 283710 607688
rect 283102 605024 283158 605033
rect 283102 604959 283158 604968
rect 283012 559700 283064 559706
rect 283012 559642 283064 559648
rect 282092 559632 282144 559638
rect 282092 559574 282144 559580
rect 283116 554130 283144 604959
rect 283194 601624 283250 601633
rect 283194 601559 283250 601568
rect 283104 554124 283156 554130
rect 283104 554066 283156 554072
rect 283208 554062 283236 601559
rect 283286 598904 283342 598913
rect 283286 598839 283342 598848
rect 283196 554056 283248 554062
rect 283196 553998 283248 554004
rect 283300 552770 283328 598839
rect 283562 589384 283618 589393
rect 283562 589319 283564 589328
rect 283616 589319 283618 589328
rect 283564 589290 283616 589296
rect 283378 583264 283434 583273
rect 283378 583199 283434 583208
rect 283288 552764 283340 552770
rect 283288 552706 283340 552712
rect 283392 549914 283420 583199
rect 283470 580544 283526 580553
rect 283470 580479 283526 580488
rect 283484 551410 283512 580479
rect 283562 571024 283618 571033
rect 283562 570959 283618 570968
rect 283576 556986 283604 570959
rect 283564 556980 283616 556986
rect 283564 556922 283616 556928
rect 283472 551404 283524 551410
rect 283472 551346 283524 551352
rect 283380 549908 283432 549914
rect 283380 549850 283432 549856
rect 282368 547256 282420 547262
rect 282368 547198 282420 547204
rect 282000 544400 282052 544406
rect 282000 544342 282052 544348
rect 281080 543108 281132 543114
rect 281080 543050 281132 543056
rect 281632 542496 281684 542502
rect 281632 542438 281684 542444
rect 281644 539963 281672 542438
rect 282380 539963 282408 547198
rect 283668 547194 283696 607679
rect 283748 547528 283800 547534
rect 283748 547470 283800 547476
rect 283656 547188 283708 547194
rect 283656 547130 283708 547136
rect 282920 542428 282972 542434
rect 282920 542370 282972 542376
rect 282932 541657 282960 542370
rect 282918 541648 282974 541657
rect 282918 541583 282974 541592
rect 283104 541204 283156 541210
rect 283104 541146 283156 541152
rect 283116 539963 283144 541146
rect 283760 539963 283788 547470
rect 284956 543046 284984 631314
rect 286324 615528 286376 615534
rect 286324 615470 286376 615476
rect 286336 559570 286364 615470
rect 286416 596216 286468 596222
rect 286416 596158 286468 596164
rect 286324 559564 286376 559570
rect 286324 559506 286376 559512
rect 286428 544610 286456 596158
rect 287704 576904 287756 576910
rect 287704 576846 287756 576852
rect 286508 571396 286560 571402
rect 286508 571338 286560 571344
rect 286520 547466 286548 571338
rect 287716 558346 287744 576846
rect 287704 558340 287756 558346
rect 287704 558282 287756 558288
rect 286508 547460 286560 547466
rect 286508 547402 286560 547408
rect 288072 545284 288124 545290
rect 288072 545226 288124 545232
rect 286692 545216 286744 545222
rect 286692 545158 286744 545164
rect 286416 544604 286468 544610
rect 286416 544546 286468 544552
rect 285220 543924 285272 543930
rect 285220 543866 285272 543872
rect 284944 543040 284996 543046
rect 284944 542982 284996 542988
rect 284484 542428 284536 542434
rect 284484 542370 284536 542376
rect 284496 539963 284524 542370
rect 285232 539963 285260 543866
rect 285956 542564 286008 542570
rect 285956 542506 286008 542512
rect 285968 539963 285996 542506
rect 286704 539963 286732 545158
rect 287336 540524 287388 540530
rect 287336 540466 287388 540472
rect 287348 539963 287376 540466
rect 288084 539963 288112 545226
rect 288452 543946 288480 633422
rect 288532 631032 288584 631038
rect 288532 630974 288584 630980
rect 288544 544082 288572 630974
rect 289084 600364 289136 600370
rect 289084 600306 289136 600312
rect 289096 545970 289124 600306
rect 289832 557534 289860 633490
rect 289832 557506 290228 557534
rect 289084 545964 289136 545970
rect 289084 545906 289136 545912
rect 288544 544054 289584 544082
rect 288452 543918 288848 543946
rect 288820 539963 288848 543918
rect 289556 539963 289584 544054
rect 290200 539963 290228 557506
rect 290924 544060 290976 544066
rect 290924 544002 290976 544008
rect 290936 539963 290964 544002
rect 291212 543946 291240 634782
rect 295984 632868 296036 632874
rect 295984 632810 296036 632816
rect 291292 632800 291344 632806
rect 291292 632742 291344 632748
rect 291304 557534 291332 632742
rect 293960 631100 294012 631106
rect 293960 631042 294012 631048
rect 291844 582412 291896 582418
rect 291844 582354 291896 582360
rect 291856 561134 291884 582354
rect 291844 561128 291896 561134
rect 291844 561070 291896 561076
rect 291304 557506 292436 557534
rect 291212 543918 291700 543946
rect 291672 539963 291700 543918
rect 292408 539963 292436 557506
rect 293972 543998 294000 631042
rect 295996 544542 296024 632810
rect 298100 631236 298152 631242
rect 298100 631178 298152 631184
rect 296812 631168 296864 631174
rect 296812 631110 296864 631116
rect 296720 630896 296772 630902
rect 296720 630838 296772 630844
rect 295984 544536 296036 544542
rect 295984 544478 296036 544484
rect 293960 543992 294012 543998
rect 293960 543934 294012 543940
rect 295248 543992 295300 543998
rect 295248 543934 295300 543940
rect 293130 542600 293186 542609
rect 293130 542535 293186 542544
rect 293144 539963 293172 542535
rect 294510 541240 294566 541249
rect 294510 541175 294566 541184
rect 293776 540660 293828 540666
rect 293776 540602 293828 540608
rect 293788 539963 293816 540602
rect 294524 539963 294552 541175
rect 295260 539963 295288 543934
rect 295984 543108 296036 543114
rect 295984 543050 296036 543056
rect 295996 539963 296024 543050
rect 296732 539963 296760 630838
rect 296824 557534 296852 631110
rect 298112 557534 298140 631178
rect 302884 619676 302936 619682
rect 302884 619618 302936 619624
rect 302240 589348 302292 589354
rect 302240 589290 302292 589296
rect 300124 586560 300176 586566
rect 300124 586502 300176 586508
rect 296824 557506 297404 557534
rect 298112 557506 298876 557534
rect 297376 539963 297404 557506
rect 298100 543176 298152 543182
rect 298100 543118 298152 543124
rect 298112 539963 298140 543118
rect 298848 539963 298876 557506
rect 300136 547262 300164 586502
rect 302252 560250 302280 589290
rect 302240 560244 302292 560250
rect 302240 560186 302292 560192
rect 302252 559706 302280 560186
rect 302240 559700 302292 559706
rect 302240 559642 302292 559648
rect 302896 552702 302924 619618
rect 304264 605872 304316 605878
rect 304264 605814 304316 605820
rect 302976 559700 303028 559706
rect 302976 559642 303028 559648
rect 302884 552696 302936 552702
rect 302884 552638 302936 552644
rect 300124 547256 300176 547262
rect 300124 547198 300176 547204
rect 300584 543380 300636 543386
rect 300584 543322 300636 543328
rect 300216 543312 300268 543318
rect 300216 543254 300268 543260
rect 299572 543040 299624 543046
rect 299572 542982 299624 542988
rect 299584 539963 299612 542982
rect 300124 542564 300176 542570
rect 300124 542506 300176 542512
rect 300136 517342 300164 542506
rect 300228 518158 300256 543254
rect 300400 542904 300452 542910
rect 300400 542846 300452 542852
rect 300308 542700 300360 542706
rect 300308 542642 300360 542648
rect 300320 520062 300348 542642
rect 300308 520056 300360 520062
rect 300308 519998 300360 520004
rect 300412 519994 300440 542846
rect 300492 541000 300544 541006
rect 300492 540942 300544 540948
rect 300400 519988 300452 519994
rect 300400 519930 300452 519936
rect 300216 518152 300268 518158
rect 300216 518094 300268 518100
rect 300504 518022 300532 540942
rect 300596 519926 300624 543322
rect 301688 542972 301740 542978
rect 301688 542914 301740 542920
rect 301594 542872 301650 542881
rect 301594 542807 301650 542816
rect 301412 542428 301464 542434
rect 301412 542370 301464 542376
rect 300676 541544 300728 541550
rect 300676 541486 300728 541492
rect 300688 529922 300716 541486
rect 301424 538214 301452 542370
rect 301504 540456 301556 540462
rect 301504 540398 301556 540404
rect 301516 539578 301544 540398
rect 301504 539572 301556 539578
rect 301504 539514 301556 539520
rect 301424 538186 301544 538214
rect 300676 529916 300728 529922
rect 300676 529858 300728 529864
rect 300584 519920 300636 519926
rect 300584 519862 300636 519868
rect 300492 518016 300544 518022
rect 300492 517958 300544 517964
rect 300124 517336 300176 517342
rect 300124 517278 300176 517284
rect 301516 517206 301544 538186
rect 301608 518809 301636 542807
rect 301700 519790 301728 542914
rect 301964 542836 302016 542842
rect 301964 542778 302016 542784
rect 301872 542768 301924 542774
rect 301872 542710 301924 542716
rect 301780 541748 301832 541754
rect 301780 541690 301832 541696
rect 301688 519784 301740 519790
rect 301688 519726 301740 519732
rect 301594 518800 301650 518809
rect 301594 518735 301650 518744
rect 301792 518498 301820 541690
rect 301884 519246 301912 542710
rect 301976 519858 302004 542778
rect 302884 542496 302936 542502
rect 302884 542438 302936 542444
rect 302056 541680 302108 541686
rect 302056 541622 302108 541628
rect 301964 519852 302016 519858
rect 301964 519794 302016 519800
rect 301872 519240 301924 519246
rect 301872 519182 301924 519188
rect 302068 518634 302096 541622
rect 302238 532400 302294 532409
rect 302238 532335 302294 532344
rect 302252 532234 302280 532335
rect 302240 532228 302292 532234
rect 302240 532170 302292 532176
rect 302896 518894 302924 542438
rect 302988 520198 303016 559642
rect 304276 547534 304304 605814
rect 304264 547528 304316 547534
rect 304264 547470 304316 547476
rect 304264 543108 304316 543114
rect 304264 543050 304316 543056
rect 303068 541476 303120 541482
rect 303068 541418 303120 541424
rect 302976 520192 303028 520198
rect 302976 520134 303028 520140
rect 302804 518866 302924 518894
rect 302056 518628 302108 518634
rect 302056 518570 302108 518576
rect 301780 518492 301832 518498
rect 301780 518434 301832 518440
rect 301504 517200 301556 517206
rect 301504 517142 301556 517148
rect 302804 517138 302832 518866
rect 302882 517440 302938 517449
rect 302882 517375 302938 517384
rect 302792 517132 302844 517138
rect 302792 517074 302844 517080
rect 302896 516186 302924 517375
rect 302884 516180 302936 516186
rect 302884 516122 302936 516128
rect 57702 509960 57758 509969
rect 41328 509924 41380 509930
rect 57702 509895 57704 509904
rect 41328 509866 41380 509872
rect 57756 509895 57758 509904
rect 57886 509960 57942 509969
rect 57886 509895 57942 509904
rect 57704 509866 57756 509872
rect 40960 469124 41012 469130
rect 40960 469066 41012 469072
rect 40868 469056 40920 469062
rect 40868 468998 40920 469004
rect 40776 465656 40828 465662
rect 40776 465598 40828 465604
rect 40788 373862 40816 465598
rect 40880 373969 40908 468998
rect 40866 373960 40922 373969
rect 40866 373895 40922 373904
rect 40776 373856 40828 373862
rect 40776 373798 40828 373804
rect 40972 371210 41000 469066
rect 41052 468784 41104 468790
rect 41052 468726 41104 468732
rect 40960 371204 41012 371210
rect 40960 371146 41012 371152
rect 40684 202836 40736 202842
rect 40684 202778 40736 202784
rect 41064 164286 41092 468726
rect 41144 460352 41196 460358
rect 41144 460294 41196 460300
rect 41052 164280 41104 164286
rect 41052 164222 41104 164228
rect 41156 57730 41184 460294
rect 41236 460284 41288 460290
rect 41236 460226 41288 460232
rect 41248 57798 41276 460226
rect 41340 382226 41368 509866
rect 302988 502489 303016 520134
rect 303080 518090 303108 541418
rect 303160 541340 303212 541346
rect 303160 541282 303212 541288
rect 303172 525774 303200 541282
rect 303160 525768 303212 525774
rect 303160 525710 303212 525716
rect 303068 518084 303120 518090
rect 303068 518026 303120 518032
rect 304276 517478 304304 543050
rect 304356 542632 304408 542638
rect 304356 542574 304408 542580
rect 304368 519110 304396 542574
rect 304448 541884 304500 541890
rect 304448 541826 304500 541832
rect 304460 535430 304488 541826
rect 304448 535424 304500 535430
rect 304448 535366 304500 535372
rect 304448 532228 304500 532234
rect 304448 532170 304500 532176
rect 304356 519104 304408 519110
rect 304356 519046 304408 519052
rect 304264 517472 304316 517478
rect 304264 517414 304316 517420
rect 304460 515438 304488 532170
rect 305656 519178 305684 700334
rect 317052 639600 317104 639606
rect 317052 639542 317104 639548
rect 316960 634976 317012 634982
rect 316960 634918 317012 634924
rect 316868 634908 316920 634914
rect 316868 634850 316920 634856
rect 313924 633004 313976 633010
rect 313924 632946 313976 632952
rect 309784 632936 309836 632942
rect 309784 632878 309836 632884
rect 307024 610020 307076 610026
rect 307024 609962 307076 609968
rect 307036 550186 307064 609962
rect 307024 550180 307076 550186
rect 307024 550122 307076 550128
rect 309796 547398 309824 632878
rect 311164 632664 311216 632670
rect 311164 632606 311216 632612
rect 311176 554266 311204 632606
rect 312544 632528 312596 632534
rect 312544 632470 312596 632476
rect 311164 554260 311216 554266
rect 311164 554202 311216 554208
rect 312556 550118 312584 632470
rect 312544 550112 312596 550118
rect 312544 550054 312596 550060
rect 309784 547392 309836 547398
rect 309784 547334 309836 547340
rect 313936 545902 313964 632946
rect 316776 632392 316828 632398
rect 316776 632334 316828 632340
rect 316684 632324 316736 632330
rect 316684 632266 316736 632272
rect 315302 632224 315358 632233
rect 315302 632159 315358 632168
rect 314016 629332 314068 629338
rect 314016 629274 314068 629280
rect 314028 551614 314056 629274
rect 315316 552906 315344 632159
rect 315304 552900 315356 552906
rect 315304 552842 315356 552848
rect 314016 551608 314068 551614
rect 314016 551550 314068 551556
rect 316696 551546 316724 632266
rect 316788 555626 316816 632334
rect 316880 559910 316908 634850
rect 316868 559904 316920 559910
rect 316868 559846 316920 559852
rect 316972 559842 317000 634918
rect 317064 568313 317092 639542
rect 364352 635526 364380 702406
rect 401140 636880 401192 636886
rect 401140 636822 401192 636828
rect 364340 635520 364392 635526
rect 364340 635462 364392 635468
rect 318800 634092 318852 634098
rect 318800 634034 318852 634040
rect 318248 632188 318300 632194
rect 318248 632130 318300 632136
rect 318064 631304 318116 631310
rect 318064 631246 318116 631252
rect 317786 629640 317842 629649
rect 317786 629575 317842 629584
rect 317800 629338 317828 629575
rect 317788 629332 317840 629338
rect 317788 629274 317840 629280
rect 317970 620120 318026 620129
rect 317970 620055 318026 620064
rect 317984 619682 318012 620055
rect 317972 619676 318024 619682
rect 317972 619618 318024 619624
rect 317970 615632 318026 615641
rect 317970 615567 318026 615576
rect 317984 615534 318012 615567
rect 317972 615528 318024 615534
rect 317972 615470 318024 615476
rect 317878 610600 317934 610609
rect 317878 610535 317934 610544
rect 317892 610026 317920 610535
rect 317880 610020 317932 610026
rect 317880 609962 317932 609968
rect 317970 606112 318026 606121
rect 317970 606047 318026 606056
rect 317984 605878 318012 606047
rect 317972 605872 318024 605878
rect 317972 605814 318024 605820
rect 317602 601080 317658 601089
rect 317602 601015 317658 601024
rect 317616 600370 317644 601015
rect 317604 600364 317656 600370
rect 317604 600306 317656 600312
rect 317602 596456 317658 596465
rect 317602 596391 317658 596400
rect 317616 596222 317644 596391
rect 317604 596216 317656 596222
rect 317604 596158 317656 596164
rect 317420 586560 317472 586566
rect 317418 586528 317420 586537
rect 317472 586528 317474 586537
rect 317418 586463 317474 586472
rect 317970 582584 318026 582593
rect 317970 582519 318026 582528
rect 317984 582418 318012 582519
rect 317972 582412 318024 582418
rect 317972 582354 318024 582360
rect 317878 577280 317934 577289
rect 317878 577215 317934 577224
rect 317892 576910 317920 577215
rect 317880 576904 317932 576910
rect 317880 576846 317932 576852
rect 317970 571840 318026 571849
rect 317970 571775 318026 571784
rect 317984 571402 318012 571775
rect 317972 571396 318024 571402
rect 317972 571338 318024 571344
rect 317050 568304 317106 568313
rect 317050 568239 317106 568248
rect 316960 559836 317012 559842
rect 316960 559778 317012 559784
rect 317418 557696 317474 557705
rect 317418 557631 317474 557640
rect 317432 557598 317460 557631
rect 317420 557592 317472 557598
rect 317420 557534 317472 557540
rect 316776 555620 316828 555626
rect 316776 555562 316828 555568
rect 317970 553480 318026 553489
rect 317970 553415 317972 553424
rect 318024 553415 318026 553424
rect 317972 553386 318024 553392
rect 316684 551540 316736 551546
rect 316684 551482 316736 551488
rect 317512 549228 317564 549234
rect 317512 549170 317564 549176
rect 317524 549137 317552 549170
rect 317510 549128 317566 549137
rect 317510 549063 317566 549072
rect 313924 545896 313976 545902
rect 313924 545838 313976 545844
rect 314200 545284 314252 545290
rect 314200 545226 314252 545232
rect 314016 545216 314068 545222
rect 314016 545158 314068 545164
rect 313924 543924 313976 543930
rect 313924 543866 313976 543872
rect 307024 540388 307076 540394
rect 307024 540330 307076 540336
rect 305644 519172 305696 519178
rect 305644 519114 305696 519120
rect 307036 518430 307064 540330
rect 312544 540320 312596 540326
rect 312544 540262 312596 540268
rect 312556 518906 312584 540262
rect 312544 518900 312596 518906
rect 312544 518842 312596 518848
rect 307024 518424 307076 518430
rect 307024 518366 307076 518372
rect 313936 515914 313964 543866
rect 314028 516118 314056 545158
rect 314108 543992 314160 543998
rect 314108 543934 314160 543940
rect 314016 516112 314068 516118
rect 314016 516054 314068 516060
rect 314120 516050 314148 543934
rect 314212 520266 314240 545226
rect 316776 545148 316828 545154
rect 316776 545090 316828 545096
rect 316684 543788 316736 543794
rect 316684 543730 316736 543736
rect 314292 540592 314344 540598
rect 314292 540534 314344 540540
rect 314200 520260 314252 520266
rect 314200 520202 314252 520208
rect 314108 516044 314160 516050
rect 314108 515986 314160 515992
rect 313924 515908 313976 515914
rect 313924 515850 313976 515856
rect 314304 515846 314332 540534
rect 314384 540524 314436 540530
rect 314384 540466 314436 540472
rect 314396 515982 314424 540466
rect 314384 515976 314436 515982
rect 314384 515918 314436 515924
rect 314292 515840 314344 515846
rect 314292 515782 314344 515788
rect 304448 515432 304500 515438
rect 304448 515374 304500 515380
rect 316696 514758 316724 543730
rect 316788 515778 316816 545090
rect 317972 543856 318024 543862
rect 317970 543824 317972 543833
rect 318024 543824 318026 543833
rect 317970 543759 318026 543768
rect 317052 543176 317104 543182
rect 317052 543118 317104 543124
rect 316866 541648 316922 541657
rect 316866 541583 316922 541592
rect 316776 515772 316828 515778
rect 316776 515714 316828 515720
rect 316684 514752 316736 514758
rect 316684 514694 316736 514700
rect 316880 514690 316908 541583
rect 316960 541204 317012 541210
rect 316960 541146 317012 541152
rect 316972 515710 317000 541146
rect 317064 517274 317092 543118
rect 318076 543017 318104 631246
rect 318154 625288 318210 625297
rect 318154 625223 318210 625232
rect 318168 544474 318196 625223
rect 318260 559978 318288 632130
rect 318812 592793 318840 634034
rect 383108 633684 383160 633690
rect 383108 633626 383160 633632
rect 337384 633004 337436 633010
rect 337384 632946 337436 632952
rect 332876 632936 332928 632942
rect 332876 632878 332928 632884
rect 319536 632732 319588 632738
rect 319536 632674 319588 632680
rect 319444 630964 319496 630970
rect 319444 630906 319496 630912
rect 319076 630828 319128 630834
rect 319076 630770 319128 630776
rect 319088 629950 319116 630770
rect 319076 629944 319128 629950
rect 319076 629886 319128 629892
rect 318798 592784 318854 592793
rect 318798 592719 318854 592728
rect 319352 562352 319404 562358
rect 318338 562320 318394 562329
rect 319352 562294 319404 562300
rect 318338 562255 318394 562264
rect 318248 559972 318300 559978
rect 318248 559914 318300 559920
rect 318352 556850 318380 562255
rect 318340 556844 318392 556850
rect 318340 556786 318392 556792
rect 319364 552838 319392 562294
rect 319352 552832 319404 552838
rect 319352 552774 319404 552780
rect 318156 544468 318208 544474
rect 318156 544410 318208 544416
rect 318340 543244 318392 543250
rect 318340 543186 318392 543192
rect 318062 543008 318118 543017
rect 318062 542943 318118 542952
rect 318246 542600 318302 542609
rect 318246 542535 318302 542544
rect 317144 541612 317196 541618
rect 317144 541554 317196 541560
rect 317156 518226 317184 541554
rect 318156 541408 318208 541414
rect 318156 541350 318208 541356
rect 317234 541240 317290 541249
rect 317234 541175 317290 541184
rect 317248 520130 317276 541175
rect 317972 541136 318024 541142
rect 317972 541078 318024 541084
rect 317984 538214 318012 541078
rect 318064 539572 318116 539578
rect 318064 539514 318116 539520
rect 318076 539345 318104 539514
rect 318062 539336 318118 539345
rect 318062 539271 318118 539280
rect 317984 538186 318104 538214
rect 317604 535424 317656 535430
rect 317604 535366 317656 535372
rect 317616 534993 317644 535366
rect 317602 534984 317658 534993
rect 317602 534919 317658 534928
rect 317604 529916 317656 529922
rect 317604 529858 317656 529864
rect 317616 529825 317644 529858
rect 317602 529816 317658 529825
rect 317602 529751 317658 529760
rect 317604 525768 317656 525774
rect 317604 525710 317656 525716
rect 317616 525473 317644 525710
rect 317602 525464 317658 525473
rect 317602 525399 317658 525408
rect 317236 520124 317288 520130
rect 317236 520066 317288 520072
rect 318076 518702 318104 538186
rect 318064 518696 318116 518702
rect 318064 518638 318116 518644
rect 318168 518566 318196 541350
rect 318156 518560 318208 518566
rect 318156 518502 318208 518508
rect 317144 518220 317196 518226
rect 317144 518162 317196 518168
rect 318260 517410 318288 542535
rect 318352 519042 318380 543186
rect 319456 543046 319484 630906
rect 319548 545766 319576 632674
rect 319720 632596 319772 632602
rect 319720 632538 319772 632544
rect 319626 632360 319682 632369
rect 319626 632295 319682 632304
rect 319640 547330 319668 632295
rect 319732 548554 319760 632538
rect 319812 632460 319864 632466
rect 319812 632402 319864 632408
rect 319824 562358 319852 632402
rect 320824 632256 320876 632262
rect 320824 632198 320876 632204
rect 319904 632120 319956 632126
rect 319904 632062 319956 632068
rect 319812 562352 319864 562358
rect 319812 562294 319864 562300
rect 319916 558362 319944 632062
rect 320836 630494 320864 632198
rect 323860 632120 323912 632126
rect 323860 632062 323912 632068
rect 323872 630972 323900 632062
rect 332888 630972 332916 632878
rect 337396 630972 337424 632946
rect 378600 632868 378652 632874
rect 378600 632810 378652 632816
rect 355416 632732 355468 632738
rect 355416 632674 355468 632680
rect 350908 632664 350960 632670
rect 350908 632606 350960 632612
rect 341892 632256 341944 632262
rect 341892 632198 341944 632204
rect 341904 630972 341932 632198
rect 346398 632088 346454 632097
rect 346398 632023 346454 632032
rect 346412 630972 346440 632023
rect 350920 630972 350948 632606
rect 355428 630972 355456 632674
rect 364432 632596 364484 632602
rect 364432 632538 364484 632544
rect 359924 632528 359976 632534
rect 359924 632470 359976 632476
rect 359936 630972 359964 632470
rect 364444 630972 364472 632538
rect 373448 632460 373500 632466
rect 373448 632402 373500 632408
rect 368940 631372 368992 631378
rect 368940 631314 368992 631320
rect 368952 630972 368980 631314
rect 373460 630972 373488 632402
rect 378612 630972 378640 632810
rect 383120 630972 383148 633626
rect 387616 632392 387668 632398
rect 387616 632334 387668 632340
rect 392122 632360 392178 632369
rect 387628 630972 387656 632334
rect 392122 632295 392178 632304
rect 396632 632324 396684 632330
rect 392136 630972 392164 632295
rect 396632 632266 396684 632272
rect 396644 630972 396672 632266
rect 401152 630972 401180 636822
rect 423680 635520 423732 635526
rect 423680 635462 423732 635468
rect 419170 632224 419226 632233
rect 419170 632159 419226 632168
rect 419184 630972 419212 632159
rect 423692 630972 423720 635462
rect 428188 632188 428240 632194
rect 428188 632130 428240 632136
rect 428200 630972 428228 632130
rect 428464 631032 428516 631038
rect 428464 630974 428516 630980
rect 328090 630864 328146 630873
rect 328146 630822 328394 630850
rect 328090 630799 328146 630808
rect 409880 630760 409932 630766
rect 405370 630728 405426 630737
rect 405426 630686 405674 630714
rect 409932 630708 410182 630714
rect 409880 630702 410182 630708
rect 409892 630686 410182 630702
rect 414400 630698 414690 630714
rect 414388 630692 414690 630698
rect 405370 630663 405426 630672
rect 414440 630686 414690 630692
rect 414388 630634 414440 630640
rect 320824 630488 320876 630494
rect 320824 630430 320876 630436
rect 428476 611318 428504 630974
rect 428464 611312 428516 611318
rect 428464 611254 428516 611260
rect 319824 558334 319944 558362
rect 319824 558278 319852 558334
rect 319812 558272 319864 558278
rect 319812 558214 319864 558220
rect 428370 558240 428426 558249
rect 428370 558175 428426 558184
rect 319812 555484 319864 555490
rect 319812 555426 319864 555432
rect 319720 548548 319772 548554
rect 319720 548490 319772 548496
rect 319824 547874 319852 555426
rect 319824 547846 319944 547874
rect 319628 547324 319680 547330
rect 319628 547266 319680 547272
rect 319536 545760 319588 545766
rect 319536 545702 319588 545708
rect 319444 543040 319496 543046
rect 319444 542982 319496 542988
rect 319534 542464 319590 542473
rect 319534 542399 319590 542408
rect 319444 541816 319496 541822
rect 319444 541758 319496 541764
rect 318432 540184 318484 540190
rect 318432 540126 318484 540132
rect 318340 519036 318392 519042
rect 318340 518978 318392 518984
rect 318444 518770 318472 540126
rect 319352 540116 319404 540122
rect 319352 540058 319404 540064
rect 319260 523728 319312 523734
rect 319260 523670 319312 523676
rect 318432 518764 318484 518770
rect 318432 518706 318484 518712
rect 319272 518294 319300 523670
rect 319364 518537 319392 540058
rect 319456 518838 319484 541758
rect 319548 519722 319576 542399
rect 319720 541272 319772 541278
rect 319720 541214 319772 541220
rect 319628 541068 319680 541074
rect 319628 541010 319680 541016
rect 319640 523734 319668 541010
rect 319628 523728 319680 523734
rect 319628 523670 319680 523676
rect 319536 519716 319588 519722
rect 319536 519658 319588 519664
rect 319732 518906 319760 541214
rect 319812 540252 319864 540258
rect 319812 540194 319864 540200
rect 319720 518900 319772 518906
rect 319720 518842 319772 518848
rect 319444 518832 319496 518838
rect 319444 518774 319496 518780
rect 319350 518528 319406 518537
rect 319350 518463 319406 518472
rect 319824 518362 319852 540194
rect 319916 518401 319944 547846
rect 427818 520296 427874 520305
rect 320022 520254 320220 520282
rect 356086 520254 356284 520282
rect 320192 519874 320220 520254
rect 324530 520118 324912 520146
rect 320100 519846 320220 519874
rect 320100 518974 320128 519846
rect 324884 518974 324912 520118
rect 328748 520118 329038 520146
rect 333256 520118 333546 520146
rect 337672 520118 338054 520146
rect 342272 520118 342562 520146
rect 346688 520118 347070 520146
rect 351288 520118 351578 520146
rect 320088 518968 320140 518974
rect 320088 518910 320140 518916
rect 324872 518968 324924 518974
rect 324872 518910 324924 518916
rect 328748 518770 328776 520118
rect 333256 518838 333284 520118
rect 333244 518832 333296 518838
rect 333244 518774 333296 518780
rect 328736 518764 328788 518770
rect 328736 518706 328788 518712
rect 337672 518401 337700 520118
rect 319902 518392 319958 518401
rect 319812 518356 319864 518362
rect 319902 518327 319958 518336
rect 337658 518392 337714 518401
rect 337658 518327 337714 518336
rect 319812 518298 319864 518304
rect 319260 518288 319312 518294
rect 319260 518230 319312 518236
rect 342272 518226 342300 520118
rect 346688 518906 346716 520118
rect 351288 519246 351316 520118
rect 351276 519240 351328 519246
rect 351276 519182 351328 519188
rect 346676 518900 346728 518906
rect 346676 518842 346728 518848
rect 356256 518537 356284 520254
rect 427818 520231 427874 520240
rect 360304 520118 360594 520146
rect 364720 520118 365102 520146
rect 369320 520118 369610 520146
rect 374472 520118 374762 520146
rect 378152 520118 379270 520146
rect 383672 520118 383778 520146
rect 387904 520118 388286 520146
rect 391952 520118 392794 520146
rect 396920 520118 397302 520146
rect 401612 520118 401810 520146
rect 406028 520118 406318 520146
rect 410536 520118 410826 520146
rect 414952 520118 415334 520146
rect 419552 520118 419842 520146
rect 423968 520118 424350 520146
rect 356242 518528 356298 518537
rect 356242 518463 356298 518472
rect 360304 518294 360332 520118
rect 364720 518362 364748 520118
rect 369320 519178 369348 520118
rect 369308 519172 369360 519178
rect 369308 519114 369360 519120
rect 374472 518673 374500 520118
rect 374458 518664 374514 518673
rect 374458 518599 374514 518608
rect 364708 518356 364760 518362
rect 364708 518298 364760 518304
rect 360292 518288 360344 518294
rect 360292 518230 360344 518236
rect 342260 518220 342312 518226
rect 342260 518162 342312 518168
rect 318248 517404 318300 517410
rect 318248 517346 318300 517352
rect 317052 517268 317104 517274
rect 317052 517210 317104 517216
rect 316960 515704 317012 515710
rect 316960 515646 317012 515652
rect 316868 514684 316920 514690
rect 316868 514626 316920 514632
rect 302974 502480 303030 502489
rect 302974 502415 303030 502424
rect 302882 487520 302938 487529
rect 302882 487455 302938 487464
rect 302896 487218 302924 487455
rect 302884 487212 302936 487218
rect 302884 487154 302936 487160
rect 59740 480134 60214 480162
rect 299782 480134 299888 480162
rect 59740 480094 59768 480134
rect 59648 480066 59768 480094
rect 189080 480072 189132 480078
rect 50804 479188 50856 479194
rect 50804 479130 50856 479136
rect 50344 479052 50396 479058
rect 50344 478994 50396 479000
rect 45376 478916 45428 478922
rect 45376 478858 45428 478864
rect 43996 473136 44048 473142
rect 43996 473078 44048 473084
rect 42340 472728 42392 472734
rect 42340 472670 42392 472676
rect 43902 472696 43958 472705
rect 42248 470076 42300 470082
rect 42248 470018 42300 470024
rect 41328 382220 41380 382226
rect 41328 382162 41380 382168
rect 42260 373046 42288 470018
rect 42352 373726 42380 472670
rect 43260 472660 43312 472666
rect 43902 472631 43958 472640
rect 43260 472602 43312 472608
rect 42614 472560 42670 472569
rect 42614 472495 42670 472504
rect 42524 470008 42576 470014
rect 42524 469950 42576 469956
rect 42432 466200 42484 466206
rect 42432 466142 42484 466148
rect 42340 373720 42392 373726
rect 42340 373662 42392 373668
rect 42248 373040 42300 373046
rect 42248 372982 42300 372988
rect 42444 267714 42472 466142
rect 42536 269074 42564 469950
rect 42524 269068 42576 269074
rect 42524 269010 42576 269016
rect 42628 268734 42656 472495
rect 42708 470348 42760 470354
rect 42708 470290 42760 470296
rect 42616 268728 42668 268734
rect 42616 268670 42668 268676
rect 42432 267708 42484 267714
rect 42432 267650 42484 267656
rect 42720 248402 42748 470290
rect 43272 373454 43300 472602
rect 43628 470552 43680 470558
rect 43628 470494 43680 470500
rect 43536 470212 43588 470218
rect 43536 470154 43588 470160
rect 43442 469840 43498 469849
rect 43442 469775 43498 469784
rect 43352 460216 43404 460222
rect 43352 460158 43404 460164
rect 43260 373448 43312 373454
rect 43260 373390 43312 373396
rect 43364 269482 43392 460158
rect 43352 269476 43404 269482
rect 43352 269418 43404 269424
rect 43456 268462 43484 469775
rect 43444 268456 43496 268462
rect 43444 268398 43496 268404
rect 43548 267073 43576 470154
rect 43534 267064 43590 267073
rect 43534 266999 43590 267008
rect 43640 264246 43668 470494
rect 43812 470484 43864 470490
rect 43812 470426 43864 470432
rect 43720 470144 43772 470150
rect 43720 470086 43772 470092
rect 43732 264314 43760 470086
rect 43824 264722 43852 470426
rect 43812 264716 43864 264722
rect 43812 264658 43864 264664
rect 43916 264450 43944 472631
rect 44008 264790 44036 473078
rect 45192 470280 45244 470286
rect 45192 470222 45244 470228
rect 44732 469872 44784 469878
rect 44732 469814 44784 469820
rect 44088 468920 44140 468926
rect 44088 468862 44140 468868
rect 43996 264784 44048 264790
rect 43996 264726 44048 264732
rect 43904 264444 43956 264450
rect 43904 264386 43956 264392
rect 43720 264308 43772 264314
rect 43720 264250 43772 264256
rect 43628 264240 43680 264246
rect 43628 264182 43680 264188
rect 42708 248396 42760 248402
rect 42708 248338 42760 248344
rect 41236 57792 41288 57798
rect 41236 57734 41288 57740
rect 41144 57724 41196 57730
rect 41144 57666 41196 57672
rect 44100 55214 44128 468862
rect 44640 409896 44692 409902
rect 44640 409838 44692 409844
rect 44652 373998 44680 409838
rect 44744 385014 44772 469814
rect 45100 468988 45152 468994
rect 45100 468930 45152 468936
rect 45008 468716 45060 468722
rect 45008 468658 45060 468664
rect 44916 468648 44968 468654
rect 44916 468590 44968 468596
rect 44824 466404 44876 466410
rect 44824 466346 44876 466352
rect 44732 385008 44784 385014
rect 44732 384950 44784 384956
rect 44640 373992 44692 373998
rect 44640 373934 44692 373940
rect 44836 269346 44864 466346
rect 44824 269340 44876 269346
rect 44824 269282 44876 269288
rect 44928 269142 44956 468590
rect 45020 269278 45048 468658
rect 45008 269272 45060 269278
rect 45008 269214 45060 269220
rect 45112 269210 45140 468930
rect 45100 269204 45152 269210
rect 45100 269146 45152 269152
rect 44916 269136 44968 269142
rect 44916 269078 44968 269084
rect 45204 268598 45232 470222
rect 45282 469976 45338 469985
rect 45282 469911 45338 469920
rect 45192 268592 45244 268598
rect 45192 268534 45244 268540
rect 45296 264382 45324 469911
rect 45388 269414 45416 478858
rect 50066 478408 50122 478417
rect 48044 478372 48096 478378
rect 50066 478343 50122 478352
rect 48044 478314 48096 478320
rect 47952 478236 48004 478242
rect 47952 478178 48004 478184
rect 45468 476944 45520 476950
rect 45468 476886 45520 476892
rect 45376 269408 45428 269414
rect 45376 269350 45428 269356
rect 45480 264858 45508 476886
rect 47768 476060 47820 476066
rect 47768 476002 47820 476008
rect 46664 475992 46716 475998
rect 46664 475934 46716 475940
rect 46388 475856 46440 475862
rect 46388 475798 46440 475804
rect 46112 472796 46164 472802
rect 46112 472738 46164 472744
rect 46020 408536 46072 408542
rect 46020 408478 46072 408484
rect 46032 375057 46060 408478
rect 46124 383654 46152 472738
rect 46296 465588 46348 465594
rect 46296 465530 46348 465536
rect 46204 462800 46256 462806
rect 46204 462742 46256 462748
rect 46112 383648 46164 383654
rect 46112 383590 46164 383596
rect 46018 375048 46074 375057
rect 46018 374983 46074 374992
rect 46216 371958 46244 462742
rect 46204 371952 46256 371958
rect 46204 371894 46256 371900
rect 46216 364334 46244 371894
rect 46308 371482 46336 465530
rect 46296 371476 46348 371482
rect 46296 371418 46348 371424
rect 46216 364306 46336 364334
rect 46308 287054 46336 364306
rect 46400 299470 46428 475798
rect 46480 475788 46532 475794
rect 46480 475730 46532 475736
rect 46388 299464 46440 299470
rect 46388 299406 46440 299412
rect 46492 298110 46520 475730
rect 46572 468852 46624 468858
rect 46572 468794 46624 468800
rect 46480 298104 46532 298110
rect 46480 298046 46532 298052
rect 46308 287026 46520 287054
rect 46492 267617 46520 287026
rect 46478 267608 46534 267617
rect 46478 267543 46534 267552
rect 45468 264852 45520 264858
rect 45468 264794 45520 264800
rect 45284 264376 45336 264382
rect 45284 264318 45336 264324
rect 46492 148510 46520 267543
rect 46584 264586 46612 468794
rect 46676 268326 46704 475934
rect 46754 475552 46810 475561
rect 46754 475487 46810 475496
rect 46664 268320 46716 268326
rect 46664 268262 46716 268268
rect 46572 264580 46624 264586
rect 46572 264522 46624 264528
rect 46480 148504 46532 148510
rect 46480 148446 46532 148452
rect 46676 145382 46704 268262
rect 46768 267374 46796 475487
rect 46848 473340 46900 473346
rect 46848 473282 46900 473288
rect 46756 267368 46808 267374
rect 46756 267310 46808 267316
rect 46860 264654 46888 473282
rect 47584 472864 47636 472870
rect 47584 472806 47636 472812
rect 47492 465520 47544 465526
rect 47492 465462 47544 465468
rect 47400 460488 47452 460494
rect 47400 460430 47452 460436
rect 47412 372026 47440 460430
rect 47400 372020 47452 372026
rect 47400 371962 47452 371968
rect 47412 371278 47440 371962
rect 47504 371890 47532 465462
rect 47596 373182 47624 472806
rect 47676 472592 47728 472598
rect 47676 472534 47728 472540
rect 47584 373176 47636 373182
rect 47584 373118 47636 373124
rect 47492 371884 47544 371890
rect 47492 371826 47544 371832
rect 47400 371272 47452 371278
rect 47400 371214 47452 371220
rect 47412 268598 47440 268629
rect 47400 268592 47452 268598
rect 47398 268560 47400 268569
rect 47452 268560 47454 268569
rect 47398 268495 47454 268504
rect 47320 268462 47348 268493
rect 47308 268456 47360 268462
rect 47306 268424 47308 268433
rect 47360 268424 47362 268433
rect 47306 268359 47362 268368
rect 47216 268252 47268 268258
rect 47216 268194 47268 268200
rect 46848 264648 46900 264654
rect 46848 264590 46900 264596
rect 47228 145450 47256 268194
rect 47320 160886 47348 268359
rect 47412 160954 47440 268495
rect 47504 267102 47532 371826
rect 47584 371272 47636 371278
rect 47584 371214 47636 371220
rect 47492 267096 47544 267102
rect 47492 267038 47544 267044
rect 47596 266830 47624 371214
rect 47688 267646 47716 472534
rect 47780 268666 47808 476002
rect 47860 475584 47912 475590
rect 47860 475526 47912 475532
rect 47768 268660 47820 268666
rect 47768 268602 47820 268608
rect 47780 268258 47808 268602
rect 47768 268252 47820 268258
rect 47768 268194 47820 268200
rect 47676 267640 47728 267646
rect 47676 267582 47728 267588
rect 47872 267209 47900 475526
rect 47964 268598 47992 478178
rect 47952 268592 48004 268598
rect 47952 268534 48004 268540
rect 48056 268530 48084 478314
rect 49514 478136 49570 478145
rect 49514 478071 49570 478080
rect 49240 475924 49292 475930
rect 49240 475866 49292 475872
rect 48136 475652 48188 475658
rect 48136 475594 48188 475600
rect 48044 268524 48096 268530
rect 48044 268466 48096 268472
rect 47858 267200 47914 267209
rect 47858 267135 47914 267144
rect 47768 267096 47820 267102
rect 47768 267038 47820 267044
rect 47780 266898 47808 267038
rect 47768 266892 47820 266898
rect 47768 266834 47820 266840
rect 47584 266824 47636 266830
rect 47584 266766 47636 266772
rect 47492 264376 47544 264382
rect 47492 264318 47544 264324
rect 47400 160948 47452 160954
rect 47400 160890 47452 160896
rect 47308 160880 47360 160886
rect 47308 160822 47360 160828
rect 47504 160750 47532 264318
rect 47492 160744 47544 160750
rect 47492 160686 47544 160692
rect 47596 145790 47624 266766
rect 47780 148578 47808 266834
rect 48148 264926 48176 475594
rect 49148 475312 49200 475318
rect 49148 475254 49200 475260
rect 49056 473068 49108 473074
rect 49056 473010 49108 473016
rect 48964 469940 49016 469946
rect 48964 469882 49016 469888
rect 48228 466132 48280 466138
rect 48228 466074 48280 466080
rect 48136 264920 48188 264926
rect 48136 264862 48188 264868
rect 47952 264444 48004 264450
rect 47952 264386 48004 264392
rect 47860 264240 47912 264246
rect 47860 264182 47912 264188
rect 47768 148572 47820 148578
rect 47768 148514 47820 148520
rect 47584 145784 47636 145790
rect 47584 145726 47636 145732
rect 47216 145444 47268 145450
rect 47216 145386 47268 145392
rect 46664 145376 46716 145382
rect 46664 145318 46716 145324
rect 47872 144809 47900 264182
rect 47858 144800 47914 144809
rect 47858 144735 47914 144744
rect 47964 144702 47992 264386
rect 48240 162178 48268 466074
rect 48872 463548 48924 463554
rect 48872 463490 48924 463496
rect 48688 460896 48740 460902
rect 48688 460838 48740 460844
rect 48700 459649 48728 460838
rect 48686 459640 48742 459649
rect 48686 459575 48742 459584
rect 48780 458312 48832 458318
rect 48780 458254 48832 458260
rect 48792 451274 48820 458254
rect 48884 456142 48912 463490
rect 48872 456136 48924 456142
rect 48872 456078 48924 456084
rect 48792 451246 48912 451274
rect 48884 412622 48912 451246
rect 48872 412616 48924 412622
rect 48872 412558 48924 412564
rect 48872 407176 48924 407182
rect 48872 407118 48924 407124
rect 48780 405748 48832 405754
rect 48780 405690 48832 405696
rect 48792 373930 48820 405690
rect 48884 375086 48912 407118
rect 48872 375080 48924 375086
rect 48872 375022 48924 375028
rect 48780 373924 48832 373930
rect 48780 373866 48832 373872
rect 48976 373522 49004 469882
rect 48964 373516 49016 373522
rect 48964 373458 49016 373464
rect 49068 373250 49096 473010
rect 49056 373244 49108 373250
rect 49056 373186 49108 373192
rect 49056 371476 49108 371482
rect 49056 371418 49108 371424
rect 49068 267481 49096 371418
rect 49160 268462 49188 475254
rect 49252 268802 49280 475866
rect 49424 466064 49476 466070
rect 49424 466006 49476 466012
rect 49332 456136 49384 456142
rect 49332 456078 49384 456084
rect 49240 268796 49292 268802
rect 49240 268738 49292 268744
rect 49148 268456 49200 268462
rect 49148 268398 49200 268404
rect 49054 267472 49110 267481
rect 49054 267407 49110 267416
rect 48228 162172 48280 162178
rect 48228 162114 48280 162120
rect 49068 148646 49096 267407
rect 49148 264308 49200 264314
rect 49148 264250 49200 264256
rect 49056 148640 49108 148646
rect 49056 148582 49108 148588
rect 49160 145314 49188 264250
rect 49252 145722 49280 268738
rect 49344 162110 49372 456078
rect 49436 164082 49464 466006
rect 49424 164076 49476 164082
rect 49424 164018 49476 164024
rect 49528 162625 49556 478071
rect 49608 460420 49660 460426
rect 49608 460362 49660 460368
rect 49514 162616 49570 162625
rect 49514 162551 49570 162560
rect 49332 162104 49384 162110
rect 49332 162046 49384 162052
rect 49240 145716 49292 145722
rect 49240 145658 49292 145664
rect 49148 145308 49200 145314
rect 49148 145250 49200 145256
rect 47952 144696 48004 144702
rect 47952 144638 48004 144644
rect 49620 59498 49648 460362
rect 49608 59492 49660 59498
rect 49608 59434 49660 59440
rect 50080 58750 50108 478343
rect 50252 475720 50304 475726
rect 50252 475662 50304 475668
rect 50160 473000 50212 473006
rect 50160 472942 50212 472948
rect 50172 373386 50200 472942
rect 50160 373380 50212 373386
rect 50160 373322 50212 373328
rect 50264 265878 50292 475662
rect 50356 267034 50384 478994
rect 50712 478644 50764 478650
rect 50712 478586 50764 478592
rect 50724 477737 50752 478586
rect 50710 477728 50766 477737
rect 50710 477663 50766 477672
rect 50434 475688 50490 475697
rect 50434 475623 50490 475632
rect 50344 267028 50396 267034
rect 50344 266970 50396 266976
rect 50344 266348 50396 266354
rect 50344 266290 50396 266296
rect 50252 265872 50304 265878
rect 50252 265814 50304 265820
rect 50356 144634 50384 266290
rect 50448 249762 50476 475623
rect 50528 466268 50580 466274
rect 50528 466210 50580 466216
rect 50436 249756 50488 249762
rect 50436 249698 50488 249704
rect 50540 164422 50568 466210
rect 50710 465896 50766 465905
rect 50710 465831 50766 465840
rect 50618 462904 50674 462913
rect 50618 462839 50674 462848
rect 50528 164416 50580 164422
rect 50528 164358 50580 164364
rect 50632 161945 50660 462839
rect 50724 163810 50752 465831
rect 50816 163946 50844 479130
rect 52000 479120 52052 479126
rect 52000 479062 52052 479068
rect 51724 478984 51776 478990
rect 51724 478926 51776 478932
rect 50896 477964 50948 477970
rect 50896 477906 50948 477912
rect 50908 477601 50936 477906
rect 50894 477592 50950 477601
rect 50894 477527 50950 477536
rect 50894 463312 50950 463321
rect 50894 463247 50950 463256
rect 50804 163940 50856 163946
rect 50804 163882 50856 163888
rect 50712 163804 50764 163810
rect 50712 163746 50764 163752
rect 50618 161936 50674 161945
rect 50618 161871 50674 161880
rect 50344 144628 50396 144634
rect 50344 144570 50396 144576
rect 50908 59430 50936 463247
rect 51632 460760 51684 460766
rect 51632 460702 51684 460708
rect 51540 460556 51592 460562
rect 51540 460498 51592 460504
rect 51446 383616 51502 383625
rect 51446 383551 51502 383560
rect 51356 267368 51408 267374
rect 51354 267336 51356 267345
rect 51408 267336 51410 267345
rect 51354 267271 51410 267280
rect 50896 59424 50948 59430
rect 50896 59366 50948 59372
rect 50068 58744 50120 58750
rect 50068 58686 50120 58692
rect 51460 57866 51488 383551
rect 51448 57860 51500 57866
rect 51448 57802 51500 57808
rect 51552 57390 51580 460498
rect 51644 459649 51672 460702
rect 51630 459640 51686 459649
rect 51630 459575 51686 459584
rect 51632 459196 51684 459202
rect 51632 459138 51684 459144
rect 51644 405006 51672 459138
rect 51632 405000 51684 405006
rect 51632 404942 51684 404948
rect 51632 404388 51684 404394
rect 51632 404330 51684 404336
rect 51644 375018 51672 404330
rect 51736 383586 51764 478926
rect 51908 478304 51960 478310
rect 51908 478246 51960 478252
rect 51816 475244 51868 475250
rect 51816 475186 51868 475192
rect 51724 383580 51776 383586
rect 51724 383522 51776 383528
rect 51632 375012 51684 375018
rect 51632 374954 51684 374960
rect 51828 268394 51856 475186
rect 51816 268388 51868 268394
rect 51816 268330 51868 268336
rect 51920 267170 51948 478246
rect 51908 267164 51960 267170
rect 51908 267106 51960 267112
rect 52012 267102 52040 479062
rect 53748 478848 53800 478854
rect 53748 478790 53800 478796
rect 52184 478712 52236 478718
rect 52184 478654 52236 478660
rect 52092 466336 52144 466342
rect 52092 466278 52144 466284
rect 52000 267096 52052 267102
rect 52000 267038 52052 267044
rect 52000 265872 52052 265878
rect 52000 265814 52052 265820
rect 51908 148504 51960 148510
rect 51908 148446 51960 148452
rect 51540 57384 51592 57390
rect 51540 57326 51592 57332
rect 51920 55758 51948 148446
rect 52012 144770 52040 265814
rect 52104 164014 52132 466278
rect 52092 164008 52144 164014
rect 52092 163950 52144 163956
rect 52196 163878 52224 478654
rect 52276 472932 52328 472938
rect 52276 472874 52328 472880
rect 52288 373590 52316 472874
rect 53656 469804 53708 469810
rect 53656 469746 53708 469752
rect 53562 466168 53618 466177
rect 53562 466103 53618 466112
rect 53196 465860 53248 465866
rect 53196 465802 53248 465808
rect 53104 465724 53156 465730
rect 53104 465666 53156 465672
rect 52920 463344 52972 463350
rect 52920 463286 52972 463292
rect 52368 460692 52420 460698
rect 52368 460634 52420 460640
rect 52380 459649 52408 460634
rect 52366 459640 52422 459649
rect 52366 459575 52422 459584
rect 52932 456142 52960 463286
rect 53012 459128 53064 459134
rect 53012 459070 53064 459076
rect 52920 456136 52972 456142
rect 52920 456078 52972 456084
rect 52368 403028 52420 403034
rect 52368 402970 52420 402976
rect 52380 374921 52408 402970
rect 52920 383580 52972 383586
rect 52920 383522 52972 383528
rect 52826 375320 52882 375329
rect 52826 375255 52882 375264
rect 52366 374912 52422 374921
rect 52366 374847 52422 374856
rect 52276 373584 52328 373590
rect 52276 373526 52328 373532
rect 52366 267336 52422 267345
rect 52366 267271 52422 267280
rect 52184 163872 52236 163878
rect 52184 163814 52236 163820
rect 52092 160880 52144 160886
rect 52092 160822 52144 160828
rect 52000 144764 52052 144770
rect 52000 144706 52052 144712
rect 52104 57458 52132 160822
rect 52380 160818 52408 267271
rect 52552 265736 52604 265742
rect 52552 265678 52604 265684
rect 52564 264722 52592 265678
rect 52736 265668 52788 265674
rect 52736 265610 52788 265616
rect 52748 264897 52776 265610
rect 52734 264888 52790 264897
rect 52734 264823 52790 264832
rect 52552 264716 52604 264722
rect 52552 264658 52604 264664
rect 52736 249756 52788 249762
rect 52736 249698 52788 249704
rect 52748 249150 52776 249698
rect 52736 249144 52788 249150
rect 52736 249086 52788 249092
rect 52748 243710 52776 249086
rect 52736 243704 52788 243710
rect 52736 243646 52788 243652
rect 52840 243642 52868 375255
rect 52932 269550 52960 383522
rect 52920 269544 52972 269550
rect 52920 269486 52972 269492
rect 53024 267374 53052 459070
rect 53012 267368 53064 267374
rect 53012 267310 53064 267316
rect 53116 267238 53144 465666
rect 53208 267306 53236 465802
rect 53288 463072 53340 463078
rect 53288 463014 53340 463020
rect 53300 458402 53328 463014
rect 53380 463004 53432 463010
rect 53380 462946 53432 462952
rect 53392 460934 53420 462946
rect 53392 460906 53512 460934
rect 53380 460828 53432 460834
rect 53380 460770 53432 460776
rect 53392 459649 53420 460770
rect 53378 459640 53434 459649
rect 53378 459575 53434 459584
rect 53300 458374 53420 458402
rect 53288 456136 53340 456142
rect 53288 456078 53340 456084
rect 53196 267300 53248 267306
rect 53196 267242 53248 267248
rect 53104 267232 53156 267238
rect 53104 267174 53156 267180
rect 53194 264888 53250 264897
rect 53194 264823 53250 264832
rect 53104 264716 53156 264722
rect 53104 264658 53156 264664
rect 53012 249076 53064 249082
rect 53012 249018 53064 249024
rect 53024 248414 53052 249018
rect 52932 248402 53052 248414
rect 52920 248396 53052 248402
rect 52972 248386 53052 248396
rect 52920 248338 52972 248344
rect 52828 243636 52880 243642
rect 52828 243578 52880 243584
rect 52828 243432 52880 243438
rect 52828 243374 52880 243380
rect 52368 160812 52420 160818
rect 52368 160754 52420 160760
rect 52184 160744 52236 160750
rect 52184 160686 52236 160692
rect 52092 57452 52144 57458
rect 52092 57394 52144 57400
rect 51908 55752 51960 55758
rect 51908 55694 51960 55700
rect 44088 55208 44140 55214
rect 44088 55150 44140 55156
rect 52196 55078 52224 160686
rect 52368 145784 52420 145790
rect 52368 145726 52420 145732
rect 52380 57254 52408 145726
rect 52840 58682 52868 243374
rect 52932 162926 52960 248338
rect 53012 243704 53064 243710
rect 53012 243646 53064 243652
rect 52920 162920 52972 162926
rect 52920 162862 52972 162868
rect 53024 161090 53052 243646
rect 53012 161084 53064 161090
rect 53012 161026 53064 161032
rect 53012 149048 53064 149054
rect 53012 148990 53064 148996
rect 53024 58818 53052 148990
rect 53116 144838 53144 264658
rect 53208 149054 53236 264823
rect 53300 162450 53328 456078
rect 53392 162518 53420 458374
rect 53380 162512 53432 162518
rect 53484 162489 53512 460906
rect 53380 162454 53432 162460
rect 53470 162480 53526 162489
rect 53288 162444 53340 162450
rect 53470 162415 53526 162424
rect 53288 162386 53340 162392
rect 53576 162246 53604 466103
rect 53668 374678 53696 469746
rect 53656 374672 53708 374678
rect 53656 374614 53708 374620
rect 53564 162240 53616 162246
rect 53564 162182 53616 162188
rect 53472 160948 53524 160954
rect 53472 160890 53524 160896
rect 53196 149048 53248 149054
rect 53196 148990 53248 148996
rect 53380 148572 53432 148578
rect 53380 148514 53432 148520
rect 53288 148368 53340 148374
rect 53288 148310 53340 148316
rect 53196 146056 53248 146062
rect 53196 145998 53248 146004
rect 53104 144832 53156 144838
rect 53104 144774 53156 144780
rect 53012 58812 53064 58818
rect 53012 58754 53064 58760
rect 52828 58676 52880 58682
rect 52828 58618 52880 58624
rect 52368 57248 52420 57254
rect 52368 57190 52420 57196
rect 52184 55072 52236 55078
rect 52184 55014 52236 55020
rect 53208 54874 53236 145998
rect 53300 55146 53328 148310
rect 53288 55140 53340 55146
rect 53288 55082 53340 55088
rect 53196 54868 53248 54874
rect 53196 54810 53248 54816
rect 53392 54738 53420 148514
rect 53484 56506 53512 160890
rect 53564 160132 53616 160138
rect 53564 160074 53616 160080
rect 53472 56500 53524 56506
rect 53472 56442 53524 56448
rect 53576 55826 53604 160074
rect 53760 57662 53788 478790
rect 54760 478440 54812 478446
rect 54760 478382 54812 478388
rect 54668 475176 54720 475182
rect 54668 475118 54720 475124
rect 54576 472524 54628 472530
rect 54576 472466 54628 472472
rect 54484 460148 54536 460154
rect 54484 460090 54536 460096
rect 54392 458992 54444 458998
rect 54392 458934 54444 458940
rect 54300 458856 54352 458862
rect 54300 458798 54352 458804
rect 54312 374066 54340 458798
rect 54404 374882 54432 458934
rect 54392 374876 54444 374882
rect 54392 374818 54444 374824
rect 54300 374060 54352 374066
rect 54300 374002 54352 374008
rect 54496 371142 54524 460090
rect 54484 371136 54536 371142
rect 54484 371078 54536 371084
rect 54484 303816 54536 303822
rect 54484 303758 54536 303764
rect 53840 268116 53892 268122
rect 53840 268058 53892 268064
rect 53852 267646 53880 268058
rect 54496 267782 54524 303758
rect 54484 267776 54536 267782
rect 54312 267724 54484 267734
rect 54312 267718 54536 267724
rect 54312 267706 54524 267718
rect 53840 267640 53892 267646
rect 53840 267582 53892 267588
rect 53852 146062 53880 267582
rect 54116 266212 54168 266218
rect 54116 266154 54168 266160
rect 53932 266076 53984 266082
rect 53932 266018 53984 266024
rect 53944 264654 53972 266018
rect 54128 264926 54156 266154
rect 54116 264920 54168 264926
rect 54116 264862 54168 264868
rect 53932 264648 53984 264654
rect 53932 264590 53984 264596
rect 54208 146260 54260 146266
rect 54208 146202 54260 146208
rect 53840 146056 53892 146062
rect 53840 145998 53892 146004
rect 54220 59566 54248 146202
rect 54312 145761 54340 267706
rect 54588 265946 54616 472466
rect 54680 266966 54708 475118
rect 54772 267442 54800 478382
rect 55128 478168 55180 478174
rect 55128 478110 55180 478116
rect 55036 463616 55088 463622
rect 55036 463558 55088 463564
rect 54852 463208 54904 463214
rect 54852 463150 54904 463156
rect 54760 267436 54812 267442
rect 54760 267378 54812 267384
rect 54668 266960 54720 266966
rect 54668 266902 54720 266908
rect 54576 265940 54628 265946
rect 54576 265882 54628 265888
rect 54484 264920 54536 264926
rect 54484 264862 54536 264868
rect 54392 162920 54444 162926
rect 54392 162862 54444 162868
rect 54298 145752 54354 145761
rect 54298 145687 54354 145696
rect 54208 59560 54260 59566
rect 54208 59502 54260 59508
rect 54404 58954 54432 162862
rect 54496 144906 54524 264862
rect 54576 264648 54628 264654
rect 54576 264590 54628 264596
rect 54588 145926 54616 264590
rect 54668 249212 54720 249218
rect 54668 249154 54720 249160
rect 54680 161362 54708 249154
rect 54864 162722 54892 463150
rect 54944 462936 54996 462942
rect 54944 462878 54996 462884
rect 54852 162716 54904 162722
rect 54852 162658 54904 162664
rect 54956 162314 54984 462878
rect 55048 162586 55076 463558
rect 55140 162858 55168 478110
rect 56508 478032 56560 478038
rect 56508 477974 56560 477980
rect 56048 470416 56100 470422
rect 56048 470358 56100 470364
rect 55864 463684 55916 463690
rect 55864 463626 55916 463632
rect 55772 459264 55824 459270
rect 55772 459206 55824 459212
rect 55680 408604 55732 408610
rect 55680 408546 55732 408552
rect 55692 371385 55720 408546
rect 55784 375358 55812 459206
rect 55876 457298 55904 463626
rect 55956 460624 56008 460630
rect 55956 460566 56008 460572
rect 55968 459649 55996 460566
rect 55954 459640 56010 459649
rect 55954 459575 56010 459584
rect 55956 458924 56008 458930
rect 55956 458866 56008 458872
rect 55864 457292 55916 457298
rect 55864 457234 55916 457240
rect 55864 405000 55916 405006
rect 55864 404942 55916 404948
rect 55772 375352 55824 375358
rect 55772 375294 55824 375300
rect 55678 371376 55734 371385
rect 55678 371311 55734 371320
rect 55876 269618 55904 404942
rect 55968 373114 55996 458866
rect 56060 380866 56088 470358
rect 56232 463480 56284 463486
rect 56232 463422 56284 463428
rect 56140 463412 56192 463418
rect 56140 463354 56192 463360
rect 56048 380860 56100 380866
rect 56048 380802 56100 380808
rect 55956 373108 56008 373114
rect 55956 373050 56008 373056
rect 56048 353388 56100 353394
rect 56048 353330 56100 353336
rect 55956 351960 56008 351966
rect 55956 351902 56008 351908
rect 55864 269612 55916 269618
rect 55864 269554 55916 269560
rect 55968 267646 55996 351902
rect 55956 267640 56008 267646
rect 55956 267582 56008 267588
rect 56060 267510 56088 353330
rect 56048 267504 56100 267510
rect 56048 267446 56100 267452
rect 56048 265940 56100 265946
rect 56048 265882 56100 265888
rect 55956 249416 56008 249422
rect 55956 249358 56008 249364
rect 55128 162852 55180 162858
rect 55128 162794 55180 162800
rect 55126 162752 55182 162761
rect 55126 162687 55182 162696
rect 55036 162580 55088 162586
rect 55036 162522 55088 162528
rect 54944 162308 54996 162314
rect 54944 162250 54996 162256
rect 54668 161356 54720 161362
rect 54668 161298 54720 161304
rect 54680 160138 54708 161298
rect 54668 160132 54720 160138
rect 54668 160074 54720 160080
rect 54944 148640 54996 148646
rect 54944 148582 54996 148588
rect 54576 145920 54628 145926
rect 54576 145862 54628 145868
rect 54852 145920 54904 145926
rect 54852 145862 54904 145868
rect 54668 145716 54720 145722
rect 54668 145658 54720 145664
rect 54484 144900 54536 144906
rect 54484 144842 54536 144848
rect 54680 59634 54708 145658
rect 54760 145376 54812 145382
rect 54760 145318 54812 145324
rect 54668 59628 54720 59634
rect 54668 59570 54720 59576
rect 54392 58948 54444 58954
rect 54392 58890 54444 58896
rect 53748 57656 53800 57662
rect 53748 57598 53800 57604
rect 54772 57186 54800 145318
rect 54760 57180 54812 57186
rect 54760 57122 54812 57128
rect 54864 55962 54892 145862
rect 54956 56574 54984 148582
rect 55036 145444 55088 145450
rect 55036 145386 55088 145392
rect 55048 59702 55076 145386
rect 55036 59696 55088 59702
rect 55036 59638 55088 59644
rect 55140 57526 55168 162687
rect 55968 161430 55996 249358
rect 56060 161474 56088 265882
rect 56152 162654 56180 463354
rect 56244 162790 56272 463422
rect 56416 463276 56468 463282
rect 56416 463218 56468 463224
rect 56428 460934 56456 463218
rect 56336 460906 56456 460934
rect 56232 162784 56284 162790
rect 56232 162726 56284 162732
rect 56140 162648 56192 162654
rect 56140 162590 56192 162596
rect 56336 162353 56364 460906
rect 56416 457292 56468 457298
rect 56416 457234 56468 457240
rect 56428 162382 56456 457234
rect 56416 162376 56468 162382
rect 56322 162344 56378 162353
rect 56416 162318 56468 162324
rect 56322 162279 56378 162288
rect 56520 162042 56548 477974
rect 58440 477896 58492 477902
rect 58440 477838 58492 477844
rect 57152 475516 57204 475522
rect 57152 475458 57204 475464
rect 57060 469736 57112 469742
rect 57060 469678 57112 469684
rect 56968 412616 57020 412622
rect 56968 412558 57020 412564
rect 56980 412321 57008 412558
rect 56966 412312 57022 412321
rect 56966 412247 57022 412256
rect 57072 410530 57100 469678
rect 56980 410502 57100 410530
rect 56980 408610 57008 410502
rect 57058 410408 57114 410417
rect 57058 410343 57114 410352
rect 57072 409902 57100 410343
rect 57060 409896 57112 409902
rect 57060 409838 57112 409844
rect 57058 408640 57114 408649
rect 56968 408604 57020 408610
rect 57058 408575 57114 408584
rect 56968 408546 57020 408552
rect 57072 408542 57100 408575
rect 57060 408536 57112 408542
rect 57060 408478 57112 408484
rect 56966 407416 57022 407425
rect 56966 407351 57022 407360
rect 56980 407182 57008 407351
rect 56968 407176 57020 407182
rect 56968 407118 57020 407124
rect 57058 405784 57114 405793
rect 57058 405719 57060 405728
rect 57112 405719 57114 405728
rect 57060 405690 57112 405696
rect 57058 404424 57114 404433
rect 57058 404359 57060 404368
rect 57112 404359 57114 404368
rect 57060 404330 57112 404336
rect 57058 403064 57114 403073
rect 57058 402999 57060 403008
rect 57112 402999 57114 403008
rect 57060 402970 57112 402976
rect 57164 389174 57192 475458
rect 57336 475448 57388 475454
rect 57336 475390 57388 475396
rect 57244 465928 57296 465934
rect 57244 465870 57296 465876
rect 56980 389146 57192 389174
rect 56600 385008 56652 385014
rect 56598 384976 56600 384985
rect 56652 384976 56654 384985
rect 56598 384911 56654 384920
rect 56600 383648 56652 383654
rect 56600 383590 56652 383596
rect 56612 383081 56640 383590
rect 56598 383072 56654 383081
rect 56598 383007 56654 383016
rect 56600 374876 56652 374882
rect 56600 374818 56652 374824
rect 56612 303822 56640 374818
rect 56980 374134 57008 389146
rect 57256 384418 57284 465870
rect 57072 384390 57284 384418
rect 57072 383654 57100 384390
rect 57348 384282 57376 475390
rect 57888 472456 57940 472462
rect 57888 472398 57940 472404
rect 57704 471300 57756 471306
rect 57704 471242 57756 471248
rect 57520 467152 57572 467158
rect 57520 467094 57572 467100
rect 57428 463140 57480 463146
rect 57428 463082 57480 463088
rect 57164 384254 57376 384282
rect 57440 384266 57468 463082
rect 57428 384260 57480 384266
rect 57060 383648 57112 383654
rect 57060 383590 57112 383596
rect 57060 380860 57112 380866
rect 57060 380802 57112 380808
rect 56968 374128 57020 374134
rect 56968 374070 57020 374076
rect 57072 373658 57100 380802
rect 57164 378690 57192 384254
rect 57428 384202 57480 384208
rect 57532 384146 57560 467094
rect 57612 464364 57664 464370
rect 57612 464306 57664 464312
rect 57348 384118 57560 384146
rect 57242 383344 57298 383353
rect 57242 383279 57298 383288
rect 57256 382226 57284 383279
rect 57244 382220 57296 382226
rect 57244 382162 57296 382168
rect 57152 378684 57204 378690
rect 57152 378626 57204 378632
rect 57060 373652 57112 373658
rect 57060 373594 57112 373600
rect 57060 352028 57112 352034
rect 57060 351970 57112 351976
rect 56874 305008 56930 305017
rect 56874 304943 56930 304952
rect 56600 303816 56652 303822
rect 56600 303758 56652 303764
rect 56888 201385 56916 304943
rect 56968 299464 57020 299470
rect 56968 299406 57020 299412
rect 56874 201376 56930 201385
rect 56874 201311 56930 201320
rect 56874 198792 56930 198801
rect 56874 198727 56930 198736
rect 56508 162036 56560 162042
rect 56508 161978 56560 161984
rect 56060 161446 56364 161474
rect 55956 161424 56008 161430
rect 55956 161366 56008 161372
rect 55968 160177 55996 161366
rect 55954 160168 56010 160177
rect 55954 160103 56010 160112
rect 56336 151814 56364 161446
rect 56508 161084 56560 161090
rect 56508 161026 56560 161032
rect 56060 151786 56364 151814
rect 56060 145994 56088 151786
rect 56232 148436 56284 148442
rect 56232 148378 56284 148384
rect 56140 147212 56192 147218
rect 56140 147154 56192 147160
rect 56048 145988 56100 145994
rect 56048 145930 56100 145936
rect 55956 144900 56008 144906
rect 55956 144842 56008 144848
rect 55864 144832 55916 144838
rect 55864 144774 55916 144780
rect 55876 59090 55904 144774
rect 55968 59362 55996 144842
rect 56060 144378 56088 145930
rect 56152 144566 56180 147154
rect 56140 144560 56192 144566
rect 56140 144502 56192 144508
rect 56244 144498 56272 148378
rect 56324 145648 56376 145654
rect 56324 145590 56376 145596
rect 56414 145616 56470 145625
rect 56336 144906 56364 145590
rect 56414 145551 56470 145560
rect 56324 144900 56376 144906
rect 56324 144842 56376 144848
rect 56428 144838 56456 145551
rect 56416 144832 56468 144838
rect 56416 144774 56468 144780
rect 56416 144560 56468 144566
rect 56416 144502 56468 144508
rect 56232 144492 56284 144498
rect 56232 144434 56284 144440
rect 56060 144350 56364 144378
rect 56232 144288 56284 144294
rect 56232 144230 56284 144236
rect 55956 59356 56008 59362
rect 55956 59298 56008 59304
rect 55864 59084 55916 59090
rect 55864 59026 55916 59032
rect 56244 58886 56272 144230
rect 56232 58880 56284 58886
rect 56232 58822 56284 58828
rect 55128 57520 55180 57526
rect 55128 57462 55180 57468
rect 54944 56568 54996 56574
rect 54944 56510 54996 56516
rect 56336 56030 56364 144350
rect 56428 56234 56456 144502
rect 56520 59158 56548 161026
rect 56888 93809 56916 198727
rect 56980 195265 57008 299406
rect 57072 267578 57100 351970
rect 57150 307728 57206 307737
rect 57150 307663 57206 307672
rect 57164 306921 57192 307663
rect 57150 306912 57206 306921
rect 57150 306847 57206 306856
rect 57060 267572 57112 267578
rect 57060 267514 57112 267520
rect 57164 209774 57192 306847
rect 57256 278769 57284 382162
rect 57348 378826 57376 384118
rect 57428 384056 57480 384062
rect 57428 383998 57480 384004
rect 57336 378820 57388 378826
rect 57336 378762 57388 378768
rect 57336 378684 57388 378690
rect 57336 378626 57388 378632
rect 57348 373318 57376 378626
rect 57336 373312 57388 373318
rect 57336 373254 57388 373260
rect 57440 306374 57468 383998
rect 57520 378820 57572 378826
rect 57520 378762 57572 378768
rect 57532 307737 57560 378762
rect 57518 307728 57574 307737
rect 57518 307663 57574 307672
rect 57440 306346 57560 306374
rect 57334 303648 57390 303657
rect 57334 303583 57390 303592
rect 57242 278760 57298 278769
rect 57242 278695 57298 278704
rect 57244 264784 57296 264790
rect 57244 264726 57296 264732
rect 57072 209746 57192 209774
rect 57072 201929 57100 209746
rect 57058 201920 57114 201929
rect 57058 201855 57114 201864
rect 56966 195256 57022 195265
rect 56966 195191 57022 195200
rect 56968 146192 57020 146198
rect 56968 146134 57020 146140
rect 56874 93800 56930 93809
rect 56874 93735 56930 93744
rect 56508 59152 56560 59158
rect 56508 59094 56560 59100
rect 56416 56228 56468 56234
rect 56416 56170 56468 56176
rect 56324 56024 56376 56030
rect 56324 55966 56376 55972
rect 54852 55956 54904 55962
rect 54852 55898 54904 55904
rect 53564 55820 53616 55826
rect 53564 55762 53616 55768
rect 56980 54942 57008 146134
rect 57072 97481 57100 201855
rect 57150 201376 57206 201385
rect 57150 201311 57206 201320
rect 57058 97472 57114 97481
rect 57058 97407 57114 97416
rect 57164 96529 57192 201311
rect 57256 146198 57284 264726
rect 57348 198801 57376 303583
rect 57532 302297 57560 306346
rect 57518 302288 57574 302297
rect 57518 302223 57574 302232
rect 57426 299568 57482 299577
rect 57426 299503 57482 299512
rect 57440 299470 57468 299503
rect 57428 299464 57480 299470
rect 57428 299406 57480 299412
rect 57426 298208 57482 298217
rect 57426 298143 57482 298152
rect 57440 298110 57468 298143
rect 57428 298104 57480 298110
rect 57428 298046 57480 298052
rect 57334 198792 57390 198801
rect 57334 198727 57390 198736
rect 57334 197432 57390 197441
rect 57334 197367 57390 197376
rect 57244 146192 57296 146198
rect 57244 146134 57296 146140
rect 57150 96520 57206 96529
rect 57150 96455 57206 96464
rect 57348 93401 57376 197367
rect 57440 193225 57468 298046
rect 57532 197441 57560 302223
rect 57624 301345 57652 464306
rect 57716 303657 57744 471242
rect 57796 459060 57848 459066
rect 57796 459002 57848 459008
rect 57702 303648 57758 303657
rect 57702 303583 57758 303592
rect 57610 301336 57666 301345
rect 57610 301271 57666 301280
rect 57624 209774 57652 301271
rect 57808 277394 57836 459002
rect 57900 305969 57928 472398
rect 57980 383648 58032 383654
rect 58452 383625 58480 477838
rect 58990 475960 59046 475969
rect 58990 475895 59046 475904
rect 58808 474020 58860 474026
rect 58808 473962 58860 473968
rect 58624 473272 58676 473278
rect 58624 473214 58676 473220
rect 58532 469668 58584 469674
rect 58532 469610 58584 469616
rect 57980 383590 58032 383596
rect 58438 383616 58494 383625
rect 57992 351966 58020 383590
rect 58438 383551 58494 383560
rect 58544 372881 58572 469610
rect 58636 374202 58664 473214
rect 58716 465792 58768 465798
rect 58716 465734 58768 465740
rect 58624 374196 58676 374202
rect 58624 374138 58676 374144
rect 58530 372872 58586 372881
rect 58530 372807 58586 372816
rect 58622 372736 58678 372745
rect 58622 372671 58678 372680
rect 58532 353320 58584 353326
rect 58532 353262 58584 353268
rect 57980 351960 58032 351966
rect 57980 351902 58032 351908
rect 57886 305960 57942 305969
rect 57886 305895 57942 305904
rect 57900 305017 57928 305895
rect 57886 305008 57942 305017
rect 57886 304943 57942 304952
rect 57886 278760 57942 278769
rect 57886 278695 57942 278704
rect 57716 277366 57836 277394
rect 57716 266354 57744 277366
rect 57796 268728 57848 268734
rect 57796 268670 57848 268676
rect 57808 267918 57836 268670
rect 57796 267912 57848 267918
rect 57796 267854 57848 267860
rect 57704 266348 57756 266354
rect 57704 266290 57756 266296
rect 57704 265804 57756 265810
rect 57704 265746 57756 265752
rect 57716 264790 57744 265746
rect 57704 264784 57756 264790
rect 57704 264726 57756 264732
rect 57624 209746 57744 209774
rect 57518 197432 57574 197441
rect 57518 197367 57574 197376
rect 57716 196081 57744 209746
rect 57702 196072 57758 196081
rect 57702 196007 57758 196016
rect 57518 195256 57574 195265
rect 57518 195191 57574 195200
rect 57426 193216 57482 193225
rect 57426 193151 57482 193160
rect 57334 93392 57390 93401
rect 57334 93327 57390 93336
rect 57440 88233 57468 193151
rect 57532 90545 57560 195191
rect 57716 91089 57744 196007
rect 57808 147626 57836 267854
rect 57900 173369 57928 278695
rect 58544 276049 58572 353262
rect 58530 276040 58586 276049
rect 58530 275975 58586 275984
rect 58636 268054 58664 372671
rect 58728 279993 58756 465734
rect 58714 279984 58770 279993
rect 58714 279919 58770 279928
rect 58820 278089 58848 473962
rect 58900 459332 58952 459338
rect 58900 459274 58952 459280
rect 58806 278080 58862 278089
rect 58806 278015 58862 278024
rect 58624 268048 58676 268054
rect 58624 267990 58676 267996
rect 58636 267734 58664 267990
rect 58636 267706 58848 267734
rect 58622 267064 58678 267073
rect 58622 266999 58678 267008
rect 58440 249756 58492 249762
rect 58440 249698 58492 249704
rect 58346 175264 58402 175273
rect 58346 175199 58402 175208
rect 57886 173360 57942 173369
rect 57886 173295 57942 173304
rect 57796 147620 57848 147626
rect 57796 147562 57848 147568
rect 57702 91080 57758 91089
rect 57702 91015 57758 91024
rect 57518 90536 57574 90545
rect 57518 90471 57574 90480
rect 57426 88224 57482 88233
rect 57426 88159 57482 88168
rect 57244 57588 57296 57594
rect 57244 57530 57296 57536
rect 56968 54936 57020 54942
rect 56968 54878 57020 54884
rect 53380 54732 53432 54738
rect 53380 54674 53432 54680
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 2792 19417 2820 20334
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 57256 3466 57284 57530
rect 57808 56370 57836 147562
rect 57900 68921 57928 173295
rect 57886 68912 57942 68921
rect 57886 68847 57942 68856
rect 57900 57934 57928 68847
rect 57888 57928 57940 57934
rect 57888 57870 57940 57876
rect 57900 57594 57928 57870
rect 57888 57588 57940 57594
rect 57888 57530 57940 57536
rect 58360 57322 58388 175199
rect 58452 160138 58480 249698
rect 58532 249688 58584 249694
rect 58532 249630 58584 249636
rect 58544 161022 58572 249630
rect 58532 161016 58584 161022
rect 58532 160958 58584 160964
rect 58440 160132 58492 160138
rect 58440 160074 58492 160080
rect 58636 147558 58664 266999
rect 58716 266144 58768 266150
rect 58716 266086 58768 266092
rect 58728 264858 58756 266086
rect 58716 264852 58768 264858
rect 58716 264794 58768 264800
rect 58624 147552 58676 147558
rect 58624 147494 58676 147500
rect 58636 147218 58664 147494
rect 58624 147212 58676 147218
rect 58624 147154 58676 147160
rect 58728 146146 58756 264794
rect 58820 146266 58848 267706
rect 58912 163538 58940 459274
rect 59004 175273 59032 475895
rect 59648 470594 59676 480066
rect 60004 478780 60056 478786
rect 60004 478722 60056 478728
rect 59728 473204 59780 473210
rect 59728 473146 59780 473152
rect 59372 470566 59676 470594
rect 59372 468586 59400 470566
rect 59360 468580 59412 468586
rect 59360 468522 59412 468528
rect 59082 466440 59138 466449
rect 59082 466375 59138 466384
rect 58990 175264 59046 175273
rect 58990 175199 59046 175208
rect 59096 164354 59124 466375
rect 59174 466304 59230 466313
rect 59174 466239 59230 466248
rect 59084 164348 59136 164354
rect 59084 164290 59136 164296
rect 59188 163674 59216 466239
rect 59268 458652 59320 458658
rect 59268 458594 59320 458600
rect 59176 163668 59228 163674
rect 59176 163610 59228 163616
rect 58900 163532 58952 163538
rect 58900 163474 58952 163480
rect 59176 161288 59228 161294
rect 59176 161230 59228 161236
rect 59084 161152 59136 161158
rect 59084 161094 59136 161100
rect 59096 160818 59124 161094
rect 59188 161022 59216 161230
rect 59176 161016 59228 161022
rect 59176 160958 59228 160964
rect 59084 160812 59136 160818
rect 59084 160754 59136 160760
rect 58808 146260 58860 146266
rect 58808 146202 58860 146208
rect 58728 146118 58940 146146
rect 58622 145888 58678 145897
rect 58912 145858 58940 146118
rect 58622 145823 58678 145832
rect 58900 145852 58952 145858
rect 58530 145752 58586 145761
rect 58530 145687 58586 145696
rect 58544 59022 58572 145687
rect 58636 144702 58664 145823
rect 58900 145794 58952 145800
rect 58808 145580 58860 145586
rect 58808 145522 58860 145528
rect 58716 145512 58768 145518
rect 58716 145454 58768 145460
rect 58728 144770 58756 145454
rect 58716 144764 58768 144770
rect 58716 144706 58768 144712
rect 58624 144696 58676 144702
rect 58624 144638 58676 144644
rect 58532 59016 58584 59022
rect 58532 58958 58584 58964
rect 58348 57316 58400 57322
rect 58348 57258 58400 57264
rect 57796 56364 57848 56370
rect 57796 56306 57848 56312
rect 58636 55010 58664 144638
rect 58728 55894 58756 144706
rect 58820 144634 58848 145522
rect 58808 144628 58860 144634
rect 58808 144570 58860 144576
rect 58820 56098 58848 144570
rect 58808 56092 58860 56098
rect 58808 56034 58860 56040
rect 58716 55888 58768 55894
rect 58716 55830 58768 55836
rect 58624 55004 58676 55010
rect 58624 54946 58676 54952
rect 58912 54806 58940 145794
rect 59096 59226 59124 160754
rect 59084 59220 59136 59226
rect 59084 59162 59136 59168
rect 58992 57520 59044 57526
rect 58992 57462 59044 57468
rect 59004 57322 59032 57462
rect 58992 57316 59044 57322
rect 58992 57258 59044 57264
rect 59188 56302 59216 160958
rect 59280 57322 59308 458594
rect 59360 375352 59412 375358
rect 59360 375294 59412 375300
rect 59372 352034 59400 375294
rect 59636 374672 59688 374678
rect 59636 374614 59688 374620
rect 59360 352028 59412 352034
rect 59360 351970 59412 351976
rect 59648 269074 59676 374614
rect 59740 373794 59768 473146
rect 59910 466032 59966 466041
rect 59820 465996 59872 466002
rect 59910 465967 59966 465976
rect 59820 465938 59872 465944
rect 59728 373788 59780 373794
rect 59728 373730 59780 373736
rect 59728 373040 59780 373046
rect 59728 372982 59780 372988
rect 59636 269068 59688 269074
rect 59636 269010 59688 269016
rect 59740 267850 59768 372982
rect 59832 353394 59860 465938
rect 59820 353388 59872 353394
rect 59820 353330 59872 353336
rect 59818 276176 59874 276185
rect 59818 276111 59874 276120
rect 59832 268841 59860 276111
rect 59818 268832 59874 268841
rect 59818 268767 59874 268776
rect 59728 267844 59780 267850
rect 59728 267786 59780 267792
rect 59740 161226 59768 267786
rect 59818 267200 59874 267209
rect 59818 267135 59874 267144
rect 59832 266393 59860 267135
rect 59818 266384 59874 266393
rect 59818 266319 59874 266328
rect 59728 161220 59780 161226
rect 59728 161162 59780 161168
rect 59360 160812 59412 160818
rect 59360 160754 59412 160760
rect 59372 160138 59400 160754
rect 59740 160342 59768 161162
rect 59728 160336 59780 160342
rect 59728 160278 59780 160284
rect 59360 160132 59412 160138
rect 59360 160074 59412 160080
rect 59372 140865 59400 160074
rect 59832 146198 59860 266319
rect 59924 163606 59952 465967
rect 60016 163742 60044 478722
rect 60568 476882 60596 480037
rect 60752 480023 61042 480051
rect 60556 476876 60608 476882
rect 60556 476818 60608 476824
rect 60752 462874 60780 480023
rect 61488 471209 61516 480037
rect 61672 480023 61962 480051
rect 62224 480023 62330 480051
rect 61474 471200 61530 471209
rect 61474 471135 61530 471144
rect 61672 470594 61700 480023
rect 62120 475380 62172 475386
rect 62120 475322 62172 475328
rect 60844 470566 61700 470594
rect 60844 465662 60872 470566
rect 62132 469130 62160 475322
rect 62120 469124 62172 469130
rect 62120 469066 62172 469072
rect 62224 469062 62252 480023
rect 62776 475114 62804 480037
rect 62960 480023 63250 480051
rect 63604 480023 63710 480051
rect 62960 475386 62988 480023
rect 62948 475380 63000 475386
rect 62948 475322 63000 475328
rect 63500 475380 63552 475386
rect 63500 475322 63552 475328
rect 62764 475108 62816 475114
rect 62764 475050 62816 475056
rect 62212 469056 62264 469062
rect 62212 468998 62264 469004
rect 60832 465656 60884 465662
rect 60832 465598 60884 465604
rect 60740 462868 60792 462874
rect 60740 462810 60792 462816
rect 63512 460494 63540 475322
rect 63500 460488 63552 460494
rect 63500 460430 63552 460436
rect 63604 460154 63632 480023
rect 64156 478106 64184 480037
rect 64248 480023 64538 480051
rect 64892 480023 64998 480051
rect 65076 480023 65458 480051
rect 65536 480023 65918 480051
rect 64144 478100 64196 478106
rect 64144 478042 64196 478048
rect 64248 475386 64276 480023
rect 64236 475380 64288 475386
rect 64236 475322 64288 475328
rect 64328 475380 64380 475386
rect 64328 475322 64380 475328
rect 64340 475114 64368 475322
rect 64328 475108 64380 475114
rect 64328 475050 64380 475056
rect 64892 462806 64920 480023
rect 64972 475108 65024 475114
rect 64972 475050 65024 475056
rect 64984 465594 65012 475050
rect 64972 465588 65024 465594
rect 64972 465530 65024 465536
rect 65076 465526 65104 480023
rect 65536 475114 65564 480023
rect 66364 478689 66392 480037
rect 66456 480023 66746 480051
rect 66824 480023 67206 480051
rect 66350 478680 66406 478689
rect 66350 478615 66406 478624
rect 65524 475108 65576 475114
rect 65524 475050 65576 475056
rect 66260 475108 66312 475114
rect 66260 475050 66312 475056
rect 65064 465520 65116 465526
rect 65064 465462 65116 465468
rect 64880 462800 64932 462806
rect 64880 462742 64932 462748
rect 63592 460148 63644 460154
rect 63592 460090 63644 460096
rect 66272 458658 66300 475050
rect 66456 470594 66484 480023
rect 66824 475114 66852 480023
rect 66812 475108 66864 475114
rect 66812 475050 66864 475056
rect 66364 470566 66484 470594
rect 66364 460562 66392 470566
rect 66352 460556 66404 460562
rect 66352 460498 66404 460504
rect 67652 459105 67680 480037
rect 67744 480023 68126 480051
rect 68204 480023 68494 480051
rect 68664 480023 68954 480051
rect 69032 480023 69414 480051
rect 69492 480023 69874 480051
rect 69952 480023 70334 480051
rect 70504 480023 70702 480051
rect 70872 480023 71162 480051
rect 71240 480023 71622 480051
rect 71792 480023 72082 480051
rect 72160 480023 72542 480051
rect 72620 480023 72910 480051
rect 67744 460057 67772 480023
rect 68204 470594 68232 480023
rect 68664 478825 68692 480023
rect 68650 478816 68706 478825
rect 68650 478751 68706 478760
rect 68926 478816 68982 478825
rect 68926 478751 68982 478760
rect 68940 478650 68968 478751
rect 68928 478644 68980 478650
rect 68928 478586 68980 478592
rect 68284 478576 68336 478582
rect 68284 478518 68336 478524
rect 67836 470566 68232 470594
rect 67836 460193 67864 470566
rect 68296 460222 68324 478518
rect 68376 478508 68428 478514
rect 68376 478450 68428 478456
rect 68388 466410 68416 478450
rect 68376 466404 68428 466410
rect 68376 466346 68428 466352
rect 68284 460216 68336 460222
rect 67822 460184 67878 460193
rect 68284 460158 68336 460164
rect 67822 460119 67878 460128
rect 67730 460048 67786 460057
rect 67730 459983 67786 459992
rect 67638 459096 67694 459105
rect 67638 459031 67694 459040
rect 69032 458969 69060 480023
rect 69492 475402 69520 480023
rect 69952 478258 69980 480023
rect 69124 475374 69520 475402
rect 69584 478230 69980 478258
rect 69124 460465 69152 475374
rect 69584 470594 69612 478230
rect 69664 478100 69716 478106
rect 69664 478042 69716 478048
rect 69216 470566 69612 470594
rect 69216 463185 69244 470566
rect 69202 463176 69258 463185
rect 69202 463111 69258 463120
rect 69110 460456 69166 460465
rect 69110 460391 69166 460400
rect 69676 460222 69704 478042
rect 70400 476128 70452 476134
rect 70400 476070 70452 476076
rect 70412 460426 70440 476070
rect 70504 463457 70532 480023
rect 70872 476134 70900 480023
rect 70860 476128 70912 476134
rect 70860 476070 70912 476076
rect 71240 475402 71268 480023
rect 71320 478644 71372 478650
rect 71320 478586 71372 478592
rect 70596 475374 71268 475402
rect 70596 468926 70624 475374
rect 71332 470594 71360 478586
rect 71056 470566 71360 470594
rect 71056 468994 71084 470566
rect 71044 468988 71096 468994
rect 71044 468930 71096 468936
rect 70584 468920 70636 468926
rect 70584 468862 70636 468868
rect 70490 463448 70546 463457
rect 70490 463383 70546 463392
rect 71792 460873 71820 480023
rect 71872 475108 71924 475114
rect 71872 475050 71924 475056
rect 71778 460864 71834 460873
rect 71778 460799 71834 460808
rect 70400 460420 70452 460426
rect 70400 460362 70452 460368
rect 71884 460358 71912 475050
rect 72160 470594 72188 480023
rect 72620 475114 72648 480023
rect 72608 475108 72660 475114
rect 72608 475050 72660 475056
rect 71976 470566 72188 470594
rect 71976 463321 72004 470566
rect 71962 463312 72018 463321
rect 71962 463247 72018 463256
rect 73356 461553 73384 480037
rect 73816 478009 73844 480037
rect 74276 478854 74304 480037
rect 74552 480023 74658 480051
rect 74736 480023 75118 480051
rect 75196 480023 75578 480051
rect 75932 480023 76038 480051
rect 76116 480023 76498 480051
rect 76576 480023 76866 480051
rect 74264 478848 74316 478854
rect 74264 478790 74316 478796
rect 73802 478000 73858 478009
rect 73802 477935 73858 477944
rect 73342 461544 73398 461553
rect 73342 461479 73398 461488
rect 71872 460352 71924 460358
rect 71872 460294 71924 460300
rect 74552 460290 74580 480023
rect 74736 475402 74764 480023
rect 74644 475374 74764 475402
rect 74644 460329 74672 475374
rect 75196 475266 75224 480023
rect 75368 478848 75420 478854
rect 75368 478790 75420 478796
rect 75276 478100 75328 478106
rect 75276 478042 75328 478048
rect 74736 475238 75224 475266
rect 74736 460601 74764 475238
rect 75288 474314 75316 478042
rect 75196 474286 75316 474314
rect 75196 466206 75224 474286
rect 75380 470594 75408 478790
rect 75826 478680 75882 478689
rect 75826 478615 75882 478624
rect 75840 477970 75868 478615
rect 75828 477964 75880 477970
rect 75828 477906 75880 477912
rect 75288 470566 75408 470594
rect 75288 468858 75316 470566
rect 75276 468852 75328 468858
rect 75276 468794 75328 468800
rect 75184 466200 75236 466206
rect 75184 466142 75236 466148
rect 75932 460737 75960 480023
rect 76116 475402 76144 480023
rect 76024 475374 76144 475402
rect 75918 460728 75974 460737
rect 76024 460698 76052 475374
rect 76576 470594 76604 480023
rect 77312 478417 77340 480037
rect 77772 478553 77800 480037
rect 77864 480023 78246 480051
rect 77758 478544 77814 478553
rect 77758 478479 77814 478488
rect 77298 478408 77354 478417
rect 77298 478343 77354 478352
rect 77864 470594 77892 480023
rect 78692 478689 78720 480037
rect 78784 480023 79074 480051
rect 78678 478680 78734 478689
rect 78678 478615 78734 478624
rect 78680 475108 78732 475114
rect 78680 475050 78732 475056
rect 76116 470566 76604 470594
rect 77312 470566 77892 470594
rect 76116 460766 76144 470566
rect 76104 460760 76156 460766
rect 76104 460702 76156 460708
rect 75918 460663 75974 460672
rect 76012 460692 76064 460698
rect 76012 460634 76064 460640
rect 77312 460630 77340 470566
rect 78692 460834 78720 475050
rect 78784 460902 78812 480023
rect 79520 478825 79548 480037
rect 79704 480023 79994 480051
rect 80164 480023 80454 480051
rect 80532 480023 80822 480051
rect 79506 478816 79562 478825
rect 79506 478751 79562 478760
rect 79704 475114 79732 480023
rect 79692 475108 79744 475114
rect 79692 475050 79744 475056
rect 80164 463049 80192 480023
rect 80532 470594 80560 480023
rect 81268 477902 81296 480037
rect 81728 478038 81756 480037
rect 81912 480023 82202 480051
rect 82280 480023 82662 480051
rect 82924 480023 83030 480051
rect 83108 480023 83490 480051
rect 83568 480023 83950 480051
rect 81716 478032 81768 478038
rect 81716 477974 81768 477980
rect 81256 477896 81308 477902
rect 81256 477838 81308 477844
rect 81532 473612 81584 473618
rect 81532 473554 81584 473560
rect 80256 470566 80560 470594
rect 80150 463040 80206 463049
rect 80150 462975 80206 462984
rect 78772 460896 78824 460902
rect 78772 460838 78824 460844
rect 78680 460828 78732 460834
rect 78680 460770 78732 460776
rect 77300 460624 77352 460630
rect 74722 460592 74778 460601
rect 77300 460566 77352 460572
rect 74722 460527 74778 460536
rect 74630 460320 74686 460329
rect 74540 460284 74592 460290
rect 74630 460255 74686 460264
rect 74540 460226 74592 460232
rect 69664 460216 69716 460222
rect 69664 460158 69716 460164
rect 69018 458960 69074 458969
rect 69018 458895 69074 458904
rect 80256 458833 80284 470566
rect 81544 466138 81572 473554
rect 81912 470594 81940 480023
rect 82280 473618 82308 480023
rect 82820 475108 82872 475114
rect 82820 475050 82872 475056
rect 82268 473612 82320 473618
rect 82268 473554 82320 473560
rect 81636 470566 81940 470594
rect 81532 466132 81584 466138
rect 81532 466074 81584 466080
rect 81636 463554 81664 470566
rect 82832 466342 82860 475050
rect 82820 466336 82872 466342
rect 82820 466278 82872 466284
rect 82924 466274 82952 480023
rect 83108 470594 83136 480023
rect 83568 475114 83596 480023
rect 84396 479194 84424 480037
rect 84384 479188 84436 479194
rect 84384 479130 84436 479136
rect 84856 478718 84884 480037
rect 84948 480023 85238 480051
rect 85698 480023 85804 480051
rect 84844 478712 84896 478718
rect 84844 478654 84896 478660
rect 83556 475108 83608 475114
rect 83556 475050 83608 475056
rect 84948 470594 84976 480023
rect 85776 476134 85804 480023
rect 85868 480023 86158 480051
rect 86328 480023 86618 480051
rect 87078 480023 87184 480051
rect 85764 476128 85816 476134
rect 85764 476070 85816 476076
rect 85868 475538 85896 480023
rect 85948 476128 86000 476134
rect 85948 476070 86000 476076
rect 83016 470566 83136 470594
rect 84304 470566 84976 470594
rect 85592 475510 85896 475538
rect 82912 466268 82964 466274
rect 82912 466210 82964 466216
rect 83016 466070 83044 470566
rect 83004 466064 83056 466070
rect 83004 466006 83056 466012
rect 84304 465905 84332 470566
rect 84290 465896 84346 465905
rect 84290 465831 84346 465840
rect 81624 463548 81676 463554
rect 81624 463490 81676 463496
rect 85592 462942 85620 475510
rect 85672 475108 85724 475114
rect 85672 475050 85724 475056
rect 85684 463350 85712 475050
rect 85960 470594 85988 476070
rect 86328 475114 86356 480023
rect 86316 475108 86368 475114
rect 86316 475050 86368 475056
rect 87052 475108 87104 475114
rect 87052 475050 87104 475056
rect 86960 475040 87012 475046
rect 86960 474982 87012 474988
rect 85776 470566 85988 470594
rect 85776 466177 85804 470566
rect 85762 466168 85818 466177
rect 85762 466103 85818 466112
rect 86972 463622 87000 474982
rect 86960 463616 87012 463622
rect 86960 463558 87012 463564
rect 85672 463344 85724 463350
rect 85672 463286 85724 463292
rect 87064 463078 87092 475050
rect 87156 463690 87184 480023
rect 87248 480023 87446 480051
rect 87616 480023 87906 480051
rect 88366 480023 88656 480051
rect 87248 475114 87276 480023
rect 87236 475108 87288 475114
rect 87236 475050 87288 475056
rect 87616 475046 87644 480023
rect 88432 475108 88484 475114
rect 88432 475050 88484 475056
rect 87604 475040 87656 475046
rect 87604 474982 87656 474988
rect 87144 463684 87196 463690
rect 87144 463626 87196 463632
rect 88444 463486 88472 475050
rect 88524 475040 88576 475046
rect 88524 474982 88576 474988
rect 88432 463480 88484 463486
rect 88432 463422 88484 463428
rect 88536 463214 88564 474982
rect 88628 463418 88656 480023
rect 88720 480023 88826 480051
rect 88904 480023 89194 480051
rect 88720 475046 88748 480023
rect 88904 475114 88932 480023
rect 89640 478174 89668 480037
rect 89732 480023 90114 480051
rect 90192 480023 90574 480051
rect 90744 480023 91034 480051
rect 89628 478168 89680 478174
rect 89628 478110 89680 478116
rect 88892 475108 88944 475114
rect 88892 475050 88944 475056
rect 88708 475040 88760 475046
rect 88708 474982 88760 474988
rect 88616 463412 88668 463418
rect 88616 463354 88668 463360
rect 89732 463282 89760 480023
rect 89812 475108 89864 475114
rect 89812 475050 89864 475056
rect 89824 466449 89852 475050
rect 90192 470594 90220 480023
rect 90744 475114 90772 480023
rect 91388 478281 91416 480037
rect 91848 478786 91876 480037
rect 91940 480023 92322 480051
rect 92676 480023 92782 480051
rect 92952 480023 93242 480051
rect 93320 480023 93610 480051
rect 91836 478780 91888 478786
rect 91836 478722 91888 478728
rect 91374 478272 91430 478281
rect 91374 478207 91430 478216
rect 90732 475108 90784 475114
rect 90732 475050 90784 475056
rect 91940 470594 91968 480023
rect 92480 475108 92532 475114
rect 92480 475050 92532 475056
rect 89916 470566 90220 470594
rect 91296 470566 91968 470594
rect 89810 466440 89866 466449
rect 89810 466375 89866 466384
rect 89916 465769 89944 470566
rect 91296 466313 91324 470566
rect 91282 466304 91338 466313
rect 91282 466239 91338 466248
rect 89902 465760 89958 465769
rect 89902 465695 89958 465704
rect 89720 463276 89772 463282
rect 89720 463218 89772 463224
rect 88524 463208 88576 463214
rect 88524 463150 88576 463156
rect 87052 463072 87104 463078
rect 87052 463014 87104 463020
rect 85580 462936 85632 462942
rect 85580 462878 85632 462884
rect 92492 459338 92520 475050
rect 92572 475040 92624 475046
rect 92572 474982 92624 474988
rect 92584 463010 92612 474982
rect 92676 466041 92704 480023
rect 92952 475114 92980 480023
rect 92940 475108 92992 475114
rect 92940 475050 92992 475056
rect 93320 475046 93348 480023
rect 94056 478145 94084 480037
rect 94148 480023 94530 480051
rect 94608 480023 94990 480051
rect 94042 478136 94098 478145
rect 94042 478071 94098 478080
rect 94148 475402 94176 480023
rect 93872 475374 94176 475402
rect 93308 475040 93360 475046
rect 93308 474982 93360 474988
rect 92662 466032 92718 466041
rect 92662 465967 92718 465976
rect 92572 463004 92624 463010
rect 92572 462946 92624 462952
rect 93872 462913 93900 475374
rect 94608 470594 94636 480023
rect 95344 478174 95372 480037
rect 95332 478168 95384 478174
rect 95332 478110 95384 478116
rect 95804 475969 95832 480037
rect 95790 475960 95846 475969
rect 95790 475895 95846 475904
rect 96264 474094 96292 480037
rect 96724 475182 96752 480037
rect 97184 478242 97212 480037
rect 97552 478378 97580 480037
rect 97540 478372 97592 478378
rect 97540 478314 97592 478320
rect 97172 478236 97224 478242
rect 97172 478178 97224 478184
rect 98012 475318 98040 480037
rect 98000 475312 98052 475318
rect 98000 475254 98052 475260
rect 98472 475250 98500 480037
rect 98932 479058 98960 480037
rect 99392 479126 99420 480037
rect 99380 479120 99432 479126
rect 99380 479062 99432 479068
rect 98920 479052 98972 479058
rect 98920 478994 98972 479000
rect 99760 478310 99788 480037
rect 100220 478990 100248 480037
rect 100312 480023 100694 480051
rect 100956 480023 101154 480051
rect 101232 480023 101522 480051
rect 101600 480023 101982 480051
rect 100208 478984 100260 478990
rect 100208 478926 100260 478932
rect 99748 478304 99800 478310
rect 99748 478246 99800 478252
rect 98460 475244 98512 475250
rect 98460 475186 98512 475192
rect 96712 475176 96764 475182
rect 96712 475118 96764 475124
rect 96252 474088 96304 474094
rect 96252 474030 96304 474036
rect 100312 470594 100340 480023
rect 100852 475312 100904 475318
rect 100852 475254 100904 475260
rect 100760 475244 100812 475250
rect 100760 475186 100812 475192
rect 93964 470566 94636 470594
rect 99484 470566 100340 470594
rect 93964 468790 93992 470566
rect 93952 468784 94004 468790
rect 93952 468726 94004 468732
rect 93858 462904 93914 462913
rect 93858 462839 93914 462848
rect 92480 459332 92532 459338
rect 92480 459274 92532 459280
rect 99484 459202 99512 470566
rect 99472 459196 99524 459202
rect 99472 459138 99524 459144
rect 100772 459134 100800 475186
rect 100864 465866 100892 475254
rect 100852 465860 100904 465866
rect 100852 465802 100904 465808
rect 100956 465730 100984 480023
rect 101232 475318 101260 480023
rect 101220 475312 101272 475318
rect 101220 475254 101272 475260
rect 101600 475250 101628 480023
rect 102428 478446 102456 480037
rect 102416 478440 102468 478446
rect 102416 478382 102468 478388
rect 102888 478106 102916 480037
rect 103072 480023 103362 480051
rect 102876 478100 102928 478106
rect 102876 478042 102928 478048
rect 101588 475244 101640 475250
rect 101588 475186 101640 475192
rect 103072 470594 103100 480023
rect 103612 475312 103664 475318
rect 103612 475254 103664 475260
rect 102244 470566 103100 470594
rect 102244 466002 102272 470566
rect 102232 465996 102284 466002
rect 102232 465938 102284 465944
rect 103624 465934 103652 475254
rect 103612 465928 103664 465934
rect 103612 465870 103664 465876
rect 100944 465724 100996 465730
rect 100944 465666 100996 465672
rect 103716 459270 103744 480037
rect 103808 480023 104190 480051
rect 103808 475318 103836 480023
rect 104636 478582 104664 480037
rect 105096 478922 105124 480037
rect 105084 478916 105136 478922
rect 105084 478858 105136 478864
rect 104624 478576 104676 478582
rect 104624 478518 104676 478524
rect 105556 478514 105584 480037
rect 105648 480023 105938 480051
rect 105544 478508 105596 478514
rect 105544 478450 105596 478456
rect 103796 475312 103848 475318
rect 103796 475254 103848 475260
rect 105648 470594 105676 480023
rect 106384 478650 106412 480037
rect 106568 480023 106858 480051
rect 106372 478644 106424 478650
rect 106372 478586 106424 478592
rect 106568 470594 106596 480023
rect 107304 478854 107332 480037
rect 107292 478848 107344 478854
rect 107292 478790 107344 478796
rect 107660 475312 107712 475318
rect 107660 475254 107712 475260
rect 105004 470566 105676 470594
rect 106384 470566 106596 470594
rect 105004 468722 105032 470566
rect 104992 468716 105044 468722
rect 104992 468658 105044 468664
rect 106384 468654 106412 470566
rect 106372 468648 106424 468654
rect 106372 468590 106424 468596
rect 107672 463010 107700 475254
rect 107660 463004 107712 463010
rect 107660 462946 107712 462952
rect 107764 462913 107792 480037
rect 107856 480023 108146 480051
rect 108224 480023 108606 480051
rect 107856 475318 107884 480023
rect 107844 475312 107896 475318
rect 107844 475254 107896 475260
rect 108224 470594 108252 480023
rect 109052 478990 109080 480037
rect 109040 478984 109092 478990
rect 109040 478926 109092 478932
rect 109512 478922 109540 480037
rect 109500 478916 109552 478922
rect 109500 478858 109552 478864
rect 109880 478242 109908 480037
rect 110064 480023 110354 480051
rect 110616 480023 110814 480051
rect 109868 478236 109920 478242
rect 109868 478178 109920 478184
rect 110064 470594 110092 480023
rect 107856 470566 108252 470594
rect 109052 470566 110092 470594
rect 107856 465730 107884 470566
rect 107844 465724 107896 465730
rect 107844 465666 107896 465672
rect 109052 463078 109080 470566
rect 110616 465798 110644 480023
rect 111260 475998 111288 480037
rect 111720 476066 111748 480037
rect 111708 476060 111760 476066
rect 111708 476002 111760 476008
rect 111248 475992 111300 475998
rect 111248 475934 111300 475940
rect 112088 475794 112116 480037
rect 112548 475862 112576 480037
rect 112640 480023 113022 480051
rect 113376 480023 113482 480051
rect 112536 475856 112588 475862
rect 112536 475798 112588 475804
rect 112076 475788 112128 475794
rect 112076 475730 112128 475736
rect 112640 470594 112668 480023
rect 111996 470566 112668 470594
rect 110604 465792 110656 465798
rect 110604 465734 110656 465740
rect 111996 464370 112024 470566
rect 111984 464364 112036 464370
rect 111984 464306 112036 464312
rect 113376 463146 113404 480023
rect 113928 471306 113956 480037
rect 114296 472462 114324 480037
rect 114284 472456 114336 472462
rect 114284 472398 114336 472404
rect 113916 471300 113968 471306
rect 113916 471242 113968 471248
rect 114756 467158 114784 480037
rect 115216 475930 115244 480037
rect 115204 475924 115256 475930
rect 115204 475866 115256 475872
rect 115676 475658 115704 480037
rect 116044 475726 116072 480037
rect 116032 475720 116084 475726
rect 116032 475662 116084 475668
rect 115664 475652 115716 475658
rect 115664 475594 115716 475600
rect 116504 473346 116532 480037
rect 116492 473340 116544 473346
rect 116492 473282 116544 473288
rect 116964 472598 116992 480037
rect 116952 472592 117004 472598
rect 116952 472534 117004 472540
rect 117424 472530 117452 480037
rect 117884 476950 117912 480037
rect 117872 476944 117924 476950
rect 117872 476886 117924 476892
rect 118252 473142 118280 480037
rect 118726 480023 118924 480051
rect 118240 473136 118292 473142
rect 118240 473078 118292 473084
rect 117412 472524 117464 472530
rect 117412 472466 117464 472472
rect 114744 467152 114796 467158
rect 114744 467094 114796 467100
rect 113364 463140 113416 463146
rect 113364 463082 113416 463088
rect 109040 463072 109092 463078
rect 109040 463014 109092 463020
rect 107750 462904 107806 462913
rect 107750 462839 107806 462848
rect 103704 459264 103756 459270
rect 103704 459206 103756 459212
rect 100760 459128 100812 459134
rect 100760 459070 100812 459076
rect 118896 459066 118924 480023
rect 119172 472705 119200 480037
rect 119632 475590 119660 480037
rect 119620 475584 119672 475590
rect 120092 475561 120120 480037
rect 120184 480023 120474 480051
rect 119620 475526 119672 475532
rect 120078 475552 120134 475561
rect 120078 475487 120134 475496
rect 119158 472696 119214 472705
rect 119158 472631 119214 472640
rect 120184 470558 120212 480023
rect 120724 476876 120776 476882
rect 120724 476818 120776 476824
rect 120736 476746 120764 476818
rect 120724 476740 120776 476746
rect 120724 476682 120776 476688
rect 120920 475697 120948 480037
rect 121380 475833 121408 480037
rect 121748 480023 121854 480051
rect 121932 480023 122222 480051
rect 122392 480023 122682 480051
rect 122852 480023 123142 480051
rect 121366 475824 121422 475833
rect 121366 475759 121422 475768
rect 120906 475688 120962 475697
rect 120906 475623 120962 475632
rect 120172 470552 120224 470558
rect 120172 470494 120224 470500
rect 121748 470490 121776 480023
rect 121736 470484 121788 470490
rect 121736 470426 121788 470432
rect 121932 470354 121960 480023
rect 121920 470348 121972 470354
rect 121920 470290 121972 470296
rect 122392 466454 122420 480023
rect 122852 470218 122880 480023
rect 123588 472569 123616 480037
rect 123680 480023 124062 480051
rect 124232 480023 124430 480051
rect 124508 480023 124890 480051
rect 124968 480023 125350 480051
rect 123574 472560 123630 472569
rect 123574 472495 123630 472504
rect 122840 470212 122892 470218
rect 122840 470154 122892 470160
rect 123680 470082 123708 480023
rect 123668 470076 123720 470082
rect 123668 470018 123720 470024
rect 124232 470014 124260 480023
rect 124508 470150 124536 480023
rect 124968 470286 124996 480023
rect 124956 470280 125008 470286
rect 124956 470222 125008 470228
rect 124496 470144 124548 470150
rect 124496 470086 124548 470092
rect 124220 470008 124272 470014
rect 124220 469950 124272 469956
rect 125796 469849 125824 480037
rect 125888 480023 126270 480051
rect 125888 469985 125916 480023
rect 126624 475425 126652 480037
rect 126610 475416 126666 475425
rect 126610 475351 126666 475360
rect 125874 469976 125930 469985
rect 125874 469911 125930 469920
rect 125782 469840 125838 469849
rect 125782 469775 125838 469784
rect 127084 468489 127112 480037
rect 127176 480023 127558 480051
rect 127728 480023 128018 480051
rect 127176 469810 127204 480023
rect 127164 469804 127216 469810
rect 127164 469746 127216 469752
rect 127728 468654 127756 480023
rect 128464 469742 128492 480037
rect 128556 480023 128846 480051
rect 128452 469736 128504 469742
rect 128452 469678 128504 469684
rect 128556 469674 128584 480023
rect 129292 472802 129320 480037
rect 129752 472870 129780 480037
rect 130028 480023 130226 480051
rect 129740 472864 129792 472870
rect 129740 472806 129792 472812
rect 129280 472796 129332 472802
rect 129280 472738 129332 472744
rect 128544 469668 128596 469674
rect 128544 469610 128596 469616
rect 127716 468648 127768 468654
rect 127716 468590 127768 468596
rect 127070 468480 127126 468489
rect 127070 468415 127126 468424
rect 121472 466426 122420 466454
rect 118884 459060 118936 459066
rect 118884 459002 118936 459008
rect 121472 458998 121500 466426
rect 121460 458992 121512 458998
rect 121460 458934 121512 458940
rect 130028 458930 130056 480023
rect 130580 473278 130608 480037
rect 130568 473272 130620 473278
rect 130568 473214 130620 473220
rect 131040 473074 131068 480037
rect 131028 473068 131080 473074
rect 131028 473010 131080 473016
rect 131500 473006 131528 480037
rect 131488 473000 131540 473006
rect 131488 472942 131540 472948
rect 131960 472734 131988 480037
rect 132420 475522 132448 480037
rect 132512 480023 132802 480051
rect 132880 480023 133262 480051
rect 133340 480023 133722 480051
rect 132408 475516 132460 475522
rect 132408 475458 132460 475464
rect 131948 472728 132000 472734
rect 131948 472670 132000 472676
rect 132512 472666 132540 480023
rect 132880 475504 132908 480023
rect 133340 476762 133368 480023
rect 132604 475476 132908 475504
rect 133064 476734 133368 476762
rect 132604 473210 132632 475476
rect 132592 473204 132644 473210
rect 132592 473146 132644 473152
rect 132500 472660 132552 472666
rect 132500 472602 132552 472608
rect 133064 470594 133092 476734
rect 133144 476672 133196 476678
rect 133144 476614 133196 476620
rect 132696 470566 133092 470594
rect 132696 469946 132724 470566
rect 132684 469940 132736 469946
rect 132684 469882 132736 469888
rect 133156 462330 133184 476614
rect 133972 475312 134024 475318
rect 133972 475254 134024 475260
rect 133984 470422 134012 475254
rect 134168 472938 134196 480037
rect 134260 480023 134642 480051
rect 134720 480023 135010 480051
rect 134156 472932 134208 472938
rect 134156 472874 134208 472880
rect 134260 470594 134288 480023
rect 134720 475318 134748 480023
rect 134708 475312 134760 475318
rect 134708 475254 134760 475260
rect 134076 470566 134288 470594
rect 133972 470416 134024 470422
rect 133972 470358 134024 470364
rect 133144 462324 133196 462330
rect 133144 462266 133196 462272
rect 130016 458924 130068 458930
rect 130016 458866 130068 458872
rect 134076 458862 134104 470566
rect 135456 458998 135484 480037
rect 135916 475454 135944 480037
rect 136376 475726 136404 480037
rect 136364 475720 136416 475726
rect 136364 475662 136416 475668
rect 136744 475590 136772 480037
rect 136836 480023 137218 480051
rect 136732 475584 136784 475590
rect 136732 475526 136784 475532
rect 135904 475448 135956 475454
rect 135904 475390 135956 475396
rect 136836 470594 136864 480023
rect 137664 475522 137692 480037
rect 138124 475658 138152 480037
rect 138216 480023 138598 480051
rect 138112 475652 138164 475658
rect 138112 475594 138164 475600
rect 137652 475516 137704 475522
rect 137652 475458 137704 475464
rect 138216 470594 138244 480023
rect 138952 478310 138980 480037
rect 138940 478304 138992 478310
rect 138940 478246 138992 478252
rect 139412 477970 139440 480037
rect 139504 480023 139886 480051
rect 140056 480023 140346 480051
rect 139400 477964 139452 477970
rect 139400 477906 139452 477912
rect 139400 475312 139452 475318
rect 139400 475254 139452 475260
rect 136652 470566 136864 470594
rect 138032 470566 138244 470594
rect 135444 458992 135496 458998
rect 135444 458934 135496 458940
rect 136652 458930 136680 470566
rect 136640 458924 136692 458930
rect 136640 458866 136692 458872
rect 138032 458862 138060 470566
rect 139412 466002 139440 475254
rect 139504 468722 139532 480023
rect 140056 475318 140084 480023
rect 140792 479058 140820 480037
rect 140976 480023 141174 480051
rect 141344 480023 141634 480051
rect 141712 480023 142094 480051
rect 142356 480023 142554 480051
rect 142632 480023 142922 480051
rect 143000 480023 143382 480051
rect 143644 480023 143842 480051
rect 143920 480023 144302 480051
rect 140780 479052 140832 479058
rect 140780 478994 140832 479000
rect 140780 475448 140832 475454
rect 140780 475390 140832 475396
rect 140044 475312 140096 475318
rect 140044 475254 140096 475260
rect 139492 468716 139544 468722
rect 139492 468658 139544 468664
rect 139400 465996 139452 466002
rect 139400 465938 139452 465944
rect 140792 465866 140820 475390
rect 140872 475312 140924 475318
rect 140872 475254 140924 475260
rect 140780 465860 140832 465866
rect 140780 465802 140832 465808
rect 140884 465798 140912 475254
rect 140976 465934 141004 480023
rect 141344 475318 141372 480023
rect 141712 475454 141740 480023
rect 141884 475720 141936 475726
rect 141884 475662 141936 475668
rect 141896 475522 141924 475662
rect 141884 475516 141936 475522
rect 141884 475458 141936 475464
rect 141700 475448 141752 475454
rect 141700 475390 141752 475396
rect 141332 475312 141384 475318
rect 141332 475254 141384 475260
rect 142252 475312 142304 475318
rect 142252 475254 142304 475260
rect 142160 475244 142212 475250
rect 142160 475186 142212 475192
rect 140964 465928 141016 465934
rect 140964 465870 141016 465876
rect 140872 465792 140924 465798
rect 140872 465734 140924 465740
rect 142172 459066 142200 475186
rect 142264 459134 142292 475254
rect 142356 463146 142384 480023
rect 142632 475318 142660 480023
rect 142620 475312 142672 475318
rect 142620 475254 142672 475260
rect 143000 475250 143028 480023
rect 143540 475312 143592 475318
rect 143540 475254 143592 475260
rect 142988 475244 143040 475250
rect 142988 475186 143040 475192
rect 142344 463140 142396 463146
rect 142344 463082 142396 463088
rect 143552 460329 143580 475254
rect 143644 469878 143672 480023
rect 143920 475318 143948 480023
rect 143908 475312 143960 475318
rect 143908 475254 143960 475260
rect 144748 474201 144776 480037
rect 145116 475425 145144 480037
rect 145102 475416 145158 475425
rect 145102 475351 145158 475360
rect 144734 474192 144790 474201
rect 144734 474127 144790 474136
rect 145576 471345 145604 480037
rect 146036 478145 146064 480037
rect 146022 478136 146078 478145
rect 146022 478071 146078 478080
rect 146496 475561 146524 480037
rect 146482 475552 146538 475561
rect 146482 475487 146538 475496
rect 146956 474337 146984 480037
rect 147324 478417 147352 480037
rect 147692 480023 147798 480051
rect 147310 478408 147366 478417
rect 147310 478343 147366 478352
rect 146942 474328 146998 474337
rect 146942 474263 146998 474272
rect 145562 471336 145618 471345
rect 145562 471271 145618 471280
rect 143632 469872 143684 469878
rect 143632 469814 143684 469820
rect 147692 463049 147720 480023
rect 148244 478281 148272 480037
rect 148230 478272 148286 478281
rect 148230 478207 148286 478216
rect 148704 475697 148732 480037
rect 149164 478582 149192 480037
rect 149532 478854 149560 480037
rect 149520 478848 149572 478854
rect 149520 478790 149572 478796
rect 149152 478576 149204 478582
rect 149152 478518 149204 478524
rect 148690 475688 148746 475697
rect 148690 475623 148746 475632
rect 149992 471617 150020 480037
rect 150452 478106 150480 480037
rect 150544 480023 150926 480051
rect 150440 478100 150492 478106
rect 150440 478042 150492 478048
rect 150440 475312 150492 475318
rect 150440 475254 150492 475260
rect 149978 471608 150034 471617
rect 149978 471543 150034 471552
rect 147678 463040 147734 463049
rect 147678 462975 147734 462984
rect 143538 460320 143594 460329
rect 143538 460255 143594 460264
rect 150452 460193 150480 475254
rect 150544 469849 150572 480023
rect 151280 478514 151308 480037
rect 151464 480023 151754 480051
rect 151268 478508 151320 478514
rect 151268 478450 151320 478456
rect 151464 475318 151492 480023
rect 152200 478786 152228 480037
rect 152188 478780 152240 478786
rect 152188 478722 152240 478728
rect 151452 475312 151504 475318
rect 151452 475254 151504 475260
rect 152660 474065 152688 480037
rect 153120 478650 153148 480037
rect 153108 478644 153160 478650
rect 153108 478586 153160 478592
rect 153488 478378 153516 480037
rect 153476 478372 153528 478378
rect 153476 478314 153528 478320
rect 152646 474056 152702 474065
rect 152646 473991 152702 474000
rect 153948 472569 153976 480037
rect 154408 478718 154436 480037
rect 154396 478712 154448 478718
rect 154396 478654 154448 478660
rect 154868 476921 154896 480037
rect 154960 480023 155342 480051
rect 155420 480023 155710 480051
rect 155972 480023 156170 480051
rect 154854 476912 154910 476921
rect 154854 476847 154910 476856
rect 154960 475402 154988 480023
rect 154592 475374 154988 475402
rect 153934 472560 153990 472569
rect 153934 472495 153990 472504
rect 150530 469840 150586 469849
rect 150530 469775 150586 469784
rect 154592 460465 154620 475374
rect 155420 470594 155448 480023
rect 154684 470566 155448 470594
rect 154684 463185 154712 470566
rect 155972 468625 156000 480023
rect 156616 478038 156644 480037
rect 156800 480023 157090 480051
rect 157352 480023 157458 480051
rect 156604 478032 156656 478038
rect 156604 477974 156656 477980
rect 156800 470594 156828 480023
rect 156064 470566 156828 470594
rect 156064 469985 156092 470566
rect 156050 469976 156106 469985
rect 156050 469911 156106 469920
rect 155958 468616 156014 468625
rect 155958 468551 156014 468560
rect 154670 463176 154726 463185
rect 154670 463111 154726 463120
rect 157352 460902 157380 480023
rect 157904 478446 157932 480037
rect 158088 480023 158378 480051
rect 157892 478440 157944 478446
rect 157892 478382 157944 478388
rect 158088 470594 158116 480023
rect 158824 472841 158852 480037
rect 159008 480023 159298 480051
rect 158810 472832 158866 472841
rect 158810 472767 158866 472776
rect 159008 470594 159036 480023
rect 159652 476882 159680 480037
rect 160126 480023 160156 480051
rect 160128 479874 160156 480023
rect 160204 480023 160586 480051
rect 160664 480023 161046 480051
rect 161506 480023 161704 480051
rect 160116 479868 160168 479874
rect 160116 479810 160168 479816
rect 159640 476876 159692 476882
rect 159640 476818 159692 476824
rect 160100 475312 160152 475318
rect 160100 475254 160152 475260
rect 157444 470566 158116 470594
rect 158732 470566 159036 470594
rect 157444 467129 157472 470566
rect 157430 467120 157486 467129
rect 157430 467055 157486 467064
rect 158732 464370 158760 470566
rect 158720 464364 158772 464370
rect 158720 464306 158772 464312
rect 160112 463214 160140 475254
rect 160204 467265 160232 480023
rect 160284 479868 160336 479874
rect 160284 479810 160336 479816
rect 160296 471481 160324 479810
rect 160664 475318 160692 480023
rect 160652 475312 160704 475318
rect 160652 475254 160704 475260
rect 161572 475312 161624 475318
rect 161572 475254 161624 475260
rect 161480 475244 161532 475250
rect 161480 475186 161532 475192
rect 160282 471472 160338 471481
rect 160282 471407 160338 471416
rect 160190 467256 160246 467265
rect 160190 467191 160246 467200
rect 160100 463208 160152 463214
rect 160100 463150 160152 463156
rect 157340 460896 157392 460902
rect 157340 460838 157392 460844
rect 154578 460456 154634 460465
rect 154578 460391 154634 460400
rect 150438 460184 150494 460193
rect 150438 460119 150494 460128
rect 142252 459128 142304 459134
rect 142252 459070 142304 459076
rect 142160 459060 142212 459066
rect 142160 459002 142212 459008
rect 134064 458856 134116 458862
rect 80242 458824 80298 458833
rect 134064 458798 134116 458804
rect 138020 458856 138072 458862
rect 161492 458833 161520 475186
rect 161584 461650 161612 475254
rect 161676 466041 161704 480023
rect 161768 480023 161874 480051
rect 161952 480023 162334 480051
rect 162504 480023 162794 480051
rect 162872 480023 163254 480051
rect 161768 475250 161796 480023
rect 161952 475318 161980 480023
rect 161940 475312 161992 475318
rect 161940 475254 161992 475260
rect 161756 475244 161808 475250
rect 161756 475186 161808 475192
rect 162504 470594 162532 480023
rect 161768 470566 162532 470594
rect 161768 468858 161796 470566
rect 161756 468852 161808 468858
rect 161756 468794 161808 468800
rect 161662 466032 161718 466041
rect 161662 465967 161718 465976
rect 162872 465905 162900 480023
rect 163608 478553 163636 480037
rect 163700 480023 164082 480051
rect 163594 478544 163650 478553
rect 163594 478479 163650 478488
rect 163700 470594 163728 480023
rect 164528 472705 164556 480037
rect 164620 480023 165002 480051
rect 165080 480023 165462 480051
rect 165724 480023 165830 480051
rect 164514 472696 164570 472705
rect 164514 472631 164570 472640
rect 164620 472546 164648 480023
rect 162964 470566 163728 470594
rect 164252 472518 164648 472546
rect 162964 468790 162992 470566
rect 162952 468784 163004 468790
rect 162952 468726 163004 468732
rect 162858 465896 162914 465905
rect 162858 465831 162914 465840
rect 161572 461644 161624 461650
rect 161572 461586 161624 461592
rect 164252 458969 164280 472518
rect 165080 470594 165108 480023
rect 165620 475312 165672 475318
rect 165620 475254 165672 475260
rect 164344 470566 165108 470594
rect 164344 460290 164372 470566
rect 165632 460601 165660 475254
rect 165724 469878 165752 480023
rect 166276 474026 166304 480037
rect 166368 480023 166750 480051
rect 166368 475318 166396 480023
rect 167196 478689 167224 480037
rect 167288 480023 167670 480051
rect 167748 480023 168038 480051
rect 168392 480023 168498 480051
rect 167182 478680 167238 478689
rect 167182 478615 167238 478624
rect 166356 475312 166408 475318
rect 166356 475254 166408 475260
rect 167000 475312 167052 475318
rect 167000 475254 167052 475260
rect 166264 474020 166316 474026
rect 166264 473962 166316 473968
rect 165712 469872 165764 469878
rect 165712 469814 165764 469820
rect 167012 460737 167040 475254
rect 167288 470594 167316 480023
rect 167748 475318 167776 480023
rect 167736 475312 167788 475318
rect 167736 475254 167788 475260
rect 167104 470566 167316 470594
rect 167104 465769 167132 470566
rect 167090 465760 167146 465769
rect 167090 465695 167146 465704
rect 168392 463282 168420 480023
rect 168944 477902 168972 480037
rect 169024 478236 169076 478242
rect 169024 478178 169076 478184
rect 168932 477896 168984 477902
rect 168932 477838 168984 477844
rect 168380 463276 168432 463282
rect 168380 463218 168432 463224
rect 166998 460728 167054 460737
rect 166998 460663 167054 460672
rect 165618 460592 165674 460601
rect 169036 460562 169064 478178
rect 169404 471306 169432 480037
rect 169772 480023 169878 480051
rect 169956 480023 170246 480051
rect 170324 480023 170706 480051
rect 171166 480023 171272 480051
rect 169392 471300 169444 471306
rect 169392 471242 169444 471248
rect 169772 463321 169800 480023
rect 169956 475402 169984 480023
rect 169864 475374 169984 475402
rect 169864 466177 169892 475374
rect 170324 470594 170352 480023
rect 171140 475720 171192 475726
rect 171140 475662 171192 475668
rect 169956 470566 170352 470594
rect 169850 466168 169906 466177
rect 169850 466103 169906 466112
rect 169956 463457 169984 470566
rect 169942 463448 169998 463457
rect 169942 463383 169998 463392
rect 169758 463312 169814 463321
rect 169758 463247 169814 463256
rect 165618 460527 165674 460536
rect 169024 460556 169076 460562
rect 169024 460498 169076 460504
rect 164332 460284 164384 460290
rect 164332 460226 164384 460232
rect 171152 459105 171180 475662
rect 171244 460873 171272 480023
rect 171336 480023 171626 480051
rect 171704 480023 171994 480051
rect 172072 480023 172454 480051
rect 171336 475726 171364 480023
rect 171324 475720 171376 475726
rect 171324 475662 171376 475668
rect 171704 475402 171732 480023
rect 171336 475374 171732 475402
rect 171230 460864 171286 460873
rect 171230 460799 171286 460808
rect 171336 459377 171364 475374
rect 172072 470594 172100 480023
rect 172900 478825 172928 480037
rect 172992 480023 173374 480051
rect 173544 480023 173834 480051
rect 173912 480023 174202 480051
rect 174280 480023 174662 480051
rect 174740 480023 175122 480051
rect 172886 478816 172942 478825
rect 172886 478751 172942 478760
rect 172520 472524 172572 472530
rect 172520 472466 172572 472472
rect 171428 470566 172100 470594
rect 171428 467158 171456 470566
rect 171416 467152 171468 467158
rect 171416 467094 171468 467100
rect 171322 459368 171378 459377
rect 171322 459303 171378 459312
rect 172532 459241 172560 472466
rect 172992 470594 173020 480023
rect 173544 472530 173572 480023
rect 173532 472524 173584 472530
rect 173532 472466 173584 472472
rect 172624 470566 173020 470594
rect 172624 461553 172652 470566
rect 172610 461544 172666 461553
rect 172610 461479 172666 461488
rect 173912 459270 173940 480023
rect 174280 475402 174308 480023
rect 174004 475374 174308 475402
rect 173900 459264 173952 459270
rect 172518 459232 172574 459241
rect 173900 459206 173952 459212
rect 174004 459202 174032 475374
rect 174740 470594 174768 480023
rect 175568 472666 175596 480037
rect 176028 474094 176056 480037
rect 176120 480023 176410 480051
rect 176672 480023 176870 480051
rect 177040 480023 177330 480051
rect 176016 474088 176068 474094
rect 176016 474030 176068 474036
rect 175556 472660 175608 472666
rect 175556 472602 175608 472608
rect 176120 470594 176148 480023
rect 174096 470566 174768 470594
rect 175292 470566 176148 470594
rect 174096 466138 174124 470566
rect 174084 466132 174136 466138
rect 174084 466074 174136 466080
rect 175292 463350 175320 470566
rect 176672 467226 176700 480023
rect 177040 470594 177068 480023
rect 177776 476950 177804 480037
rect 178052 480023 178158 480051
rect 178236 480023 178618 480051
rect 178696 480023 179078 480051
rect 177764 476944 177816 476950
rect 177764 476886 177816 476892
rect 176764 470566 177068 470594
rect 176764 469946 176792 470566
rect 176752 469940 176804 469946
rect 176752 469882 176804 469888
rect 176660 467220 176712 467226
rect 176660 467162 176712 467168
rect 175280 463344 175332 463350
rect 175280 463286 175332 463292
rect 178052 459406 178080 480023
rect 178132 475312 178184 475318
rect 178132 475254 178184 475260
rect 178144 460358 178172 475254
rect 178236 468994 178264 480023
rect 178592 477964 178644 477970
rect 178592 477906 178644 477912
rect 178604 470594 178632 477906
rect 178696 475318 178724 480023
rect 178684 475312 178736 475318
rect 178684 475254 178736 475260
rect 179420 475312 179472 475318
rect 179420 475254 179472 475260
rect 178604 470566 178724 470594
rect 178224 468988 178276 468994
rect 178224 468930 178276 468936
rect 178696 468926 178724 470566
rect 178684 468920 178736 468926
rect 178684 468862 178736 468868
rect 178316 462324 178368 462330
rect 178316 462266 178368 462272
rect 178328 461417 178356 462266
rect 178314 461408 178370 461417
rect 178314 461343 178370 461352
rect 178328 461106 178356 461343
rect 178316 461100 178368 461106
rect 178316 461042 178368 461048
rect 179432 460426 179460 475254
rect 179524 461718 179552 480037
rect 179984 478009 180012 480037
rect 180076 480023 180366 480051
rect 180826 480023 181024 480051
rect 179970 478000 180026 478009
rect 179970 477935 180026 477944
rect 180076 475318 180104 480023
rect 180064 475312 180116 475318
rect 180064 475254 180116 475260
rect 180892 475312 180944 475318
rect 180892 475254 180944 475260
rect 180800 475244 180852 475250
rect 180800 475186 180852 475192
rect 179604 468580 179656 468586
rect 179604 468522 179656 468528
rect 179616 461786 179644 468522
rect 179604 461780 179656 461786
rect 179604 461722 179656 461728
rect 179512 461712 179564 461718
rect 179616 461689 179644 461722
rect 179512 461654 179564 461660
rect 179602 461680 179658 461689
rect 179602 461615 179658 461624
rect 179420 460420 179472 460426
rect 179420 460362 179472 460368
rect 178132 460352 178184 460358
rect 178132 460294 178184 460300
rect 178040 459400 178092 459406
rect 178040 459342 178092 459348
rect 180812 459338 180840 475186
rect 180904 463418 180932 475254
rect 180996 463486 181024 480023
rect 181088 480023 181286 480051
rect 181456 480023 181746 480051
rect 182206 480023 182496 480051
rect 181088 475250 181116 480023
rect 181456 475318 181484 480023
rect 181444 475312 181496 475318
rect 181444 475254 181496 475260
rect 182364 475312 182416 475318
rect 182364 475254 182416 475260
rect 181076 475244 181128 475250
rect 181076 475186 181128 475192
rect 182180 475244 182232 475250
rect 182180 475186 182232 475192
rect 180984 463480 181036 463486
rect 180984 463422 181036 463428
rect 180892 463412 180944 463418
rect 180892 463354 180944 463360
rect 182192 461854 182220 475186
rect 182272 475176 182324 475182
rect 182272 475118 182324 475124
rect 182284 465594 182312 475118
rect 182376 466206 182404 475254
rect 182468 466410 182496 480023
rect 182560 475250 182588 480037
rect 182744 480023 183034 480051
rect 183112 480023 183494 480051
rect 183664 480023 183954 480051
rect 182744 475318 182772 480023
rect 182824 478168 182876 478174
rect 182824 478110 182876 478116
rect 182732 475312 182784 475318
rect 182732 475254 182784 475260
rect 182548 475244 182600 475250
rect 182548 475186 182600 475192
rect 182456 466404 182508 466410
rect 182456 466346 182508 466352
rect 182364 466200 182416 466206
rect 182364 466142 182416 466148
rect 182272 465588 182324 465594
rect 182272 465530 182324 465536
rect 182180 461848 182232 461854
rect 182180 461790 182232 461796
rect 182836 460057 182864 478110
rect 183112 475182 183140 480023
rect 183560 475312 183612 475318
rect 183560 475254 183612 475260
rect 183100 475176 183152 475182
rect 183100 475118 183152 475124
rect 183572 466313 183600 475254
rect 183558 466304 183614 466313
rect 183558 466239 183614 466248
rect 183664 465662 183692 480023
rect 184308 475726 184336 480037
rect 184400 480023 184782 480051
rect 184952 480023 185242 480051
rect 185320 480023 185702 480051
rect 185872 480023 186162 480051
rect 184296 475720 184348 475726
rect 184296 475662 184348 475668
rect 184400 475318 184428 480023
rect 184388 475312 184440 475318
rect 184388 475254 184440 475260
rect 183652 465656 183704 465662
rect 183652 465598 183704 465604
rect 184952 460494 184980 480023
rect 185032 475312 185084 475318
rect 185032 475254 185084 475260
rect 185044 463690 185072 475254
rect 185320 470594 185348 480023
rect 185872 475318 185900 480023
rect 186516 478174 186544 480037
rect 186608 480023 186990 480051
rect 187160 480023 187450 480051
rect 186504 478168 186556 478174
rect 186504 478110 186556 478116
rect 185860 475312 185912 475318
rect 185860 475254 185912 475260
rect 185136 470566 185348 470594
rect 185136 467294 185164 470566
rect 185124 467288 185176 467294
rect 185124 467230 185176 467236
rect 186608 466454 186636 480023
rect 187160 470014 187188 480023
rect 187148 470008 187200 470014
rect 187148 469950 187200 469956
rect 187896 468586 187924 480037
rect 187988 480023 188370 480051
rect 188448 480023 188738 480051
rect 187884 468580 187936 468586
rect 187884 468522 187936 468528
rect 187988 467362 188016 480023
rect 187976 467356 188028 467362
rect 187976 467298 188028 467304
rect 188448 466454 188476 480023
rect 189356 480072 189408 480078
rect 189198 480023 189228 480051
rect 189080 480014 189132 480020
rect 186332 466426 186636 466454
rect 187712 466426 188476 466454
rect 185032 463684 185084 463690
rect 185032 463626 185084 463632
rect 186332 463554 186360 466426
rect 186320 463548 186372 463554
rect 186320 463490 186372 463496
rect 184940 460488 184992 460494
rect 184940 460430 184992 460436
rect 182822 460048 182878 460057
rect 182822 459983 182878 459992
rect 187712 459542 187740 466426
rect 189092 460630 189120 480014
rect 189200 479890 189228 480023
rect 196298 480066 196664 480094
rect 189408 480023 189658 480051
rect 189736 480023 190118 480051
rect 190486 480023 190592 480051
rect 189356 480014 189408 480020
rect 189200 479862 189396 479890
rect 189368 476114 189396 479862
rect 189184 476086 189396 476114
rect 189184 460766 189212 476086
rect 189736 466454 189764 480023
rect 190460 471232 190512 471238
rect 190460 471174 190512 471180
rect 189276 466426 189764 466454
rect 189276 462874 189304 466426
rect 190472 463622 190500 471174
rect 190460 463616 190512 463622
rect 190460 463558 190512 463564
rect 190564 462942 190592 480023
rect 190656 480023 190946 480051
rect 191024 480023 191406 480051
rect 191866 480023 191972 480051
rect 190656 471238 190684 480023
rect 190644 471232 190696 471238
rect 190644 471174 190696 471180
rect 191024 466454 191052 480023
rect 191840 471232 191892 471238
rect 191840 471174 191892 471180
rect 190656 466426 191052 466454
rect 190656 466342 190684 466426
rect 190644 466336 190696 466342
rect 190644 466278 190696 466284
rect 190552 462936 190604 462942
rect 190552 462878 190604 462884
rect 189264 462868 189316 462874
rect 189264 462810 189316 462816
rect 191852 461922 191880 471174
rect 191944 466274 191972 480023
rect 192036 480023 192326 480051
rect 192404 480023 192694 480051
rect 192864 480023 193154 480051
rect 193416 480023 193614 480051
rect 193784 480023 194074 480051
rect 194152 480023 194534 480051
rect 191932 466268 191984 466274
rect 191932 466210 191984 466216
rect 192036 466070 192064 480023
rect 192404 466454 192432 480023
rect 192864 471238 192892 480023
rect 193220 471368 193272 471374
rect 193220 471310 193272 471316
rect 192852 471232 192904 471238
rect 192852 471174 192904 471180
rect 192128 466426 192432 466454
rect 192024 466064 192076 466070
rect 192024 466006 192076 466012
rect 192128 465526 192156 466426
rect 192116 465520 192168 465526
rect 192116 465462 192168 465468
rect 191840 461916 191892 461922
rect 191840 461858 191892 461864
rect 190918 461000 190974 461009
rect 190918 460935 190920 460944
rect 190972 460935 190974 460944
rect 190920 460906 190972 460912
rect 189172 460760 189224 460766
rect 189172 460702 189224 460708
rect 189080 460624 189132 460630
rect 189080 460566 189132 460572
rect 187700 459536 187752 459542
rect 187700 459478 187752 459484
rect 193232 459474 193260 471310
rect 193312 471232 193364 471238
rect 193312 471174 193364 471180
rect 193324 460698 193352 471174
rect 193416 462602 193444 480023
rect 193784 471238 193812 480023
rect 193864 478304 193916 478310
rect 193864 478246 193916 478252
rect 193772 471232 193824 471238
rect 193772 471174 193824 471180
rect 193404 462596 193456 462602
rect 193404 462538 193456 462544
rect 193876 460834 193904 478246
rect 194152 471374 194180 480023
rect 194888 477630 194916 480037
rect 194980 480023 195362 480051
rect 194876 477624 194928 477630
rect 194876 477566 194928 477572
rect 194140 471368 194192 471374
rect 194140 471310 194192 471316
rect 194980 466454 195008 480023
rect 195808 477562 195836 480037
rect 195796 477556 195848 477562
rect 195796 477498 195848 477504
rect 194612 466426 195008 466454
rect 193864 460828 193916 460834
rect 193864 460770 193916 460776
rect 193312 460692 193364 460698
rect 193312 460634 193364 460640
rect 193220 459468 193272 459474
rect 193220 459410 193272 459416
rect 180800 459332 180852 459338
rect 180800 459274 180852 459280
rect 172518 459167 172574 459176
rect 173992 459196 174044 459202
rect 173992 459138 174044 459144
rect 171138 459096 171194 459105
rect 171138 459031 171194 459040
rect 164238 458960 164294 458969
rect 164238 458895 164294 458904
rect 138020 458798 138072 458804
rect 161478 458824 161534 458833
rect 80242 458759 80298 458768
rect 194612 458794 194640 466426
rect 161478 458759 161534 458768
rect 194600 458788 194652 458794
rect 194600 458730 194652 458736
rect 66260 458652 66312 458658
rect 66260 458594 66312 458600
rect 163410 374640 163466 374649
rect 163410 374575 163466 374584
rect 165986 374640 166042 374649
rect 165986 374575 165988 374584
rect 163424 374542 163452 374575
rect 166040 374575 166042 374584
rect 165988 374546 166040 374552
rect 163412 374536 163464 374542
rect 93582 374504 93638 374513
rect 93582 374439 93638 374448
rect 103518 374504 103574 374513
rect 103518 374439 103574 374448
rect 116030 374504 116086 374513
rect 116030 374439 116086 374448
rect 143538 374504 143594 374513
rect 143538 374439 143594 374448
rect 146206 374504 146262 374513
rect 146206 374439 146262 374448
rect 153474 374504 153530 374513
rect 153474 374439 153530 374448
rect 156510 374504 156566 374513
rect 156510 374439 156566 374448
rect 158534 374504 158590 374513
rect 158534 374439 158536 374448
rect 93596 374202 93624 374439
rect 93584 374196 93636 374202
rect 93584 374138 93636 374144
rect 103532 374134 103560 374439
rect 103520 374128 103572 374134
rect 103520 374070 103572 374076
rect 116044 374066 116072 374439
rect 143552 374066 143580 374439
rect 146220 374134 146248 374439
rect 153488 374406 153516 374439
rect 153476 374400 153528 374406
rect 153476 374342 153528 374348
rect 156524 374270 156552 374439
rect 158588 374439 158590 374448
rect 160926 374504 160982 374513
rect 163412 374478 163464 374484
rect 160926 374439 160982 374448
rect 158536 374410 158588 374416
rect 160940 374338 160968 374439
rect 160928 374332 160980 374338
rect 160928 374274 160980 374280
rect 156512 374264 156564 374270
rect 148966 374232 149022 374241
rect 156512 374206 156564 374212
rect 148966 374167 148968 374176
rect 149020 374167 149022 374176
rect 148968 374138 149020 374144
rect 146208 374128 146260 374134
rect 146208 374070 146260 374076
rect 116032 374060 116084 374066
rect 116032 374002 116084 374008
rect 143540 374060 143592 374066
rect 143540 374002 143592 374008
rect 107844 373788 107896 373794
rect 107844 373730 107896 373736
rect 136456 373788 136508 373794
rect 136456 373730 136508 373736
rect 100852 373720 100904 373726
rect 100850 373688 100852 373697
rect 107856 373697 107884 373730
rect 131028 373720 131080 373726
rect 100904 373688 100906 373697
rect 100850 373623 100906 373632
rect 107842 373688 107898 373697
rect 107842 373623 107898 373632
rect 113546 373688 113602 373697
rect 113546 373623 113602 373632
rect 118330 373688 118386 373697
rect 118330 373623 118332 373632
rect 113560 373590 113588 373623
rect 118384 373623 118386 373632
rect 121366 373688 121422 373697
rect 121366 373623 121422 373632
rect 125782 373688 125838 373697
rect 125782 373623 125838 373632
rect 128910 373688 128966 373697
rect 128910 373623 128912 373632
rect 118332 373594 118384 373600
rect 113548 373584 113600 373590
rect 105450 373552 105506 373561
rect 105450 373487 105506 373496
rect 110418 373552 110474 373561
rect 113548 373526 113600 373532
rect 110418 373487 110420 373496
rect 105464 373454 105492 373487
rect 110472 373487 110474 373496
rect 110420 373458 110472 373464
rect 121380 373454 121408 373623
rect 125796 373522 125824 373623
rect 128964 373623 128966 373632
rect 131026 373688 131028 373697
rect 136468 373697 136496 373730
rect 131080 373688 131082 373697
rect 131026 373623 131082 373632
rect 133694 373688 133750 373697
rect 133694 373623 133750 373632
rect 136454 373688 136510 373697
rect 136454 373623 136510 373632
rect 139214 373688 139270 373697
rect 139214 373623 139270 373632
rect 141606 373688 141662 373697
rect 141606 373623 141662 373632
rect 151726 373688 151782 373697
rect 151726 373623 151782 373632
rect 128912 373594 128964 373600
rect 133708 373590 133736 373623
rect 133696 373584 133748 373590
rect 133696 373526 133748 373532
rect 125784 373516 125836 373522
rect 125784 373458 125836 373464
rect 105452 373448 105504 373454
rect 88338 373416 88394 373425
rect 88338 373351 88394 373360
rect 96066 373416 96122 373425
rect 96066 373351 96122 373360
rect 98274 373416 98330 373425
rect 105452 373390 105504 373396
rect 121368 373448 121420 373454
rect 121368 373390 121420 373396
rect 122930 373416 122986 373425
rect 98274 373351 98276 373360
rect 88352 373182 88380 373351
rect 96080 373250 96108 373351
rect 98328 373351 98330 373360
rect 99380 373380 99432 373386
rect 98276 373322 98328 373328
rect 122930 373351 122986 373360
rect 99380 373322 99432 373328
rect 96068 373244 96120 373250
rect 96068 373186 96120 373192
rect 88340 373176 88392 373182
rect 88340 373118 88392 373124
rect 90178 373144 90234 373153
rect 90178 373079 90180 373088
rect 90232 373079 90234 373088
rect 92386 373144 92442 373153
rect 92386 373079 92442 373088
rect 90180 373050 90232 373056
rect 60738 372872 60794 372881
rect 60738 372807 60794 372816
rect 60752 353326 60780 372807
rect 77206 372600 77262 372609
rect 77206 372535 77262 372544
rect 81990 372600 82046 372609
rect 81990 372535 82046 372544
rect 84750 372600 84806 372609
rect 84750 372535 84752 372544
rect 77220 372298 77248 372535
rect 78494 372464 78550 372473
rect 78494 372399 78550 372408
rect 79966 372464 80022 372473
rect 79966 372399 80022 372408
rect 80150 372464 80206 372473
rect 80150 372399 80206 372408
rect 77208 372292 77260 372298
rect 77208 372234 77260 372240
rect 78508 372026 78536 372399
rect 78496 372020 78548 372026
rect 78496 371962 78548 371968
rect 77022 371920 77078 371929
rect 77022 371855 77078 371864
rect 77036 369714 77064 371855
rect 78508 371278 78536 371962
rect 79980 371958 80008 372399
rect 79968 371952 80020 371958
rect 79968 371894 80020 371900
rect 79980 371414 80008 371894
rect 80164 371890 80192 372399
rect 80152 371884 80204 371890
rect 80152 371826 80204 371832
rect 79968 371408 80020 371414
rect 79968 371350 80020 371356
rect 80164 371346 80192 371826
rect 82004 371482 82032 372535
rect 84804 372535 84806 372544
rect 86774 372600 86830 372609
rect 86774 372535 86830 372544
rect 88062 372600 88118 372609
rect 88062 372535 88118 372544
rect 89350 372600 89406 372609
rect 89350 372535 89406 372544
rect 90730 372600 90786 372609
rect 90730 372535 90786 372544
rect 92202 372600 92258 372609
rect 92202 372535 92258 372544
rect 84752 372506 84804 372512
rect 86788 372502 86816 372535
rect 86776 372496 86828 372502
rect 85486 372464 85542 372473
rect 86776 372438 86828 372444
rect 85486 372399 85542 372408
rect 85500 371822 85528 372399
rect 85488 371816 85540 371822
rect 85488 371758 85540 371764
rect 88076 371686 88104 372535
rect 89364 372434 89392 372535
rect 89352 372428 89404 372434
rect 89352 372370 89404 372376
rect 88064 371680 88116 371686
rect 88064 371622 88116 371628
rect 90744 371482 90772 372535
rect 92216 372026 92244 372535
rect 92400 372366 92428 373079
rect 93582 372600 93638 372609
rect 93582 372535 93638 372544
rect 92388 372360 92440 372366
rect 92388 372302 92440 372308
rect 93596 372230 93624 372535
rect 99392 372298 99420 373322
rect 122944 373318 122972 373351
rect 122932 373312 122984 373318
rect 122932 373254 122984 373260
rect 139228 373250 139256 373623
rect 139216 373244 139268 373250
rect 139216 373186 139268 373192
rect 141620 373182 141648 373623
rect 141608 373176 141660 373182
rect 141608 373118 141660 373124
rect 151740 373114 151768 373623
rect 191748 373312 191800 373318
rect 191748 373254 191800 373260
rect 151728 373108 151780 373114
rect 151728 373050 151780 373056
rect 102046 372600 102102 372609
rect 102046 372535 102102 372544
rect 112902 372600 112958 372609
rect 112902 372535 112958 372544
rect 114466 372600 114522 372609
rect 114466 372535 114522 372544
rect 99380 372292 99432 372298
rect 99380 372234 99432 372240
rect 93584 372224 93636 372230
rect 93584 372166 93636 372172
rect 92204 372020 92256 372026
rect 92204 371962 92256 371968
rect 95238 371648 95294 371657
rect 95238 371583 95294 371592
rect 99286 371648 99342 371657
rect 99286 371583 99342 371592
rect 100482 371648 100538 371657
rect 100482 371583 100538 371592
rect 81992 371476 82044 371482
rect 81992 371418 82044 371424
rect 90732 371476 90784 371482
rect 90732 371418 90784 371424
rect 80152 371340 80204 371346
rect 80152 371282 80204 371288
rect 78496 371272 78548 371278
rect 78496 371214 78548 371220
rect 95252 369753 95280 371583
rect 97722 371512 97778 371521
rect 97722 371447 97778 371456
rect 95238 369744 95294 369753
rect 77024 369708 77076 369714
rect 95238 369679 95294 369688
rect 77024 369650 77076 369656
rect 97736 369034 97764 371447
rect 99300 369306 99328 371583
rect 99288 369300 99340 369306
rect 99288 369242 99340 369248
rect 100496 369170 100524 371583
rect 101126 371512 101182 371521
rect 101126 371447 101182 371456
rect 100484 369164 100536 369170
rect 100484 369106 100536 369112
rect 97724 369028 97776 369034
rect 97724 368970 97776 368976
rect 101140 368898 101168 371447
rect 102060 371074 102088 372535
rect 104622 372192 104678 372201
rect 104622 372127 104678 372136
rect 102048 371068 102100 371074
rect 102048 371010 102100 371016
rect 104636 369617 104664 372127
rect 112916 371822 112944 372535
rect 114480 372298 114508 372535
rect 114468 372292 114520 372298
rect 114468 372234 114520 372240
rect 105176 371816 105228 371822
rect 105176 371758 105228 371764
rect 112904 371816 112956 371822
rect 112904 371758 112956 371764
rect 104622 369608 104678 369617
rect 104622 369543 104678 369552
rect 105188 368966 105216 371758
rect 106094 371648 106150 371657
rect 106094 371583 106150 371592
rect 182822 371648 182878 371657
rect 182822 371583 182878 371592
rect 183466 371648 183522 371657
rect 183466 371583 183522 371592
rect 106108 369238 106136 371583
rect 107566 371376 107622 371385
rect 107566 371311 107622 371320
rect 106096 369232 106148 369238
rect 106096 369174 106148 369180
rect 105176 368960 105228 368966
rect 105176 368902 105228 368908
rect 101128 368892 101180 368898
rect 101128 368834 101180 368840
rect 107580 367810 107608 371311
rect 182836 371210 182864 371583
rect 182824 371204 182876 371210
rect 182824 371146 182876 371152
rect 107568 367804 107620 367810
rect 107568 367746 107620 367752
rect 182836 360874 182864 371146
rect 183480 371142 183508 371583
rect 183468 371136 183520 371142
rect 183468 371078 183520 371084
rect 183480 370530 183508 371078
rect 183468 370524 183520 370530
rect 183468 370466 183520 370472
rect 182824 360868 182876 360874
rect 182824 360810 182876 360816
rect 179144 356040 179196 356046
rect 179144 355982 179196 355988
rect 179156 355337 179184 355982
rect 191760 355366 191788 373254
rect 196636 370598 196664 480066
rect 196728 370666 196756 480037
rect 196820 480023 197110 480051
rect 197570 480023 197600 480051
rect 196820 370734 196848 480023
rect 197572 479874 197600 480023
rect 197648 480023 198030 480051
rect 198108 480023 198490 480051
rect 197560 479868 197612 479874
rect 197560 479810 197612 479816
rect 197452 478100 197504 478106
rect 197452 478042 197504 478048
rect 197360 478032 197412 478038
rect 197358 478000 197360 478009
rect 197412 478000 197414 478009
rect 197358 477935 197414 477944
rect 197464 477873 197492 478042
rect 197450 477864 197506 477873
rect 197450 477799 197506 477808
rect 196992 477624 197044 477630
rect 196992 477566 197044 477572
rect 196900 477556 196952 477562
rect 196900 477498 196952 477504
rect 196808 370728 196860 370734
rect 196808 370670 196860 370676
rect 196716 370660 196768 370666
rect 196716 370602 196768 370608
rect 196624 370592 196676 370598
rect 196624 370534 196676 370540
rect 196912 370530 196940 477498
rect 195980 370524 196032 370530
rect 195980 370466 196032 370472
rect 196900 370524 196952 370530
rect 196900 370466 196952 370472
rect 195992 368490 196020 370466
rect 197004 370462 197032 477566
rect 197648 476114 197676 480023
rect 198108 476114 198136 480023
rect 198280 479868 198332 479874
rect 198280 479810 198332 479816
rect 198188 478168 198240 478174
rect 198188 478110 198240 478116
rect 197464 476086 197676 476114
rect 197740 476086 198136 476114
rect 197084 465996 197136 466002
rect 197084 465938 197136 465944
rect 197096 374202 197124 465938
rect 197084 374196 197136 374202
rect 197084 374138 197136 374144
rect 197266 373416 197322 373425
rect 197266 373351 197322 373360
rect 196992 370456 197044 370462
rect 196992 370398 197044 370404
rect 195980 368484 196032 368490
rect 195980 368426 196032 368432
rect 196716 368484 196768 368490
rect 196716 368426 196768 368432
rect 191472 355360 191524 355366
rect 179142 355328 179198 355337
rect 179142 355263 179198 355272
rect 191470 355328 191472 355337
rect 191748 355360 191800 355366
rect 191524 355328 191526 355337
rect 191748 355302 191800 355308
rect 191470 355263 191526 355272
rect 179694 354784 179750 354793
rect 179694 354719 179696 354728
rect 179748 354719 179750 354728
rect 179696 354690 179748 354696
rect 60740 353320 60792 353326
rect 60740 353262 60792 353268
rect 107566 269920 107622 269929
rect 107566 269855 107622 269864
rect 110970 269920 111026 269929
rect 110970 269855 111026 269864
rect 107580 269686 107608 269855
rect 108302 269784 108358 269793
rect 108302 269719 108358 269728
rect 60832 269680 60884 269686
rect 107568 269680 107620 269686
rect 60832 269622 60884 269628
rect 83094 269648 83150 269657
rect 60740 269068 60792 269074
rect 60740 269010 60792 269016
rect 60752 268977 60780 269010
rect 60844 269006 60872 269622
rect 83094 269583 83150 269592
rect 93582 269648 93638 269657
rect 93582 269583 93638 269592
rect 94502 269648 94558 269657
rect 107568 269622 107620 269628
rect 94502 269583 94558 269592
rect 60922 269104 60978 269113
rect 60922 269039 60978 269048
rect 76010 269104 76066 269113
rect 76010 269039 76066 269048
rect 77114 269104 77170 269113
rect 77114 269039 77170 269048
rect 60832 269000 60884 269006
rect 60738 268968 60794 268977
rect 60832 268942 60884 268948
rect 60738 268903 60794 268912
rect 60752 249218 60780 268903
rect 60844 249694 60872 268942
rect 60936 268705 60964 269039
rect 61014 268832 61070 268841
rect 61014 268767 61070 268776
rect 60922 268696 60978 268705
rect 60922 268631 60978 268640
rect 60936 249762 60964 268631
rect 60924 249756 60976 249762
rect 60924 249698 60976 249704
rect 60832 249688 60884 249694
rect 60832 249630 60884 249636
rect 61028 249422 61056 268767
rect 76024 268326 76052 269039
rect 77128 268666 77156 269039
rect 83108 268802 83136 269583
rect 90730 269104 90786 269113
rect 90730 269039 90786 269048
rect 83096 268796 83148 268802
rect 83096 268738 83148 268744
rect 77116 268660 77168 268666
rect 77116 268602 77168 268608
rect 90744 268598 90772 269039
rect 90732 268592 90784 268598
rect 90732 268534 90784 268540
rect 93596 268530 93624 269583
rect 93584 268524 93636 268530
rect 93584 268466 93636 268472
rect 76012 268320 76064 268326
rect 76012 268262 76064 268268
rect 64880 268252 64932 268258
rect 64880 268194 64932 268200
rect 62120 268184 62172 268190
rect 62120 268126 62172 268132
rect 62132 266393 62160 268126
rect 64892 267345 64920 268194
rect 94516 268190 94544 269583
rect 108316 269550 108344 269719
rect 108670 269648 108726 269657
rect 110984 269618 111012 269855
rect 133418 269784 133474 269793
rect 133418 269719 133474 269728
rect 135902 269784 135958 269793
rect 135902 269719 135958 269728
rect 138478 269784 138534 269793
rect 138478 269719 138534 269728
rect 108670 269583 108726 269592
rect 110972 269612 111024 269618
rect 108304 269544 108356 269550
rect 108304 269486 108356 269492
rect 95882 269104 95938 269113
rect 95882 269039 95938 269048
rect 96066 269104 96122 269113
rect 96066 269039 96122 269048
rect 98458 269104 98514 269113
rect 98458 269039 98514 269048
rect 99378 269104 99434 269113
rect 99378 269039 99434 269048
rect 95896 268258 95924 269039
rect 96080 268462 96108 269039
rect 96068 268456 96120 268462
rect 96068 268398 96120 268404
rect 98472 268394 98500 269039
rect 98460 268388 98512 268394
rect 98460 268330 98512 268336
rect 95884 268252 95936 268258
rect 95884 268194 95936 268200
rect 94504 268184 94556 268190
rect 85394 268152 85450 268161
rect 92386 268152 92442 268161
rect 85394 268087 85450 268096
rect 86960 268116 87012 268122
rect 82084 268048 82136 268054
rect 82084 267990 82136 267996
rect 64878 267336 64934 267345
rect 64878 267271 64934 267280
rect 77298 266928 77354 266937
rect 77298 266863 77354 266872
rect 80058 266928 80114 266937
rect 80058 266863 80060 266872
rect 77312 266830 77340 266863
rect 80112 266863 80114 266872
rect 80060 266834 80112 266840
rect 77300 266824 77352 266830
rect 77300 266766 77352 266772
rect 62118 266384 62174 266393
rect 62118 266319 62174 266328
rect 63500 266280 63552 266286
rect 63500 266222 63552 266228
rect 63512 264450 63540 266222
rect 78588 265872 78640 265878
rect 78588 265814 78640 265820
rect 63500 264444 63552 264450
rect 63500 264386 63552 264392
rect 78600 264382 78628 265814
rect 78588 264376 78640 264382
rect 78588 264318 78640 264324
rect 82096 264314 82124 267990
rect 84198 267744 84254 267753
rect 84198 267679 84254 267688
rect 84212 266218 84240 267679
rect 84200 266212 84252 266218
rect 84200 266154 84252 266160
rect 85408 266014 85436 268087
rect 94504 268126 94556 268132
rect 92386 268087 92442 268096
rect 86960 268058 87012 268064
rect 86972 267753 87000 268058
rect 86958 267744 87014 267753
rect 86958 267679 87014 267688
rect 88338 267200 88394 267209
rect 88338 267135 88394 267144
rect 88352 266966 88380 267135
rect 88340 266960 88392 266966
rect 88340 266902 88392 266908
rect 91098 266656 91154 266665
rect 91098 266591 91154 266600
rect 85578 266384 85634 266393
rect 85578 266319 85634 266328
rect 88338 266384 88394 266393
rect 88338 266319 88394 266328
rect 89718 266384 89774 266393
rect 89718 266319 89774 266328
rect 85592 266082 85620 266319
rect 85580 266076 85632 266082
rect 85580 266018 85632 266024
rect 85396 266008 85448 266014
rect 85396 265950 85448 265956
rect 88352 265946 88380 266319
rect 89732 266150 89760 266319
rect 89720 266144 89772 266150
rect 89720 266086 89772 266092
rect 88340 265940 88392 265946
rect 88340 265882 88392 265888
rect 91112 265810 91140 266591
rect 92400 266354 92428 268087
rect 99392 267986 99420 269039
rect 103518 268152 103574 268161
rect 103518 268087 103574 268096
rect 99380 267980 99432 267986
rect 99380 267922 99432 267928
rect 102692 267776 102744 267782
rect 102690 267744 102692 267753
rect 102744 267744 102746 267753
rect 102690 267679 102746 267688
rect 100758 267200 100814 267209
rect 100758 267135 100814 267144
rect 100772 267034 100800 267135
rect 103532 267102 103560 268087
rect 108684 268054 108712 269583
rect 110972 269554 111024 269560
rect 133432 269482 133460 269719
rect 133420 269476 133472 269482
rect 133420 269418 133472 269424
rect 135916 269414 135944 269719
rect 135904 269408 135956 269414
rect 135904 269350 135956 269356
rect 138492 269346 138520 269719
rect 140870 269648 140926 269657
rect 140870 269583 140926 269592
rect 143538 269648 143594 269657
rect 143538 269583 143594 269592
rect 145930 269648 145986 269657
rect 145930 269583 145986 269592
rect 138480 269340 138532 269346
rect 138480 269282 138532 269288
rect 140884 269278 140912 269583
rect 140872 269272 140924 269278
rect 140872 269214 140924 269220
rect 143552 269210 143580 269583
rect 143540 269204 143592 269210
rect 143540 269146 143592 269152
rect 145944 269142 145972 269583
rect 145932 269136 145984 269142
rect 145932 269078 145984 269084
rect 196624 269068 196676 269074
rect 196624 269010 196676 269016
rect 128358 268152 128414 268161
rect 128358 268087 128414 268096
rect 153566 268152 153622 268161
rect 153566 268087 153622 268096
rect 108672 268048 108724 268054
rect 108672 267990 108724 267996
rect 113270 268016 113326 268025
rect 113270 267951 113326 267960
rect 105268 267912 105320 267918
rect 105268 267854 105320 267860
rect 105280 267753 105308 267854
rect 106372 267844 106424 267850
rect 106372 267786 106424 267792
rect 106384 267753 106412 267786
rect 105266 267744 105322 267753
rect 105266 267679 105322 267688
rect 106370 267744 106426 267753
rect 106370 267679 106426 267688
rect 113178 267744 113234 267753
rect 113178 267679 113234 267688
rect 113192 267238 113220 267679
rect 113180 267232 113232 267238
rect 104898 267200 104954 267209
rect 113180 267174 113232 267180
rect 104898 267135 104900 267144
rect 104952 267135 104954 267144
rect 104900 267106 104952 267112
rect 103520 267096 103572 267102
rect 103520 267038 103572 267044
rect 100760 267028 100812 267034
rect 100760 266970 100812 266976
rect 100758 266520 100814 266529
rect 100758 266455 100814 266464
rect 92478 266384 92534 266393
rect 92388 266348 92440 266354
rect 92478 266319 92534 266328
rect 96618 266384 96674 266393
rect 96618 266319 96674 266328
rect 97998 266384 98054 266393
rect 97998 266319 98054 266328
rect 92388 266290 92440 266296
rect 92492 266286 92520 266319
rect 92480 266280 92532 266286
rect 92480 266222 92532 266228
rect 91100 265804 91152 265810
rect 91100 265746 91152 265752
rect 82084 264308 82136 264314
rect 82084 264250 82136 264256
rect 96632 264246 96660 266319
rect 96620 264240 96672 264246
rect 96620 264182 96672 264188
rect 82820 250572 82872 250578
rect 82820 250514 82872 250520
rect 67548 250504 67600 250510
rect 67548 250446 67600 250452
rect 61016 249416 61068 249422
rect 61016 249358 61068 249364
rect 60740 249212 60792 249218
rect 60740 249154 60792 249160
rect 67560 249150 67588 250446
rect 67548 249144 67600 249150
rect 67548 249086 67600 249092
rect 82832 249082 82860 250514
rect 98012 250510 98040 266319
rect 100772 265742 100800 266455
rect 100850 266384 100906 266393
rect 100850 266319 100906 266328
rect 111798 266384 111854 266393
rect 111798 266319 111854 266328
rect 100760 265736 100812 265742
rect 100760 265678 100812 265684
rect 100864 250578 100892 266319
rect 111812 265878 111840 266319
rect 111800 265872 111852 265878
rect 111800 265814 111852 265820
rect 113284 265674 113312 267951
rect 117136 267776 117188 267782
rect 117134 267744 117136 267753
rect 117188 267744 117190 267753
rect 117134 267679 117190 267688
rect 122838 267744 122894 267753
rect 122838 267679 122840 267688
rect 122892 267679 122894 267688
rect 122840 267650 122892 267656
rect 125598 267608 125654 267617
rect 128372 267578 128400 268087
rect 129738 267744 129794 267753
rect 129738 267679 129794 267688
rect 129752 267646 129780 267679
rect 153580 267646 153608 268087
rect 196636 267782 196664 269010
rect 196624 267776 196676 267782
rect 155958 267744 156014 267753
rect 155958 267679 156014 267688
rect 158534 267744 158590 267753
rect 158534 267679 158536 267688
rect 129740 267640 129792 267646
rect 129740 267582 129792 267588
rect 153568 267640 153620 267646
rect 153568 267582 153620 267588
rect 155972 267578 156000 267679
rect 158588 267679 158590 267688
rect 163502 267744 163558 267753
rect 196624 267718 196676 267724
rect 163502 267679 163558 267688
rect 158536 267650 158588 267656
rect 125598 267543 125654 267552
rect 128360 267572 128412 267578
rect 125612 267510 125640 267543
rect 128360 267514 128412 267520
rect 155960 267572 156012 267578
rect 155960 267514 156012 267520
rect 163516 267510 163544 267679
rect 125600 267504 125652 267510
rect 117318 267472 117374 267481
rect 117318 267407 117374 267416
rect 120078 267472 120134 267481
rect 163504 267504 163556 267510
rect 125600 267446 125652 267452
rect 160926 267472 160982 267481
rect 120078 267407 120080 267416
rect 117332 267374 117360 267407
rect 120132 267407 120134 267416
rect 163504 267446 163556 267452
rect 166170 267472 166226 267481
rect 160926 267407 160982 267416
rect 166170 267407 166172 267416
rect 120080 267378 120132 267384
rect 160940 267374 160968 267407
rect 166224 267407 166226 267416
rect 183466 267472 183522 267481
rect 183466 267407 183522 267416
rect 166172 267378 166224 267384
rect 117320 267368 117372 267374
rect 115938 267336 115994 267345
rect 117320 267310 117372 267316
rect 160928 267368 160980 267374
rect 160928 267310 160980 267316
rect 183282 267336 183338 267345
rect 115938 267271 115940 267280
rect 115992 267271 115994 267280
rect 183282 267271 183338 267280
rect 115940 267242 115992 267248
rect 183296 267034 183324 267271
rect 183480 267170 183508 267407
rect 183468 267164 183520 267170
rect 183468 267106 183520 267112
rect 183284 267028 183336 267034
rect 183284 266970 183336 266976
rect 147678 266384 147734 266393
rect 147678 266319 147734 266328
rect 113272 265668 113324 265674
rect 113272 265610 113324 265616
rect 147692 264586 147720 266319
rect 147680 264580 147732 264586
rect 147680 264522 147732 264528
rect 180248 250640 180300 250646
rect 180248 250582 180300 250588
rect 100852 250572 100904 250578
rect 100852 250514 100904 250520
rect 98000 250504 98052 250510
rect 98000 250446 98052 250452
rect 179328 250504 179380 250510
rect 179328 250446 179380 250452
rect 179340 249937 179368 250446
rect 180260 249937 180288 250582
rect 179326 249928 179382 249937
rect 179326 249863 179382 249872
rect 180246 249928 180302 249937
rect 180246 249863 180302 249872
rect 190918 249928 190974 249937
rect 190918 249863 190974 249872
rect 190932 249830 190960 249863
rect 190920 249824 190972 249830
rect 190920 249766 190972 249772
rect 82820 249076 82872 249082
rect 82820 249018 82872 249024
rect 96066 164792 96122 164801
rect 96066 164727 96122 164736
rect 140870 164792 140926 164801
rect 140870 164727 140926 164736
rect 96080 164422 96108 164727
rect 103518 164656 103574 164665
rect 103518 164591 103574 164600
rect 105910 164656 105966 164665
rect 105910 164591 105966 164600
rect 117042 164656 117098 164665
rect 117042 164591 117098 164600
rect 96068 164416 96120 164422
rect 96068 164358 96120 164364
rect 98458 164248 98514 164257
rect 98458 164183 98514 164192
rect 101034 164248 101090 164257
rect 101034 164183 101090 164192
rect 98472 164082 98500 164183
rect 98460 164076 98512 164082
rect 98460 164018 98512 164024
rect 101048 164014 101076 164183
rect 101036 164008 101088 164014
rect 101036 163950 101088 163956
rect 103532 163946 103560 164591
rect 103520 163940 103572 163946
rect 103520 163882 103572 163888
rect 105924 163878 105952 164591
rect 108210 164248 108266 164257
rect 108210 164183 108266 164192
rect 105912 163872 105964 163878
rect 105912 163814 105964 163820
rect 108224 163810 108252 164183
rect 117056 163810 117084 164591
rect 140884 164354 140912 164727
rect 153382 164656 153438 164665
rect 153382 164591 153438 164600
rect 163318 164656 163374 164665
rect 163318 164591 163374 164600
rect 140872 164348 140924 164354
rect 140872 164290 140924 164296
rect 145930 164248 145986 164257
rect 145930 164183 145986 164192
rect 148506 164248 148562 164257
rect 148506 164183 148562 164192
rect 150898 164248 150954 164257
rect 150898 164183 150954 164192
rect 108212 163804 108264 163810
rect 108212 163746 108264 163752
rect 116216 163804 116268 163810
rect 116216 163746 116268 163752
rect 117044 163804 117096 163810
rect 117044 163746 117096 163752
rect 60004 163736 60056 163742
rect 60004 163678 60056 163684
rect 59912 163600 59964 163606
rect 59912 163542 59964 163548
rect 99378 163160 99434 163169
rect 99378 163095 99434 163104
rect 113546 163160 113602 163169
rect 113546 163095 113602 163104
rect 73804 162920 73856 162926
rect 73804 162862 73856 162868
rect 60004 160336 60056 160342
rect 60004 160278 60056 160284
rect 59912 146940 59964 146946
rect 59912 146882 59964 146888
rect 59820 146192 59872 146198
rect 59820 146134 59872 146140
rect 59358 140856 59414 140865
rect 59358 140791 59414 140800
rect 59832 59294 59860 146134
rect 59924 145314 59952 146882
rect 59912 145308 59964 145314
rect 59912 145250 59964 145256
rect 59820 59288 59872 59294
rect 59820 59230 59872 59236
rect 59268 57316 59320 57322
rect 59268 57258 59320 57264
rect 59924 56438 59952 145250
rect 59912 56432 59964 56438
rect 59912 56374 59964 56380
rect 59176 56296 59228 56302
rect 59176 56238 59228 56244
rect 60016 56166 60044 160278
rect 73816 146305 73844 162862
rect 75918 162752 75974 162761
rect 75918 162687 75974 162696
rect 77298 162752 77354 162761
rect 77298 162687 77354 162696
rect 78678 162752 78734 162761
rect 78678 162687 78734 162696
rect 80058 162752 80114 162761
rect 80058 162687 80114 162696
rect 81438 162752 81494 162761
rect 81438 162687 81494 162696
rect 82818 162752 82874 162761
rect 82818 162687 82874 162696
rect 84198 162752 84254 162761
rect 84198 162687 84254 162696
rect 85578 162752 85634 162761
rect 85578 162687 85634 162696
rect 86958 162752 87014 162761
rect 86958 162687 87014 162696
rect 88430 162752 88486 162761
rect 88430 162687 88486 162696
rect 89810 162752 89866 162761
rect 89810 162687 89866 162696
rect 90730 162752 90786 162761
rect 90730 162687 90786 162696
rect 91190 162752 91246 162761
rect 91190 162687 91246 162696
rect 92478 162752 92534 162761
rect 92478 162687 92534 162696
rect 93674 162752 93730 162761
rect 93674 162687 93730 162696
rect 93858 162752 93914 162761
rect 93858 162687 93914 162696
rect 95238 162752 95294 162761
rect 95238 162687 95294 162696
rect 96894 162752 96950 162761
rect 96894 162687 96950 162696
rect 97998 162752 98054 162761
rect 97998 162687 98054 162696
rect 73802 146296 73858 146305
rect 73802 146231 73858 146240
rect 75932 145382 75960 162687
rect 76010 162208 76066 162217
rect 76010 162143 76066 162152
rect 76024 145450 76052 162143
rect 77312 145790 77340 162687
rect 78692 148510 78720 162687
rect 80072 148578 80100 162687
rect 81452 148646 81480 162687
rect 81440 148640 81492 148646
rect 81440 148582 81492 148588
rect 80060 148572 80112 148578
rect 80060 148514 80112 148520
rect 78680 148504 78732 148510
rect 78680 148446 78732 148452
rect 77300 145784 77352 145790
rect 77300 145726 77352 145732
rect 82832 145722 82860 162687
rect 82820 145716 82872 145722
rect 82820 145658 82872 145664
rect 84212 145518 84240 162687
rect 84290 161528 84346 161537
rect 84290 161463 84346 161472
rect 84304 145654 84332 161463
rect 85592 145926 85620 162687
rect 86972 146062 87000 162687
rect 88338 162208 88394 162217
rect 88338 162143 88394 162152
rect 88352 162042 88380 162143
rect 88340 162036 88392 162042
rect 88340 161978 88392 161984
rect 87604 161492 87656 161498
rect 87604 161434 87656 161440
rect 86960 146056 87012 146062
rect 87616 146033 87644 161434
rect 86960 145998 87012 146004
rect 87602 146024 87658 146033
rect 88444 145994 88472 162687
rect 87602 145959 87658 145968
rect 88432 145988 88484 145994
rect 88432 145930 88484 145936
rect 85580 145920 85632 145926
rect 85580 145862 85632 145868
rect 89824 145858 89852 162687
rect 90744 162110 90772 162687
rect 91098 162208 91154 162217
rect 91098 162143 91154 162152
rect 90732 162104 90784 162110
rect 90732 162046 90784 162052
rect 89812 145852 89864 145858
rect 89812 145794 89864 145800
rect 84292 145648 84344 145654
rect 84292 145590 84344 145596
rect 91112 145586 91140 162143
rect 91204 146130 91232 162687
rect 91192 146124 91244 146130
rect 91192 146066 91244 146072
rect 92492 145897 92520 162687
rect 93688 162178 93716 162687
rect 93676 162172 93728 162178
rect 93676 162114 93728 162120
rect 93872 146198 93900 162687
rect 95252 161090 95280 162687
rect 96908 161498 96936 162687
rect 96896 161492 96948 161498
rect 96896 161434 96948 161440
rect 95240 161084 95292 161090
rect 95240 161026 95292 161032
rect 98012 161022 98040 162687
rect 98000 161016 98052 161022
rect 98000 160958 98052 160964
rect 99392 146266 99420 163095
rect 100758 162752 100814 162761
rect 100758 162687 100814 162696
rect 102138 162752 102194 162761
rect 102138 162687 102194 162696
rect 103518 162752 103574 162761
rect 103518 162687 103574 162696
rect 104898 162752 104954 162761
rect 104898 162687 104954 162696
rect 106278 162752 106334 162761
rect 106278 162687 106334 162696
rect 107658 162752 107714 162761
rect 107658 162687 107714 162696
rect 109038 162752 109094 162761
rect 109038 162687 109094 162696
rect 110418 162752 110474 162761
rect 110418 162687 110474 162696
rect 111798 162752 111854 162761
rect 111798 162687 111854 162696
rect 99380 146260 99432 146266
rect 99380 146202 99432 146208
rect 93860 146192 93912 146198
rect 93860 146134 93912 146140
rect 92478 145888 92534 145897
rect 92478 145823 92534 145832
rect 100772 145625 100800 162687
rect 100850 162208 100906 162217
rect 100850 162143 100906 162152
rect 100864 146305 100892 162143
rect 100850 146296 100906 146305
rect 100850 146231 100906 146240
rect 102152 145761 102180 162687
rect 103532 147558 103560 162687
rect 104912 147626 104940 162687
rect 106292 161226 106320 162687
rect 106370 162208 106426 162217
rect 106370 162143 106426 162152
rect 106384 161294 106412 162143
rect 106372 161288 106424 161294
rect 106372 161230 106424 161236
rect 106280 161220 106332 161226
rect 106280 161162 106332 161168
rect 104900 147620 104952 147626
rect 104900 147562 104952 147568
rect 103520 147552 103572 147558
rect 103520 147494 103572 147500
rect 107672 146946 107700 162687
rect 109052 160954 109080 162687
rect 109040 160948 109092 160954
rect 109040 160890 109092 160896
rect 110432 160886 110460 162687
rect 110972 162240 111024 162246
rect 110970 162208 110972 162217
rect 111024 162208 111026 162217
rect 110970 162143 111026 162152
rect 110420 160880 110472 160886
rect 110420 160822 110472 160828
rect 111812 160750 111840 162687
rect 113560 162314 113588 163095
rect 114466 162752 114522 162761
rect 114466 162687 114522 162696
rect 114742 162752 114798 162761
rect 114742 162687 114798 162696
rect 115938 162752 115994 162761
rect 115938 162687 115994 162696
rect 113548 162308 113600 162314
rect 113548 162250 113600 162256
rect 114480 161474 114508 162687
rect 114650 162072 114706 162081
rect 114650 162007 114706 162016
rect 114480 161446 114600 161474
rect 111800 160744 111852 160750
rect 111800 160686 111852 160692
rect 114572 149054 114600 161446
rect 114560 149048 114612 149054
rect 114560 148990 114612 148996
rect 114664 148374 114692 162007
rect 114756 161362 114784 162687
rect 115952 162450 115980 162687
rect 115940 162444 115992 162450
rect 115940 162386 115992 162392
rect 114744 161356 114796 161362
rect 114744 161298 114796 161304
rect 116228 148442 116256 163746
rect 145944 163742 145972 164183
rect 145932 163736 145984 163742
rect 145932 163678 145984 163684
rect 148520 163674 148548 164183
rect 148508 163668 148560 163674
rect 148508 163610 148560 163616
rect 150912 163606 150940 164183
rect 150900 163600 150952 163606
rect 150900 163542 150952 163548
rect 153396 163538 153424 164591
rect 163332 164286 163360 164591
rect 163320 164280 163372 164286
rect 163320 164222 163372 164228
rect 196636 163810 196664 267718
rect 196728 267170 196756 368426
rect 197280 356046 197308 373351
rect 197464 370938 197492 476086
rect 197740 471322 197768 476086
rect 197556 471294 197768 471322
rect 197556 371006 197584 471294
rect 197636 468648 197688 468654
rect 197636 468590 197688 468596
rect 197544 371000 197596 371006
rect 197544 370942 197596 370948
rect 197452 370932 197504 370938
rect 197452 370874 197504 370880
rect 197452 360868 197504 360874
rect 197452 360810 197504 360816
rect 197268 356040 197320 356046
rect 197268 355982 197320 355988
rect 197280 354674 197308 355982
rect 197280 354646 197400 354674
rect 196716 267164 196768 267170
rect 196716 267106 196768 267112
rect 196624 163804 196676 163810
rect 196624 163746 196676 163752
rect 153384 163532 153436 163538
rect 153384 163474 153436 163480
rect 196728 163470 196756 267106
rect 197372 250986 197400 354646
rect 197464 267034 197492 360810
rect 197544 354748 197596 354754
rect 197544 354690 197596 354696
rect 197556 267734 197584 354690
rect 197648 269074 197676 468590
rect 198200 466454 198228 478110
rect 198016 466426 198228 466454
rect 197728 460556 197780 460562
rect 197728 460498 197780 460504
rect 197636 269068 197688 269074
rect 197636 269010 197688 269016
rect 197556 267706 197676 267734
rect 197452 267028 197504 267034
rect 197452 266970 197504 266976
rect 197360 250980 197412 250986
rect 197360 250922 197412 250928
rect 196716 163464 196768 163470
rect 196716 163406 196768 163412
rect 197360 163464 197412 163470
rect 197360 163406 197412 163412
rect 128358 163160 128414 163169
rect 128358 163095 128414 163104
rect 117318 162752 117374 162761
rect 117318 162687 117374 162696
rect 118330 162752 118386 162761
rect 118330 162687 118386 162696
rect 118698 162752 118754 162761
rect 118698 162687 118754 162696
rect 120722 162752 120778 162761
rect 120722 162687 120778 162696
rect 122838 162752 122894 162761
rect 122838 162687 122894 162696
rect 125874 162752 125930 162761
rect 128372 162722 128400 163095
rect 133420 162852 133472 162858
rect 133420 162794 133472 162800
rect 130844 162784 130896 162790
rect 130842 162752 130844 162761
rect 133432 162761 133460 162794
rect 130896 162752 130898 162761
rect 125874 162687 125930 162696
rect 128360 162716 128412 162722
rect 117332 161430 117360 162687
rect 118344 162382 118372 162687
rect 118332 162376 118384 162382
rect 118332 162318 118384 162324
rect 117320 161424 117372 161430
rect 117320 161366 117372 161372
rect 118712 160818 118740 162687
rect 120736 162518 120764 162687
rect 122852 162586 122880 162687
rect 125888 162654 125916 162687
rect 130842 162687 130898 162696
rect 133418 162752 133474 162761
rect 133418 162687 133474 162696
rect 183466 162752 183522 162761
rect 183466 162687 183522 162696
rect 128360 162658 128412 162664
rect 125876 162648 125928 162654
rect 125876 162590 125928 162596
rect 122840 162580 122892 162586
rect 122840 162522 122892 162528
rect 120724 162512 120776 162518
rect 120724 162454 120776 162460
rect 183190 162480 183246 162489
rect 183190 162415 183246 162424
rect 183204 162178 183232 162415
rect 183480 162314 183508 162687
rect 197372 162314 197400 163406
rect 183468 162308 183520 162314
rect 183468 162250 183520 162256
rect 197360 162308 197412 162314
rect 197360 162250 197412 162256
rect 183192 162172 183244 162178
rect 183192 162114 183244 162120
rect 118700 160812 118752 160818
rect 118700 160754 118752 160760
rect 116216 148436 116268 148442
rect 116216 148378 116268 148384
rect 114652 148368 114704 148374
rect 114652 148310 114704 148316
rect 107660 146940 107712 146946
rect 107660 146882 107712 146888
rect 179052 146260 179104 146266
rect 179052 146202 179104 146208
rect 102138 145752 102194 145761
rect 102138 145687 102194 145696
rect 100758 145616 100814 145625
rect 91100 145580 91152 145586
rect 100758 145551 100814 145560
rect 91100 145522 91152 145528
rect 84200 145512 84252 145518
rect 84200 145454 84252 145460
rect 76012 145444 76064 145450
rect 76012 145386 76064 145392
rect 75920 145376 75972 145382
rect 75920 145318 75972 145324
rect 179064 144945 179092 146202
rect 179696 146192 179748 146198
rect 179696 146134 179748 146140
rect 179708 144945 179736 146134
rect 191748 145580 191800 145586
rect 191748 145522 191800 145528
rect 191760 145489 191788 145522
rect 191746 145480 191802 145489
rect 191746 145415 191802 145424
rect 179050 144936 179106 144945
rect 179050 144871 179106 144880
rect 179694 144936 179750 144945
rect 179694 144871 179750 144880
rect 77114 59800 77170 59809
rect 77114 59735 77170 59744
rect 83094 59800 83150 59809
rect 83094 59735 83150 59744
rect 99470 59800 99526 59809
rect 99470 59735 99526 59744
rect 113546 59800 113602 59809
rect 113546 59735 113602 59744
rect 120906 59800 120962 59809
rect 120906 59735 120962 59744
rect 77128 59702 77156 59735
rect 77116 59696 77168 59702
rect 77116 59638 77168 59644
rect 83108 59634 83136 59735
rect 94502 59664 94558 59673
rect 83096 59628 83148 59634
rect 94502 59599 94558 59608
rect 83096 59570 83148 59576
rect 84200 59356 84252 59362
rect 84200 59298 84252 59304
rect 84212 58041 84240 59298
rect 94516 59294 94544 59599
rect 99484 59566 99512 59735
rect 102782 59664 102838 59673
rect 102782 59599 102838 59608
rect 113270 59664 113326 59673
rect 113270 59599 113326 59608
rect 99472 59560 99524 59566
rect 99472 59502 99524 59508
rect 95882 59392 95938 59401
rect 95882 59327 95938 59336
rect 98090 59392 98146 59401
rect 98090 59327 98146 59336
rect 100758 59392 100814 59401
rect 100758 59327 100814 59336
rect 101770 59392 101826 59401
rect 101770 59327 101826 59336
rect 94504 59288 94556 59294
rect 94504 59230 94556 59236
rect 95896 59226 95924 59327
rect 95884 59220 95936 59226
rect 95884 59162 95936 59168
rect 98104 59158 98132 59327
rect 98092 59152 98144 59158
rect 98092 59094 98144 59100
rect 100772 59090 100800 59327
rect 100760 59084 100812 59090
rect 100760 59026 100812 59032
rect 101784 58954 101812 59327
rect 102796 59022 102824 59599
rect 102784 59016 102836 59022
rect 102784 58958 102836 58964
rect 101772 58948 101824 58954
rect 101772 58890 101824 58896
rect 113284 58818 113312 59599
rect 113560 59498 113588 59735
rect 116950 59664 117006 59673
rect 116950 59599 117006 59608
rect 113548 59492 113600 59498
rect 113548 59434 113600 59440
rect 116964 58886 116992 59599
rect 120920 59430 120948 59735
rect 120908 59424 120960 59430
rect 120908 59366 120960 59372
rect 148506 59256 148562 59265
rect 148506 59191 148562 59200
rect 150898 59256 150954 59265
rect 150898 59191 150954 59200
rect 116952 58880 117004 58886
rect 116952 58822 117004 58828
rect 113272 58812 113324 58818
rect 113272 58754 113324 58760
rect 148520 58750 148548 59191
rect 148508 58744 148560 58750
rect 148508 58686 148560 58692
rect 150912 58682 150940 59191
rect 150900 58676 150952 58682
rect 150900 58618 150952 58624
rect 84198 58032 84254 58041
rect 84198 57967 84254 57976
rect 76010 57896 76066 57905
rect 76010 57831 76066 57840
rect 78218 57896 78274 57905
rect 78218 57831 78274 57840
rect 79506 57896 79562 57905
rect 79506 57831 79562 57840
rect 80058 57896 80114 57905
rect 80058 57831 80114 57840
rect 81806 57896 81862 57905
rect 81806 57831 81862 57840
rect 85394 57896 85450 57905
rect 85394 57831 85450 57840
rect 86498 57896 86554 57905
rect 86498 57831 86554 57840
rect 86958 57896 87014 57905
rect 86958 57831 87014 57840
rect 88338 57896 88394 57905
rect 88338 57831 88394 57840
rect 88706 57896 88762 57905
rect 88706 57831 88762 57840
rect 89718 57896 89774 57905
rect 89718 57831 89774 57840
rect 90730 57896 90786 57905
rect 90730 57831 90786 57840
rect 91190 57896 91246 57905
rect 91190 57831 91246 57840
rect 92110 57896 92166 57905
rect 92110 57831 92166 57840
rect 92478 57896 92534 57905
rect 92478 57831 92534 57840
rect 103794 57896 103850 57905
rect 103794 57831 103850 57840
rect 104990 57896 105046 57905
rect 104990 57831 105046 57840
rect 106370 57896 106426 57905
rect 106370 57831 106426 57840
rect 106738 57896 106794 57905
rect 106738 57831 106794 57840
rect 108026 57896 108082 57905
rect 108026 57831 108082 57840
rect 109222 57896 109278 57905
rect 109222 57831 109278 57840
rect 111154 57896 111210 57905
rect 111154 57831 111210 57840
rect 115754 57896 115810 57905
rect 115754 57831 115810 57840
rect 123482 57896 123538 57905
rect 123482 57831 123538 57840
rect 125874 57896 125930 57905
rect 125874 57831 125930 57840
rect 128358 57896 128414 57905
rect 128358 57831 128414 57840
rect 130842 57896 130898 57905
rect 130842 57831 130898 57840
rect 133418 57896 133474 57905
rect 133418 57831 133474 57840
rect 145562 57896 145618 57905
rect 145562 57831 145564 57840
rect 76024 57186 76052 57831
rect 78232 57254 78260 57831
rect 78220 57248 78272 57254
rect 78220 57190 78272 57196
rect 76012 57180 76064 57186
rect 76012 57122 76064 57128
rect 60004 56160 60056 56166
rect 60004 56102 60056 56108
rect 79520 55758 79548 57831
rect 79508 55752 79560 55758
rect 79508 55694 79560 55700
rect 58900 54800 58952 54806
rect 58900 54742 58952 54748
rect 80072 54738 80100 57831
rect 81820 56574 81848 57831
rect 81808 56568 81860 56574
rect 81808 56510 81860 56516
rect 85408 55894 85436 57831
rect 86512 55962 86540 57831
rect 86500 55956 86552 55962
rect 86500 55898 86552 55904
rect 85396 55888 85448 55894
rect 85396 55830 85448 55836
rect 86972 54874 87000 57831
rect 88352 57390 88380 57831
rect 88340 57384 88392 57390
rect 88340 57326 88392 57332
rect 88720 56030 88748 57831
rect 88708 56024 88760 56030
rect 88708 55966 88760 55972
rect 86960 54868 87012 54874
rect 86960 54810 87012 54816
rect 89732 54806 89760 57831
rect 90744 57322 90772 57831
rect 90732 57316 90784 57322
rect 90732 57258 90784 57264
rect 91204 54942 91232 57831
rect 92124 56098 92152 57831
rect 92112 56092 92164 56098
rect 92112 56034 92164 56040
rect 92492 55010 92520 57831
rect 103808 56234 103836 57831
rect 105004 56370 105032 57831
rect 104992 56364 105044 56370
rect 104992 56306 105044 56312
rect 103796 56228 103848 56234
rect 103796 56170 103848 56176
rect 106384 56166 106412 57831
rect 106752 56302 106780 57831
rect 108040 56438 108068 57831
rect 109236 56506 109264 57831
rect 111168 57458 111196 57831
rect 111798 57624 111854 57633
rect 111798 57559 111854 57568
rect 113178 57624 113234 57633
rect 113178 57559 113234 57568
rect 111156 57452 111208 57458
rect 111156 57394 111208 57400
rect 109224 56500 109276 56506
rect 109224 56442 109276 56448
rect 108028 56432 108080 56438
rect 108028 56374 108080 56380
rect 106740 56296 106792 56302
rect 106740 56238 106792 56244
rect 106372 56160 106424 56166
rect 106372 56102 106424 56108
rect 111812 55078 111840 57559
rect 113192 55146 113220 57559
rect 115768 55826 115796 57831
rect 123496 57730 123524 57831
rect 123484 57724 123536 57730
rect 123484 57666 123536 57672
rect 115938 57624 115994 57633
rect 115938 57559 115994 57568
rect 118698 57624 118754 57633
rect 118698 57559 118754 57568
rect 115756 55820 115808 55826
rect 115756 55762 115808 55768
rect 115952 55214 115980 57559
rect 115940 55208 115992 55214
rect 115940 55150 115992 55156
rect 113180 55140 113232 55146
rect 113180 55082 113232 55088
rect 111800 55072 111852 55078
rect 111800 55014 111852 55020
rect 92480 55004 92532 55010
rect 92480 54946 92532 54952
rect 91192 54936 91244 54942
rect 91192 54878 91244 54884
rect 89720 54800 89772 54806
rect 118712 54777 118740 57559
rect 125888 57526 125916 57831
rect 128372 57594 128400 57831
rect 130856 57662 130884 57831
rect 133432 57798 133460 57831
rect 145616 57831 145618 57840
rect 153290 57896 153346 57905
rect 153290 57831 153346 57840
rect 183282 57896 183338 57905
rect 183282 57831 183284 57840
rect 145564 57802 145616 57808
rect 133420 57792 133472 57798
rect 133420 57734 133472 57740
rect 130844 57656 130896 57662
rect 130844 57598 130896 57604
rect 128360 57588 128412 57594
rect 128360 57530 128412 57536
rect 125876 57520 125928 57526
rect 125876 57462 125928 57468
rect 153304 56273 153332 57831
rect 183336 57831 183338 57840
rect 183284 57802 183336 57808
rect 197372 57798 197400 162250
rect 197464 162178 197492 266970
rect 197544 250980 197596 250986
rect 197544 250922 197596 250928
rect 197556 250510 197584 250922
rect 197648 250646 197676 267706
rect 197740 267510 197768 460498
rect 197912 459128 197964 459134
rect 197912 459070 197964 459076
rect 197820 458992 197872 458998
rect 197820 458934 197872 458940
rect 197832 373454 197860 458934
rect 197924 374542 197952 459070
rect 197912 374536 197964 374542
rect 197912 374478 197964 374484
rect 197820 373448 197872 373454
rect 197820 373390 197872 373396
rect 198016 268394 198044 466426
rect 198096 390584 198148 390590
rect 198096 390526 198148 390532
rect 198108 373114 198136 390526
rect 198188 389224 198240 389230
rect 198188 389166 198240 389172
rect 198200 373658 198228 389166
rect 198188 373652 198240 373658
rect 198188 373594 198240 373600
rect 198096 373108 198148 373114
rect 198096 373050 198148 373056
rect 198292 370802 198320 479810
rect 198740 471368 198792 471374
rect 198740 471310 198792 471316
rect 198844 471322 198872 480037
rect 199028 480023 199318 480051
rect 199488 480023 199778 480051
rect 199028 471374 199056 480023
rect 199108 479052 199160 479058
rect 199108 478994 199160 479000
rect 199016 471368 199068 471374
rect 198646 375320 198702 375329
rect 198646 375255 198702 375264
rect 198280 370796 198332 370802
rect 198280 370738 198332 370744
rect 198004 268388 198056 268394
rect 198004 268330 198056 268336
rect 197728 267504 197780 267510
rect 197728 267446 197780 267452
rect 197636 250640 197688 250646
rect 197636 250582 197688 250588
rect 197544 250504 197596 250510
rect 197544 250446 197596 250452
rect 197452 162172 197504 162178
rect 197452 162114 197504 162120
rect 197464 57866 197492 162114
rect 197556 146266 197584 250446
rect 197544 146260 197596 146266
rect 197544 146202 197596 146208
rect 197648 146198 197676 250582
rect 198004 173188 198056 173194
rect 198004 173130 198056 173136
rect 197636 146192 197688 146198
rect 197636 146134 197688 146140
rect 198016 145586 198044 173130
rect 198004 145580 198056 145586
rect 198004 145522 198056 145528
rect 198660 58818 198688 375255
rect 198752 371210 198780 471310
rect 198844 471294 198964 471322
rect 199016 471310 199068 471316
rect 198832 471232 198884 471238
rect 198832 471174 198884 471180
rect 198740 371204 198792 371210
rect 198740 371146 198792 371152
rect 198844 370394 198872 471174
rect 198936 371142 198964 471294
rect 199016 460216 199068 460222
rect 199016 460158 199068 460164
rect 199028 458386 199056 460158
rect 199016 458380 199068 458386
rect 199016 458322 199068 458328
rect 199028 454753 199056 458322
rect 199014 454744 199070 454753
rect 199014 454679 199070 454688
rect 198924 371136 198976 371142
rect 198924 371078 198976 371084
rect 198832 370388 198884 370394
rect 198832 370330 198884 370336
rect 199028 349625 199056 454679
rect 199120 390590 199148 478994
rect 199384 475584 199436 475590
rect 199384 475526 199436 475532
rect 199200 475244 199252 475250
rect 199200 475186 199252 475192
rect 199212 390930 199240 475186
rect 199396 466454 199424 475526
rect 199488 471238 199516 480023
rect 200224 478242 200252 480037
rect 200408 480023 200698 480051
rect 200212 478236 200264 478242
rect 200212 478178 200264 478184
rect 199476 471232 199528 471238
rect 199476 471174 199528 471180
rect 200408 466454 200436 480023
rect 200764 478576 200816 478582
rect 200762 478544 200764 478553
rect 200816 478544 200818 478553
rect 200762 478479 200818 478488
rect 200488 478372 200540 478378
rect 200488 478314 200540 478320
rect 200500 477601 200528 478314
rect 200486 477592 200542 477601
rect 200486 477527 200542 477536
rect 200488 475652 200540 475658
rect 200488 475594 200540 475600
rect 199396 466426 199516 466454
rect 199384 462868 199436 462874
rect 199384 462810 199436 462816
rect 199292 458924 199344 458930
rect 199292 458866 199344 458872
rect 199200 390924 199252 390930
rect 199200 390866 199252 390872
rect 199198 390824 199254 390833
rect 199198 390759 199254 390768
rect 199108 390584 199160 390590
rect 199108 390526 199160 390532
rect 199212 373994 199240 390759
rect 199120 373966 199240 373994
rect 199120 373862 199148 373966
rect 199108 373856 199160 373862
rect 199108 373798 199160 373804
rect 199120 370682 199148 373798
rect 199304 373726 199332 458866
rect 199396 374202 199424 462810
rect 199488 389230 199516 466426
rect 200224 466426 200436 466454
rect 199568 459060 199620 459066
rect 199568 459002 199620 459008
rect 199476 389224 199528 389230
rect 199476 389166 199528 389172
rect 199474 389056 199530 389065
rect 199474 388991 199530 389000
rect 199384 374196 199436 374202
rect 199384 374138 199436 374144
rect 199488 373969 199516 388991
rect 199580 374610 199608 459002
rect 199658 393816 199714 393825
rect 199658 393751 199714 393760
rect 199672 393378 199700 393751
rect 199660 393372 199712 393378
rect 199660 393314 199712 393320
rect 199844 390924 199896 390930
rect 199844 390866 199896 390872
rect 199856 388521 199884 390866
rect 199842 388512 199898 388521
rect 199842 388447 199898 388456
rect 199568 374604 199620 374610
rect 199568 374546 199620 374552
rect 199474 373960 199530 373969
rect 199530 373918 199608 373946
rect 199474 373895 199530 373904
rect 199292 373720 199344 373726
rect 199292 373662 199344 373668
rect 199120 370654 199516 370682
rect 199384 365696 199436 365702
rect 199384 365638 199436 365644
rect 199396 365022 199424 365638
rect 199384 365016 199436 365022
rect 199384 364958 199436 364964
rect 198738 349616 198794 349625
rect 198738 349551 198794 349560
rect 199014 349616 199070 349625
rect 199014 349551 199070 349560
rect 198752 244225 198780 349551
rect 198830 289776 198886 289785
rect 198830 289711 198886 289720
rect 198738 244216 198794 244225
rect 198738 244151 198794 244160
rect 198844 184385 198872 289711
rect 199396 287054 199424 364958
rect 199488 359514 199516 370654
rect 199580 365702 199608 373918
rect 199568 365696 199620 365702
rect 199568 365638 199620 365644
rect 199660 362228 199712 362234
rect 199660 362170 199712 362176
rect 199476 359508 199528 359514
rect 199476 359450 199528 359456
rect 199028 287026 199424 287054
rect 199028 284889 199056 287026
rect 199488 286385 199516 359450
rect 199568 356720 199620 356726
rect 199568 356662 199620 356668
rect 199474 286376 199530 286385
rect 199474 286311 199530 286320
rect 199014 284880 199070 284889
rect 199014 284815 199070 284824
rect 198922 283112 198978 283121
rect 198922 283047 198978 283056
rect 198830 184376 198886 184385
rect 198830 184311 198886 184320
rect 198936 180794 198964 283047
rect 198844 180766 198964 180794
rect 198738 179480 198794 179489
rect 198738 179415 198794 179424
rect 198752 74905 198780 179415
rect 198844 178673 198872 180766
rect 199028 179489 199056 284815
rect 199488 283642 199516 286311
rect 199212 283614 199516 283642
rect 199212 277394 199240 283614
rect 199580 283121 199608 356662
rect 199672 289785 199700 362170
rect 199750 358048 199806 358057
rect 199750 357983 199806 357992
rect 199658 289776 199714 289785
rect 199658 289711 199714 289720
rect 199764 287745 199792 357983
rect 199856 356726 199884 388447
rect 200224 374814 200252 466426
rect 200396 463072 200448 463078
rect 200396 463014 200448 463020
rect 200304 463004 200356 463010
rect 200304 462946 200356 462952
rect 200212 374808 200264 374814
rect 200212 374750 200264 374756
rect 200026 373280 200082 373289
rect 200026 373215 200082 373224
rect 200040 362234 200068 373215
rect 200028 362228 200080 362234
rect 200028 362170 200080 362176
rect 199844 356720 199896 356726
rect 199844 356662 199896 356668
rect 199750 287736 199806 287745
rect 199750 287671 199806 287680
rect 199566 283112 199622 283121
rect 199566 283047 199622 283056
rect 199764 277394 199792 287671
rect 199120 277366 199240 277394
rect 199304 277366 199792 277394
rect 199120 181393 199148 277366
rect 199198 244216 199254 244225
rect 199198 244151 199254 244160
rect 199106 181384 199162 181393
rect 199106 181319 199162 181328
rect 199014 179480 199070 179489
rect 199014 179415 199070 179424
rect 198830 178664 198886 178673
rect 198830 178599 198886 178608
rect 198738 74896 198794 74905
rect 198738 74831 198794 74840
rect 198844 73681 198872 178599
rect 199120 76401 199148 181319
rect 199212 139233 199240 244151
rect 199304 182753 199332 277366
rect 200316 267646 200344 462946
rect 200304 267640 200356 267646
rect 200304 267582 200356 267588
rect 200408 267442 200436 463014
rect 200500 373794 200528 475594
rect 200764 467356 200816 467362
rect 200764 467298 200816 467304
rect 200580 465928 200632 465934
rect 200580 465870 200632 465876
rect 200592 374406 200620 465870
rect 200672 458856 200724 458862
rect 200672 458798 200724 458804
rect 200580 374400 200632 374406
rect 200580 374342 200632 374348
rect 200488 373788 200540 373794
rect 200488 373730 200540 373736
rect 200684 373250 200712 458798
rect 200672 373244 200724 373250
rect 200672 373186 200724 373192
rect 200396 267436 200448 267442
rect 200396 267378 200448 267384
rect 200776 266801 200804 467298
rect 200856 466132 200908 466138
rect 200856 466074 200908 466080
rect 200868 269550 200896 466074
rect 200948 459536 201000 459542
rect 200948 459478 201000 459484
rect 200960 280158 200988 459478
rect 201052 374746 201080 480037
rect 201406 375320 201462 375329
rect 201406 375255 201462 375264
rect 201040 374740 201092 374746
rect 201040 374682 201092 374688
rect 200948 280152 201000 280158
rect 200948 280094 201000 280100
rect 200856 269544 200908 269550
rect 200856 269486 200908 269492
rect 200762 266792 200818 266801
rect 200762 266727 200818 266736
rect 199382 184376 199438 184385
rect 199382 184311 199438 184320
rect 199290 182744 199346 182753
rect 199290 182679 199346 182688
rect 199198 139224 199254 139233
rect 199198 139159 199254 139168
rect 199304 77761 199332 182679
rect 199396 79393 199424 184311
rect 199382 79384 199438 79393
rect 199382 79319 199438 79328
rect 199290 77752 199346 77761
rect 199290 77687 199346 77696
rect 199106 76392 199162 76401
rect 199106 76327 199162 76336
rect 198830 73672 198886 73681
rect 198830 73607 198886 73616
rect 201420 58886 201448 375255
rect 201512 374882 201540 480037
rect 201592 478508 201644 478514
rect 201592 478450 201644 478456
rect 201604 478417 201632 478450
rect 201590 478408 201646 478417
rect 201590 478343 201646 478352
rect 201972 478174 202000 480037
rect 201960 478168 202012 478174
rect 201960 478110 202012 478116
rect 202432 477630 202460 480037
rect 202906 480023 203104 480051
rect 202420 477624 202472 477630
rect 202420 477566 202472 477572
rect 201684 475516 201736 475522
rect 201684 475458 201736 475464
rect 201592 461780 201644 461786
rect 201592 461722 201644 461728
rect 201604 461038 201632 461722
rect 201592 461032 201644 461038
rect 201592 460974 201644 460980
rect 201500 374876 201552 374882
rect 201500 374818 201552 374824
rect 201604 354754 201632 460974
rect 201696 373522 201724 475458
rect 202880 471232 202932 471238
rect 202880 471174 202932 471180
rect 202328 468988 202380 468994
rect 202328 468930 202380 468936
rect 201776 465860 201828 465866
rect 201776 465802 201828 465808
rect 201788 374474 201816 465802
rect 202144 463208 202196 463214
rect 202144 463150 202196 463156
rect 201776 374468 201828 374474
rect 201776 374410 201828 374416
rect 201684 373516 201736 373522
rect 201684 373458 201736 373464
rect 201592 354748 201644 354754
rect 201592 354690 201644 354696
rect 202156 162110 202184 463150
rect 202234 459368 202290 459377
rect 202234 459303 202290 459312
rect 202248 164286 202276 459303
rect 202340 267510 202368 468930
rect 202420 465588 202472 465594
rect 202420 465530 202472 465536
rect 202432 268598 202460 465530
rect 202512 462596 202564 462602
rect 202512 462538 202564 462544
rect 202524 369782 202552 462538
rect 202604 460760 202656 460766
rect 202604 460702 202656 460708
rect 202616 383586 202644 460702
rect 202604 383580 202656 383586
rect 202604 383522 202656 383528
rect 202892 369850 202920 471174
rect 202972 465724 203024 465730
rect 202972 465666 203024 465672
rect 202880 369844 202932 369850
rect 202880 369786 202932 369792
rect 202512 369776 202564 369782
rect 202512 369718 202564 369724
rect 202420 268592 202472 268598
rect 202420 268534 202472 268540
rect 202984 267578 203012 465666
rect 203076 374678 203104 480023
rect 203168 480023 203274 480051
rect 203352 480023 203734 480051
rect 203904 480023 204194 480051
rect 204272 480023 204654 480051
rect 203168 471238 203196 480023
rect 203156 471232 203208 471238
rect 203156 471174 203208 471180
rect 203156 471096 203208 471102
rect 203156 471038 203208 471044
rect 203064 374672 203116 374678
rect 203064 374614 203116 374620
rect 203168 374542 203196 471038
rect 203352 466454 203380 480023
rect 203904 471102 203932 480023
rect 203892 471096 203944 471102
rect 203892 471038 203944 471044
rect 203260 466426 203380 466454
rect 203260 413982 203288 466426
rect 203524 464364 203576 464370
rect 203524 464306 203576 464312
rect 203340 460828 203392 460834
rect 203340 460770 203392 460776
rect 203248 413976 203300 413982
rect 203248 413918 203300 413924
rect 203248 393372 203300 393378
rect 203248 393314 203300 393320
rect 203156 374536 203208 374542
rect 203156 374478 203208 374484
rect 203168 369714 203196 374478
rect 203260 373289 203288 393314
rect 203246 373280 203302 373289
rect 203246 373215 203302 373224
rect 203352 373182 203380 460770
rect 203340 373176 203392 373182
rect 203340 373118 203392 373124
rect 203156 369708 203208 369714
rect 203156 369650 203208 369656
rect 202972 267572 203024 267578
rect 202972 267514 203024 267520
rect 202328 267504 202380 267510
rect 202328 267446 202380 267452
rect 203536 173806 203564 464306
rect 203800 462936 203852 462942
rect 203800 462878 203852 462884
rect 203616 461848 203668 461854
rect 203616 461790 203668 461796
rect 203628 268734 203656 461790
rect 203708 459400 203760 459406
rect 203708 459342 203760 459348
rect 203616 268728 203668 268734
rect 203616 268670 203668 268676
rect 203720 267442 203748 459342
rect 203812 369374 203840 462878
rect 204272 373658 204300 480023
rect 204444 475448 204496 475454
rect 204444 475390 204496 475396
rect 204352 471232 204404 471238
rect 204352 471174 204404 471180
rect 204364 405006 204392 471174
rect 204352 405000 204404 405006
rect 204352 404942 204404 404948
rect 204260 373652 204312 373658
rect 204260 373594 204312 373600
rect 204272 373386 204300 373594
rect 204456 373590 204484 475390
rect 205008 474162 205036 480037
rect 205192 480023 205482 480051
rect 205744 480023 205942 480051
rect 206020 480023 206402 480051
rect 206480 480023 206862 480051
rect 207230 480023 207336 480051
rect 204996 474156 205048 474162
rect 204996 474098 205048 474104
rect 205192 471238 205220 480023
rect 205640 478644 205692 478650
rect 205640 478586 205692 478592
rect 205652 478553 205680 478586
rect 205638 478544 205694 478553
rect 205638 478479 205694 478488
rect 205640 478440 205692 478446
rect 205640 478382 205692 478388
rect 205652 477737 205680 478382
rect 205638 477728 205694 477737
rect 205638 477663 205694 477672
rect 205744 475538 205772 480023
rect 206020 475538 206048 480023
rect 206100 478984 206152 478990
rect 206100 478926 206152 478932
rect 205652 475510 205772 475538
rect 205836 475510 206048 475538
rect 205652 475182 205680 475510
rect 205732 475380 205784 475386
rect 205732 475322 205784 475328
rect 205640 475176 205692 475182
rect 205640 475118 205692 475124
rect 205180 471232 205232 471238
rect 205180 471174 205232 471180
rect 204996 469940 205048 469946
rect 204996 469882 205048 469888
rect 204902 466168 204958 466177
rect 204902 466103 204958 466112
rect 204536 465792 204588 465798
rect 204536 465734 204588 465740
rect 204548 374270 204576 465734
rect 204536 374264 204588 374270
rect 204536 374206 204588 374212
rect 204444 373584 204496 373590
rect 204444 373526 204496 373532
rect 204260 373380 204312 373386
rect 204260 373322 204312 373328
rect 203800 369368 203852 369374
rect 203800 369310 203852 369316
rect 203708 267436 203760 267442
rect 203708 267378 203760 267384
rect 203524 173800 203576 173806
rect 203524 173742 203576 173748
rect 202236 164280 202288 164286
rect 202236 164222 202288 164228
rect 204916 162790 204944 466103
rect 205008 267306 205036 469882
rect 205086 466032 205142 466041
rect 205086 465967 205142 465976
rect 204996 267300 205048 267306
rect 204996 267242 205048 267248
rect 205100 164354 205128 465967
rect 205180 465656 205232 465662
rect 205180 465598 205232 465604
rect 205192 268530 205220 465598
rect 205364 461916 205416 461922
rect 205364 461858 205416 461864
rect 205272 459264 205324 459270
rect 205272 459206 205324 459212
rect 205284 278730 205312 459206
rect 205376 369442 205404 461858
rect 205744 409154 205772 475322
rect 205836 457502 205864 475510
rect 205916 475176 205968 475182
rect 205916 475118 205968 475124
rect 205928 469946 205956 475118
rect 206112 470594 206140 478926
rect 206376 477896 206428 477902
rect 206376 477838 206428 477844
rect 206020 470566 206140 470594
rect 205916 469940 205968 469946
rect 205916 469882 205968 469888
rect 205916 468920 205968 468926
rect 205916 468862 205968 468868
rect 205824 457496 205876 457502
rect 205824 457438 205876 457444
rect 205732 409148 205784 409154
rect 205732 409090 205784 409096
rect 205546 375320 205602 375329
rect 205546 375255 205602 375264
rect 205364 369436 205416 369442
rect 205364 369378 205416 369384
rect 205272 278724 205324 278730
rect 205272 278666 205324 278672
rect 205180 268524 205232 268530
rect 205180 268466 205232 268472
rect 205088 164348 205140 164354
rect 205088 164290 205140 164296
rect 204904 162784 204956 162790
rect 204904 162726 204956 162732
rect 202144 162104 202196 162110
rect 202144 162046 202196 162052
rect 204904 145580 204956 145586
rect 204904 145522 204956 145528
rect 204916 67658 204944 145522
rect 204904 67652 204956 67658
rect 204904 67594 204956 67600
rect 201408 58880 201460 58886
rect 201408 58822 201460 58828
rect 198648 58812 198700 58818
rect 198648 58754 198700 58760
rect 204916 57934 204944 67594
rect 204904 57928 204956 57934
rect 204904 57870 204956 57876
rect 197452 57860 197504 57866
rect 197452 57802 197504 57808
rect 205560 57798 205588 375255
rect 205928 374066 205956 468862
rect 205916 374060 205968 374066
rect 205916 374002 205968 374008
rect 206020 267714 206048 470566
rect 206192 458788 206244 458794
rect 206192 458730 206244 458736
rect 206204 369714 206232 458730
rect 206284 413976 206336 413982
rect 206284 413918 206336 413924
rect 206296 385014 206324 413918
rect 206284 385008 206336 385014
rect 206284 384950 206336 384956
rect 206284 382288 206336 382294
rect 206284 382230 206336 382236
rect 206296 373318 206324 382230
rect 206284 373312 206336 373318
rect 206284 373254 206336 373260
rect 206192 369708 206244 369714
rect 206192 369650 206244 369656
rect 206008 267708 206060 267714
rect 206008 267650 206060 267656
rect 206388 163538 206416 477838
rect 206480 475386 206508 480023
rect 207112 478916 207164 478922
rect 207112 478858 207164 478864
rect 206468 475380 206520 475386
rect 206468 475322 206520 475328
rect 206560 466404 206612 466410
rect 206560 466346 206612 466352
rect 206466 465896 206522 465905
rect 206466 465831 206522 465840
rect 206376 163532 206428 163538
rect 206376 163474 206428 163480
rect 206480 162382 206508 465831
rect 206572 268870 206600 466346
rect 206652 463344 206704 463350
rect 206652 463286 206704 463292
rect 206560 268864 206612 268870
rect 206560 268806 206612 268812
rect 206664 267102 206692 463286
rect 206744 461712 206796 461718
rect 206744 461654 206796 461660
rect 206756 267578 206784 461654
rect 207020 460964 207072 460970
rect 207020 460906 207072 460912
rect 206926 408640 206982 408649
rect 206926 408575 206982 408584
rect 206834 374640 206890 374649
rect 206834 374575 206890 374584
rect 206744 267572 206796 267578
rect 206744 267514 206796 267520
rect 206652 267096 206704 267102
rect 206652 267038 206704 267044
rect 206468 162376 206520 162382
rect 206468 162318 206520 162324
rect 206848 58750 206876 374575
rect 206940 59022 206968 408575
rect 207032 383654 207060 460906
rect 207020 383648 207072 383654
rect 207020 383590 207072 383596
rect 207032 382294 207060 383590
rect 207020 382288 207072 382294
rect 207020 382230 207072 382236
rect 207124 267374 207152 478858
rect 207204 475380 207256 475386
rect 207204 475322 207256 475328
rect 207216 373833 207244 475322
rect 207308 467362 207336 480023
rect 207400 480023 207690 480051
rect 207768 480023 208150 480051
rect 207296 467356 207348 467362
rect 207296 467298 207348 467304
rect 207400 458250 207428 480023
rect 207768 475386 207796 480023
rect 208400 478848 208452 478854
rect 208400 478790 208452 478796
rect 208412 478009 208440 478790
rect 208398 478000 208454 478009
rect 208398 477935 208454 477944
rect 208596 477562 208624 480037
rect 208688 480023 209070 480051
rect 208584 477556 208636 477562
rect 208584 477498 208636 477504
rect 207756 475380 207808 475386
rect 207756 475322 207808 475328
rect 207664 471300 207716 471306
rect 207664 471242 207716 471248
rect 207480 468716 207532 468722
rect 207480 468658 207532 468664
rect 207388 458244 207440 458250
rect 207388 458186 207440 458192
rect 207492 374134 207520 468658
rect 207480 374128 207532 374134
rect 207480 374070 207532 374076
rect 207202 373824 207258 373833
rect 207202 373759 207258 373768
rect 207216 373182 207244 373759
rect 207204 373176 207256 373182
rect 207204 373118 207256 373124
rect 207112 267368 207164 267374
rect 207112 267310 207164 267316
rect 207676 162722 207704 471242
rect 208688 470594 208716 480023
rect 209424 478378 209452 480037
rect 209412 478372 209464 478378
rect 209412 478314 209464 478320
rect 209596 478304 209648 478310
rect 209596 478246 209648 478252
rect 209504 477624 209556 477630
rect 209504 477566 209556 477572
rect 208412 470566 208716 470594
rect 207848 467220 207900 467226
rect 207848 467162 207900 467168
rect 207754 459232 207810 459241
rect 207754 459167 207810 459176
rect 207768 175234 207796 459167
rect 207860 267238 207888 467162
rect 207940 466200 207992 466206
rect 207940 466142 207992 466148
rect 207952 268802 207980 466142
rect 208032 465520 208084 465526
rect 208032 465462 208084 465468
rect 208044 369578 208072 465462
rect 208124 458244 208176 458250
rect 208124 458186 208176 458192
rect 208136 417450 208164 458186
rect 208124 417444 208176 417450
rect 208124 417386 208176 417392
rect 208216 384328 208268 384334
rect 208216 384270 208268 384276
rect 208228 372502 208256 384270
rect 208306 382392 208362 382401
rect 208306 382327 208362 382336
rect 208216 372496 208268 372502
rect 208216 372438 208268 372444
rect 208122 372328 208178 372337
rect 208122 372263 208178 372272
rect 208032 369572 208084 369578
rect 208032 369514 208084 369520
rect 207940 268796 207992 268802
rect 207940 268738 207992 268744
rect 207848 267232 207900 267238
rect 207848 267174 207900 267180
rect 208136 264314 208164 372263
rect 208228 372026 208256 372438
rect 208216 372020 208268 372026
rect 208216 371962 208268 371968
rect 208124 264308 208176 264314
rect 208124 264250 208176 264256
rect 207756 175228 207808 175234
rect 207756 175170 207808 175176
rect 207664 162716 207716 162722
rect 207664 162658 207716 162664
rect 206928 59016 206980 59022
rect 206928 58958 206980 58964
rect 206836 58744 206888 58750
rect 206836 58686 206888 58692
rect 208320 57934 208348 382327
rect 208412 372570 208440 470566
rect 209228 470008 209280 470014
rect 209228 469950 209280 469956
rect 209044 467152 209096 467158
rect 209044 467094 209096 467100
rect 208492 463140 208544 463146
rect 208492 463082 208544 463088
rect 208504 374338 208532 463082
rect 208860 460692 208912 460698
rect 208860 460634 208912 460640
rect 208492 374332 208544 374338
rect 208492 374274 208544 374280
rect 208400 372564 208452 372570
rect 208400 372506 208452 372512
rect 208768 371884 208820 371890
rect 208768 371826 208820 371832
rect 208780 371482 208808 371826
rect 208768 371476 208820 371482
rect 208768 371418 208820 371424
rect 208872 369510 208900 460634
rect 208952 371748 209004 371754
rect 208952 371690 209004 371696
rect 208964 371482 208992 371690
rect 208952 371476 209004 371482
rect 208952 371418 209004 371424
rect 208860 369504 208912 369510
rect 208860 369446 208912 369452
rect 208964 265577 208992 371418
rect 208950 265568 209006 265577
rect 208950 265503 209006 265512
rect 209056 162858 209084 467094
rect 209136 463276 209188 463282
rect 209136 463218 209188 463224
rect 209148 163674 209176 463218
rect 209240 267481 209268 469950
rect 209412 468580 209464 468586
rect 209412 468522 209464 468528
rect 209320 459332 209372 459338
rect 209320 459274 209372 459280
rect 209332 269142 209360 459274
rect 209320 269136 209372 269142
rect 209320 269078 209372 269084
rect 209424 267617 209452 468522
rect 209516 374474 209544 477566
rect 209504 374468 209556 374474
rect 209504 374410 209556 374416
rect 209608 373561 209636 478246
rect 209780 475380 209832 475386
rect 209780 475322 209832 475328
rect 209686 374640 209742 374649
rect 209686 374575 209742 374584
rect 209594 373552 209650 373561
rect 209594 373487 209650 373496
rect 209502 372192 209558 372201
rect 209502 372127 209558 372136
rect 209516 371521 209544 372127
rect 209594 371920 209650 371929
rect 209594 371855 209650 371864
rect 209608 371657 209636 371855
rect 209594 371648 209650 371657
rect 209594 371583 209650 371592
rect 209502 371512 209558 371521
rect 209502 371447 209558 371456
rect 209410 267608 209466 267617
rect 209410 267543 209466 267552
rect 209226 267472 209282 267481
rect 209226 267407 209282 267416
rect 209516 264246 209544 371447
rect 209504 264240 209556 264246
rect 209504 264182 209556 264188
rect 209608 250578 209636 371583
rect 209596 250572 209648 250578
rect 209596 250514 209648 250520
rect 209136 163668 209188 163674
rect 209136 163610 209188 163616
rect 209044 162852 209096 162858
rect 209044 162794 209096 162800
rect 208308 57928 208360 57934
rect 208308 57870 208360 57876
rect 183468 57792 183520 57798
rect 183466 57760 183468 57769
rect 197360 57792 197412 57798
rect 183520 57760 183522 57769
rect 197360 57734 197412 57740
rect 205548 57792 205600 57798
rect 205548 57734 205600 57740
rect 183466 57695 183522 57704
rect 155958 57624 156014 57633
rect 155958 57559 156014 57568
rect 160098 57624 160154 57633
rect 160098 57559 160154 57568
rect 165618 57624 165674 57633
rect 209700 57594 209728 374575
rect 209792 372434 209820 475322
rect 209780 372428 209832 372434
rect 209780 372370 209832 372376
rect 209884 371686 209912 480037
rect 209976 480023 210358 480051
rect 210436 480023 210818 480051
rect 209976 475386 210004 480023
rect 210240 478780 210292 478786
rect 210240 478722 210292 478728
rect 210252 478281 210280 478722
rect 210238 478272 210294 478281
rect 210238 478207 210294 478216
rect 209964 475380 210016 475386
rect 209964 475322 210016 475328
rect 210436 470594 210464 480023
rect 211172 477562 211200 480037
rect 211264 480023 211646 480051
rect 211816 480023 212106 480051
rect 210792 477556 210844 477562
rect 210792 477498 210844 477504
rect 211160 477556 211212 477562
rect 211160 477498 211212 477504
rect 210608 474088 210660 474094
rect 210608 474030 210660 474036
rect 209976 470566 210464 470594
rect 209976 371890 210004 470566
rect 210424 468852 210476 468858
rect 210424 468794 210476 468800
rect 210056 461100 210108 461106
rect 210056 461042 210108 461048
rect 210068 460970 210096 461042
rect 210056 460964 210108 460970
rect 210056 460906 210108 460912
rect 210068 373425 210096 460906
rect 210332 460624 210384 460630
rect 210332 460566 210384 460572
rect 210240 374400 210292 374406
rect 210240 374342 210292 374348
rect 210148 373448 210200 373454
rect 210054 373416 210110 373425
rect 210148 373390 210200 373396
rect 210054 373351 210110 373360
rect 210056 372428 210108 372434
rect 210056 372370 210108 372376
rect 209964 371884 210016 371890
rect 209964 371826 210016 371832
rect 210068 371822 210096 372370
rect 210056 371816 210108 371822
rect 210056 371758 210108 371764
rect 209872 371680 209924 371686
rect 209872 371622 209924 371628
rect 210056 371408 210108 371414
rect 210056 371350 210108 371356
rect 210068 370870 210096 371350
rect 210056 370864 210108 370870
rect 210056 370806 210108 370812
rect 210160 369034 210188 373390
rect 210148 369028 210200 369034
rect 210148 368970 210200 368976
rect 210252 368966 210280 374342
rect 210344 369102 210372 460566
rect 210332 369096 210384 369102
rect 210332 369038 210384 369044
rect 210240 368960 210292 368966
rect 210240 368902 210292 368908
rect 210436 162178 210464 468794
rect 210514 458960 210570 458969
rect 210514 458895 210570 458904
rect 210528 162450 210556 458895
rect 210620 266966 210648 474030
rect 210700 463480 210752 463486
rect 210700 463422 210752 463428
rect 210712 269278 210740 463422
rect 210804 374406 210832 477498
rect 211264 475402 211292 480023
rect 211344 478712 211396 478718
rect 211342 478680 211344 478689
rect 211396 478680 211398 478689
rect 211342 478615 211398 478624
rect 211172 475374 211292 475402
rect 211066 374640 211122 374649
rect 211066 374575 211122 374584
rect 210792 374400 210844 374406
rect 210792 374342 210844 374348
rect 210976 372564 211028 372570
rect 210976 372506 211028 372512
rect 210988 372230 211016 372506
rect 210976 372224 211028 372230
rect 210976 372166 211028 372172
rect 210976 371612 211028 371618
rect 210976 371554 211028 371560
rect 210988 370870 211016 371554
rect 210976 370864 211028 370870
rect 210976 370806 211028 370812
rect 210884 369028 210936 369034
rect 210884 368970 210936 368976
rect 210792 368960 210844 368966
rect 210792 368902 210844 368908
rect 210700 269272 210752 269278
rect 210700 269214 210752 269220
rect 210608 266960 210660 266966
rect 210608 266902 210660 266908
rect 210698 265160 210754 265169
rect 210698 265095 210754 265104
rect 210516 162444 210568 162450
rect 210516 162386 210568 162392
rect 210424 162172 210476 162178
rect 210424 162114 210476 162120
rect 210712 144702 210740 265095
rect 210804 264382 210832 368902
rect 210896 264994 210924 368970
rect 210988 265033 211016 370806
rect 210974 265024 211030 265033
rect 210884 264988 210936 264994
rect 210974 264959 211030 264968
rect 210884 264930 210936 264936
rect 210792 264376 210844 264382
rect 210792 264318 210844 264324
rect 210700 144696 210752 144702
rect 210700 144638 210752 144644
rect 211080 57866 211108 374575
rect 211172 374490 211200 475374
rect 211816 470594 211844 480023
rect 212264 478236 212316 478242
rect 212264 478178 212316 478184
rect 211988 476944 212040 476950
rect 211988 476886 212040 476892
rect 211264 470566 211844 470594
rect 211264 379514 211292 470566
rect 211804 469872 211856 469878
rect 211804 469814 211856 469820
rect 211620 459468 211672 459474
rect 211620 459410 211672 459416
rect 211264 379486 211476 379514
rect 211172 374462 211292 374490
rect 211158 373688 211214 373697
rect 211158 373623 211214 373632
rect 211172 372638 211200 373623
rect 211160 372632 211212 372638
rect 211160 372574 211212 372580
rect 211264 372366 211292 374462
rect 211448 373697 211476 379486
rect 211434 373688 211490 373697
rect 211434 373623 211490 373632
rect 211252 372360 211304 372366
rect 211252 372302 211304 372308
rect 211264 372162 211292 372302
rect 211252 372156 211304 372162
rect 211252 372098 211304 372104
rect 211632 369646 211660 459410
rect 211710 371784 211766 371793
rect 211710 371719 211766 371728
rect 211620 369640 211672 369646
rect 211620 369582 211672 369588
rect 211526 270600 211582 270609
rect 211526 270535 211582 270544
rect 211540 160886 211568 270535
rect 211724 270502 211752 371719
rect 211712 270496 211764 270502
rect 211618 270464 211674 270473
rect 211712 270438 211764 270444
rect 211618 270399 211674 270408
rect 211528 160880 211580 160886
rect 211528 160822 211580 160828
rect 211632 58954 211660 270399
rect 211816 162586 211844 469814
rect 211894 463312 211950 463321
rect 211894 463247 211950 463256
rect 211908 163606 211936 463247
rect 212000 267170 212028 476886
rect 212080 463684 212132 463690
rect 212080 463626 212132 463632
rect 212092 267345 212120 463626
rect 212172 463412 212224 463418
rect 212172 463354 212224 463360
rect 212184 269210 212212 463354
rect 212276 370870 212304 478178
rect 212552 475522 212580 480037
rect 212644 480023 213026 480051
rect 213104 480023 213394 480051
rect 213472 480023 213854 480051
rect 214024 480023 214314 480051
rect 214392 480023 214774 480051
rect 214944 480023 215234 480051
rect 215404 480023 215602 480051
rect 215680 480023 216062 480051
rect 216232 480023 216522 480051
rect 212540 475516 212592 475522
rect 212540 475458 212592 475464
rect 212540 475380 212592 475386
rect 212540 475322 212592 475328
rect 212552 373454 212580 475322
rect 212540 373448 212592 373454
rect 212540 373390 212592 373396
rect 212644 373046 212672 480023
rect 213104 475386 213132 480023
rect 213092 475380 213144 475386
rect 213092 475322 213144 475328
rect 212724 475312 212776 475318
rect 213472 475266 213500 480023
rect 213920 475380 213972 475386
rect 213920 475322 213972 475328
rect 212724 475254 212776 475260
rect 212736 373153 212764 475254
rect 212828 475238 213500 475266
rect 212722 373144 212778 373153
rect 212722 373079 212778 373088
rect 212632 373040 212684 373046
rect 212632 372982 212684 372988
rect 212356 372564 212408 372570
rect 212356 372506 212408 372512
rect 212368 371958 212396 372506
rect 212356 371952 212408 371958
rect 212356 371894 212408 371900
rect 212264 370864 212316 370870
rect 212264 370806 212316 370812
rect 212264 369164 212316 369170
rect 212264 369106 212316 369112
rect 212172 269204 212224 269210
rect 212172 269146 212224 269152
rect 212078 267336 212134 267345
rect 212078 267271 212134 267280
rect 211988 267164 212040 267170
rect 211988 267106 212040 267112
rect 212078 265840 212134 265849
rect 212078 265775 212134 265784
rect 212092 265033 212120 265775
rect 212170 265568 212226 265577
rect 212170 265503 212226 265512
rect 212078 265024 212134 265033
rect 212078 264959 212134 264968
rect 211896 163600 211948 163606
rect 211896 163542 211948 163548
rect 211804 162580 211856 162586
rect 211804 162522 211856 162528
rect 212092 147626 212120 264959
rect 212184 148918 212212 265503
rect 212276 265062 212304 369106
rect 212264 265056 212316 265062
rect 212264 264998 212316 265004
rect 212368 264926 212396 371894
rect 212448 371476 212500 371482
rect 212448 371418 212500 371424
rect 212460 265713 212488 371418
rect 212644 369753 212672 372982
rect 212828 372910 212856 475238
rect 213184 472660 213236 472666
rect 213184 472602 213236 472608
rect 213092 373380 213144 373386
rect 213092 373322 213144 373328
rect 212816 372904 212868 372910
rect 212816 372846 212868 372852
rect 212828 369854 212856 372846
rect 212736 369826 212856 369854
rect 212630 369744 212686 369753
rect 212630 369679 212686 369688
rect 212736 369306 212764 369826
rect 212724 369300 212776 369306
rect 212724 369242 212776 369248
rect 213104 368898 213132 373322
rect 213092 368892 213144 368898
rect 213092 368834 213144 368840
rect 213104 354674 213132 368834
rect 213012 354646 213132 354674
rect 212908 270496 212960 270502
rect 212908 270438 212960 270444
rect 212920 269414 212948 270438
rect 212908 269408 212960 269414
rect 212908 269350 212960 269356
rect 212446 265704 212502 265713
rect 212446 265639 212502 265648
rect 212460 265033 212488 265639
rect 212446 265024 212502 265033
rect 212446 264959 212502 264968
rect 212356 264920 212408 264926
rect 212356 264862 212408 264868
rect 212172 148912 212224 148918
rect 212172 148854 212224 148860
rect 212080 147620 212132 147626
rect 212080 147562 212132 147568
rect 211620 58948 211672 58954
rect 211620 58890 211672 58896
rect 211068 57860 211120 57866
rect 211068 57802 211120 57808
rect 165618 57559 165674 57568
rect 209688 57588 209740 57594
rect 153290 56264 153346 56273
rect 153290 56199 153346 56208
rect 155972 54913 156000 57559
rect 160112 55049 160140 57559
rect 165632 55185 165660 57559
rect 209688 57530 209740 57536
rect 165618 55176 165674 55185
rect 165618 55111 165674 55120
rect 160098 55040 160154 55049
rect 160098 54975 160154 54984
rect 155958 54904 156014 54913
rect 155958 54839 156014 54848
rect 89720 54742 89772 54748
rect 118698 54768 118754 54777
rect 80060 54732 80112 54738
rect 212184 54738 212212 148854
rect 212368 144770 212396 264862
rect 212920 148510 212948 269350
rect 213012 265130 213040 354646
rect 213092 272604 213144 272610
rect 213092 272546 213144 272552
rect 213104 265946 213132 272546
rect 213196 266898 213224 472602
rect 213460 463548 213512 463554
rect 213460 463490 213512 463496
rect 213276 461644 213328 461650
rect 213276 461586 213328 461592
rect 213184 266892 213236 266898
rect 213184 266834 213236 266840
rect 213092 265940 213144 265946
rect 213092 265882 213144 265888
rect 213000 265124 213052 265130
rect 213000 265066 213052 265072
rect 213090 265024 213146 265033
rect 213090 264959 213146 264968
rect 213104 151814 213132 264959
rect 213184 251184 213236 251190
rect 213184 251126 213236 251132
rect 213196 249830 213224 251126
rect 213184 249824 213236 249830
rect 213184 249766 213236 249772
rect 213196 173194 213224 249766
rect 213184 173188 213236 173194
rect 213184 173130 213236 173136
rect 213288 162042 213316 461586
rect 213366 458824 213422 458833
rect 213366 458759 213422 458768
rect 213380 163742 213408 458759
rect 213472 268462 213500 463490
rect 213552 460352 213604 460358
rect 213552 460294 213604 460300
rect 213460 268456 213512 268462
rect 213460 268398 213512 268404
rect 213564 267374 213592 460294
rect 213932 374626 213960 475322
rect 213840 374598 213960 374626
rect 213840 373946 213868 374598
rect 213920 374536 213972 374542
rect 213920 374478 213972 374484
rect 213932 374066 213960 374478
rect 213920 374060 213972 374066
rect 213920 374002 213972 374008
rect 213840 373918 213960 373946
rect 213736 373176 213788 373182
rect 213736 373118 213788 373124
rect 213644 372020 213696 372026
rect 213644 371962 213696 371968
rect 213656 371346 213684 371962
rect 213644 371340 213696 371346
rect 213644 371282 213696 371288
rect 213656 272610 213684 371282
rect 213644 272604 213696 272610
rect 213644 272546 213696 272552
rect 213748 269226 213776 373118
rect 213932 372978 213960 373918
rect 213920 372972 213972 372978
rect 213920 372914 213972 372920
rect 213932 371074 213960 372914
rect 214024 372842 214052 480023
rect 214392 470594 214420 480023
rect 214564 477556 214616 477562
rect 214564 477498 214616 477504
rect 214116 470566 214420 470594
rect 214116 373386 214144 470566
rect 214380 373516 214432 373522
rect 214380 373458 214432 373464
rect 214104 373380 214156 373386
rect 214104 373322 214156 373328
rect 214012 372836 214064 372842
rect 214012 372778 214064 372784
rect 213920 371068 213972 371074
rect 213920 371010 213972 371016
rect 213826 369200 213882 369209
rect 214024 369170 214052 372778
rect 214392 371754 214420 373458
rect 214576 372230 214604 477498
rect 214944 475386 214972 480023
rect 214932 475380 214984 475386
rect 214932 475322 214984 475328
rect 215300 475380 215352 475386
rect 215300 475322 215352 475328
rect 214656 467288 214708 467294
rect 214656 467230 214708 467236
rect 214564 372224 214616 372230
rect 214564 372166 214616 372172
rect 214380 371748 214432 371754
rect 214380 371690 214432 371696
rect 213826 369135 213882 369144
rect 214012 369164 214064 369170
rect 213656 269198 213776 269226
rect 213656 269074 213684 269198
rect 213734 269104 213790 269113
rect 213644 269068 213696 269074
rect 213734 269039 213790 269048
rect 213644 269010 213696 269016
rect 213552 267368 213604 267374
rect 213552 267310 213604 267316
rect 213644 266144 213696 266150
rect 213644 266086 213696 266092
rect 213656 265946 213684 266086
rect 213644 265940 213696 265946
rect 213644 265882 213696 265888
rect 213460 264240 213512 264246
rect 213460 264182 213512 264188
rect 213368 163736 213420 163742
rect 213368 163678 213420 163684
rect 213276 162036 213328 162042
rect 213276 161978 213328 161984
rect 213368 160880 213420 160886
rect 213368 160822 213420 160828
rect 213380 160682 213408 160822
rect 213368 160676 213420 160682
rect 213368 160618 213420 160624
rect 213104 151786 213316 151814
rect 213288 148850 213316 151786
rect 213276 148844 213328 148850
rect 213276 148786 213328 148792
rect 212908 148504 212960 148510
rect 212908 148446 212960 148452
rect 212356 144764 212408 144770
rect 212356 144706 212408 144712
rect 118698 54703 118754 54712
rect 212172 54732 212224 54738
rect 80060 54674 80112 54680
rect 212172 54674 212224 54680
rect 213288 54534 213316 148786
rect 213380 55894 213408 160618
rect 213472 144838 213500 264182
rect 213552 149048 213604 149054
rect 213552 148990 213604 148996
rect 213564 148510 213592 148990
rect 213552 148504 213604 148510
rect 213552 148446 213604 148452
rect 213460 144832 213512 144838
rect 213460 144774 213512 144780
rect 213368 55888 213420 55894
rect 213368 55830 213420 55836
rect 213564 55214 213592 148446
rect 213656 144906 213684 265882
rect 213644 144900 213696 144906
rect 213644 144842 213696 144848
rect 213748 57662 213776 269039
rect 213736 57656 213788 57662
rect 213736 57598 213788 57604
rect 213840 57186 213868 369135
rect 214012 369106 214064 369112
rect 214288 269068 214340 269074
rect 214288 269010 214340 269016
rect 214300 267918 214328 269010
rect 214288 267912 214340 267918
rect 214288 267854 214340 267860
rect 214300 258074 214328 267854
rect 214392 265674 214420 371690
rect 214564 355360 214616 355366
rect 214564 355302 214616 355308
rect 214576 278322 214604 355302
rect 214564 278316 214616 278322
rect 214564 278258 214616 278264
rect 214576 276622 214604 278258
rect 214564 276616 214616 276622
rect 214564 276558 214616 276564
rect 214668 266762 214696 467230
rect 214840 466336 214892 466342
rect 214840 466278 214892 466284
rect 214748 460420 214800 460426
rect 214748 460362 214800 460368
rect 214760 269346 214788 460362
rect 214852 369170 214880 466278
rect 215208 459672 215260 459678
rect 215208 459614 215260 459620
rect 215116 374060 215168 374066
rect 215116 374002 215168 374008
rect 215024 372496 215076 372502
rect 215024 372438 215076 372444
rect 214930 372056 214986 372065
rect 214930 371991 214986 372000
rect 214840 369164 214892 369170
rect 214840 369106 214892 369112
rect 214838 368384 214894 368393
rect 214838 368319 214894 368328
rect 214852 367810 214880 368319
rect 214840 367804 214892 367810
rect 214840 367746 214892 367752
rect 214748 269340 214800 269346
rect 214748 269282 214800 269288
rect 214656 266756 214708 266762
rect 214656 266698 214708 266704
rect 214564 266484 214616 266490
rect 214564 266426 214616 266432
rect 214380 265668 214432 265674
rect 214380 265610 214432 265616
rect 214300 258046 214512 258074
rect 214484 145518 214512 258046
rect 214576 151814 214604 266426
rect 214656 266416 214708 266422
rect 214656 266358 214708 266364
rect 214668 160750 214696 266358
rect 214852 265606 214880 367746
rect 214944 267034 214972 371991
rect 214932 267028 214984 267034
rect 214932 266970 214984 266976
rect 214944 266490 214972 266970
rect 214932 266484 214984 266490
rect 214932 266426 214984 266432
rect 215036 265742 215064 372438
rect 215128 267073 215156 374002
rect 215220 372473 215248 459614
rect 215312 373794 215340 475322
rect 215300 373788 215352 373794
rect 215300 373730 215352 373736
rect 215300 373652 215352 373658
rect 215300 373594 215352 373600
rect 215312 373250 215340 373594
rect 215300 373244 215352 373250
rect 215300 373186 215352 373192
rect 215404 372774 215432 480023
rect 215680 470594 215708 480023
rect 216128 475720 216180 475726
rect 216128 475662 216180 475668
rect 215944 474020 215996 474026
rect 215944 473962 215996 473968
rect 215496 470566 215708 470594
rect 215496 373994 215524 470566
rect 215850 374368 215906 374377
rect 215850 374303 215906 374312
rect 215864 373994 215892 374303
rect 215496 373966 215892 373994
rect 215392 372768 215444 372774
rect 215392 372710 215444 372716
rect 215206 372464 215262 372473
rect 215206 372399 215262 372408
rect 215404 371249 215432 372710
rect 215390 371240 215446 371249
rect 215390 371175 215446 371184
rect 215300 276616 215352 276622
rect 215300 276558 215352 276564
rect 215114 267064 215170 267073
rect 215114 266999 215170 267008
rect 215024 265736 215076 265742
rect 215024 265678 215076 265684
rect 214840 265600 214892 265606
rect 214840 265542 214892 265548
rect 214748 264988 214800 264994
rect 214748 264930 214800 264936
rect 214656 160744 214708 160750
rect 214656 160686 214708 160692
rect 214760 159390 214788 264930
rect 215024 264376 215076 264382
rect 215024 264318 215076 264324
rect 214932 264308 214984 264314
rect 214932 264250 214984 264256
rect 214748 159384 214800 159390
rect 214748 159326 214800 159332
rect 214576 151786 214880 151814
rect 214852 148986 214880 151786
rect 214840 148980 214892 148986
rect 214840 148922 214892 148928
rect 214562 145888 214618 145897
rect 214562 145823 214618 145832
rect 214472 145512 214524 145518
rect 214472 145454 214524 145460
rect 213828 57180 213880 57186
rect 213828 57122 213880 57128
rect 214484 56574 214512 145454
rect 214576 144702 214604 145823
rect 214654 145752 214710 145761
rect 214654 145687 214710 145696
rect 214668 144838 214696 145687
rect 214748 145580 214800 145586
rect 214748 145522 214800 145528
rect 214760 144906 214788 145522
rect 214748 144900 214800 144906
rect 214748 144842 214800 144848
rect 214656 144832 214708 144838
rect 214656 144774 214708 144780
rect 214564 144696 214616 144702
rect 214564 144638 214616 144644
rect 214472 56568 214524 56574
rect 214472 56510 214524 56516
rect 213552 55208 213604 55214
rect 213552 55150 213604 55156
rect 213276 54528 213328 54534
rect 213276 54470 213328 54476
rect 214576 54466 214604 144638
rect 214668 55078 214696 144774
rect 214760 56030 214788 144842
rect 214748 56024 214800 56030
rect 214748 55966 214800 55972
rect 214852 55146 214880 148922
rect 214944 146305 214972 264250
rect 214930 146296 214986 146305
rect 214930 146231 214986 146240
rect 214944 56370 214972 146231
rect 215036 145246 215064 264318
rect 215128 145382 215156 266999
rect 215312 251190 215340 276558
rect 215404 266422 215432 371175
rect 215864 369617 215892 373966
rect 215850 369608 215906 369617
rect 215850 369543 215906 369552
rect 215392 266416 215444 266422
rect 215392 266358 215444 266364
rect 215574 266384 215630 266393
rect 215574 266319 215630 266328
rect 215300 251184 215352 251190
rect 215300 251126 215352 251132
rect 215208 158772 215260 158778
rect 215208 158714 215260 158720
rect 215116 145376 215168 145382
rect 215116 145318 215168 145324
rect 215024 145240 215076 145246
rect 215024 145182 215076 145188
rect 214932 56364 214984 56370
rect 214932 56306 214984 56312
rect 214840 55140 214892 55146
rect 214840 55082 214892 55088
rect 214656 55072 214708 55078
rect 214656 55014 214708 55020
rect 215036 54670 215064 145182
rect 215220 59498 215248 158714
rect 215588 145450 215616 266319
rect 215760 265124 215812 265130
rect 215760 265066 215812 265072
rect 215668 265056 215720 265062
rect 215668 264998 215720 265004
rect 215680 160002 215708 264998
rect 215772 160070 215800 265066
rect 215864 251190 215892 369543
rect 215852 251184 215904 251190
rect 215852 251126 215904 251132
rect 215864 161474 215892 251126
rect 215956 162518 215984 473962
rect 216036 468784 216088 468790
rect 216036 468726 216088 468732
rect 215944 162512 215996 162518
rect 215944 162454 215996 162460
rect 216048 162246 216076 468726
rect 216140 267646 216168 475662
rect 216232 475386 216260 480023
rect 216680 478372 216732 478378
rect 216680 478314 216732 478320
rect 216220 475380 216272 475386
rect 216220 475322 216272 475328
rect 216312 466268 216364 466274
rect 216312 466210 216364 466216
rect 216220 460488 216272 460494
rect 216220 460430 216272 460436
rect 216232 268666 216260 460430
rect 216324 369306 216352 466210
rect 216588 459604 216640 459610
rect 216588 459546 216640 459552
rect 216496 373244 216548 373250
rect 216496 373186 216548 373192
rect 216404 371408 216456 371414
rect 216404 371350 216456 371356
rect 216312 369300 216364 369306
rect 216312 369242 216364 369248
rect 216220 268660 216272 268666
rect 216220 268602 216272 268608
rect 216128 267640 216180 267646
rect 216128 267582 216180 267588
rect 216416 267209 216444 371350
rect 216402 267200 216458 267209
rect 216402 267135 216458 267144
rect 216312 265736 216364 265742
rect 216312 265678 216364 265684
rect 216220 265668 216272 265674
rect 216220 265610 216272 265616
rect 216036 162240 216088 162246
rect 216036 162182 216088 162188
rect 215864 161446 216076 161474
rect 216048 161362 216076 161446
rect 216036 161356 216088 161362
rect 216036 161298 216088 161304
rect 215760 160064 215812 160070
rect 215760 160006 215812 160012
rect 215668 159996 215720 160002
rect 215668 159938 215720 159944
rect 215680 158778 215708 159938
rect 215772 159254 215800 160006
rect 215760 159248 215812 159254
rect 215760 159190 215812 159196
rect 215668 158772 215720 158778
rect 215668 158714 215720 158720
rect 215852 148368 215904 148374
rect 215852 148310 215904 148316
rect 215864 147626 215892 148310
rect 215852 147620 215904 147626
rect 215852 147562 215904 147568
rect 215864 147506 215892 147562
rect 215864 147478 215984 147506
rect 215850 145616 215906 145625
rect 215850 145551 215906 145560
rect 215576 145444 215628 145450
rect 215576 145386 215628 145392
rect 215864 144770 215892 145551
rect 215852 144764 215904 144770
rect 215852 144706 215904 144712
rect 215208 59492 215260 59498
rect 215208 59434 215260 59440
rect 215864 55758 215892 144706
rect 215956 56506 215984 147478
rect 216048 59430 216076 161298
rect 216128 160744 216180 160750
rect 216128 160686 216180 160692
rect 216036 59424 216088 59430
rect 216036 59366 216088 59372
rect 216140 59090 216168 160686
rect 216232 145722 216260 265610
rect 216220 145716 216272 145722
rect 216220 145658 216272 145664
rect 216128 59084 216180 59090
rect 216128 59026 216180 59032
rect 215944 56500 215996 56506
rect 215944 56442 215996 56448
rect 215852 55752 215904 55758
rect 215852 55694 215904 55700
rect 216232 54806 216260 145658
rect 216324 145654 216352 265678
rect 216416 265169 216444 267135
rect 216508 266937 216536 373186
rect 216600 371385 216628 459546
rect 216692 384334 216720 478314
rect 216968 477601 216996 480037
rect 217324 478168 217376 478174
rect 217324 478110 217376 478116
rect 216954 477592 217010 477601
rect 216954 477527 217010 477536
rect 217336 477442 217364 478110
rect 217428 477601 217456 480037
rect 217796 477601 217824 480037
rect 218164 480023 218270 480051
rect 218440 480023 218730 480051
rect 218808 480023 219190 480051
rect 217414 477592 217470 477601
rect 217414 477527 217470 477536
rect 217782 477592 217838 477601
rect 217782 477527 217838 477536
rect 217336 477414 217456 477442
rect 217324 474156 217376 474162
rect 217324 474098 217376 474104
rect 216772 409148 216824 409154
rect 216772 409090 216824 409096
rect 216784 408785 216812 409090
rect 216770 408776 216826 408785
rect 216770 408711 216826 408720
rect 216680 384328 216732 384334
rect 216680 384270 216732 384276
rect 216680 383648 216732 383654
rect 216680 383590 216732 383596
rect 216692 383353 216720 383590
rect 216678 383344 216734 383353
rect 216678 383279 216734 383288
rect 216784 375057 216812 408711
rect 216864 405000 216916 405006
rect 216862 404968 216864 404977
rect 216916 404968 216918 404977
rect 216862 404903 216918 404912
rect 216876 383602 216904 404903
rect 217336 403209 217364 474098
rect 217322 403200 217378 403209
rect 217322 403135 217378 403144
rect 217336 393314 217364 403135
rect 217152 393286 217364 393314
rect 216956 385008 217008 385014
rect 216954 384976 216956 384985
rect 217008 384976 217010 384985
rect 216954 384911 217010 384920
rect 216876 383574 216996 383602
rect 216862 375320 216918 375329
rect 216862 375255 216918 375264
rect 216770 375048 216826 375057
rect 216770 374983 216826 374992
rect 216586 371376 216642 371385
rect 216586 371311 216642 371320
rect 216586 369200 216642 369209
rect 216586 369135 216642 369144
rect 216494 266928 216550 266937
rect 216494 266863 216550 266872
rect 216508 266393 216536 266863
rect 216494 266384 216550 266393
rect 216494 266319 216550 266328
rect 216402 265160 216458 265169
rect 216402 265095 216458 265104
rect 216494 251152 216550 251161
rect 216494 251087 216550 251096
rect 216404 159248 216456 159254
rect 216404 159190 216456 159196
rect 216312 145648 216364 145654
rect 216312 145590 216364 145596
rect 216220 54800 216272 54806
rect 216220 54742 216272 54748
rect 215024 54664 215076 54670
rect 215024 54606 215076 54612
rect 216324 54602 216352 145590
rect 216416 59566 216444 159190
rect 216404 59560 216456 59566
rect 216404 59502 216456 59508
rect 216508 57390 216536 251087
rect 216496 57384 216548 57390
rect 216496 57326 216548 57332
rect 216600 57322 216628 369135
rect 216678 307728 216734 307737
rect 216678 307663 216734 307672
rect 216692 287054 216720 307663
rect 216784 303793 216812 374983
rect 216876 374921 216904 375255
rect 216968 375018 216996 383574
rect 217048 383580 217100 383586
rect 217048 383522 217100 383528
rect 217060 383081 217088 383522
rect 217046 383072 217102 383081
rect 217046 383007 217102 383016
rect 217152 375329 217180 393286
rect 217232 375352 217284 375358
rect 217138 375320 217194 375329
rect 217232 375294 217284 375300
rect 217138 375255 217194 375264
rect 217244 375086 217272 375294
rect 217232 375080 217284 375086
rect 217232 375022 217284 375028
rect 216956 375012 217008 375018
rect 216956 374954 217008 374960
rect 216862 374912 216918 374921
rect 216862 374847 216918 374856
rect 216770 303784 216826 303793
rect 216770 303719 216826 303728
rect 216876 299441 216904 374847
rect 216968 299985 216996 374954
rect 217140 372904 217192 372910
rect 217140 372846 217192 372852
rect 217048 372632 217100 372638
rect 217048 372574 217100 372580
rect 217060 305969 217088 372574
rect 217046 305960 217102 305969
rect 217046 305895 217102 305904
rect 216954 299976 217010 299985
rect 216954 299911 217010 299920
rect 216862 299432 216918 299441
rect 216862 299367 216918 299376
rect 216692 287026 216812 287054
rect 216680 280152 216732 280158
rect 216680 280094 216732 280100
rect 216692 279993 216720 280094
rect 216678 279984 216734 279993
rect 216678 279919 216734 279928
rect 216678 278352 216734 278361
rect 216678 278287 216680 278296
rect 216732 278287 216734 278296
rect 216680 278258 216732 278264
rect 216784 267734 216812 287026
rect 216864 278724 216916 278730
rect 216864 278666 216916 278672
rect 216876 278089 216904 278666
rect 216862 278080 216918 278089
rect 216862 278015 216918 278024
rect 216692 267706 216812 267734
rect 216692 202881 216720 267706
rect 216772 266212 216824 266218
rect 216772 266154 216824 266160
rect 216678 202872 216734 202881
rect 216678 202807 216734 202816
rect 216680 175228 216732 175234
rect 216680 175170 216732 175176
rect 216692 175001 216720 175170
rect 216678 174992 216734 175001
rect 216678 174927 216734 174936
rect 216678 173360 216734 173369
rect 216678 173295 216734 173304
rect 216692 173194 216720 173295
rect 216680 173188 216732 173194
rect 216680 173130 216732 173136
rect 216784 146062 216812 266154
rect 216862 202872 216918 202881
rect 216862 202807 216918 202816
rect 216876 201929 216904 202807
rect 216862 201920 216918 201929
rect 216862 201855 216918 201864
rect 216772 146056 216824 146062
rect 216772 145998 216824 146004
rect 216876 96937 216904 201855
rect 217060 200977 217088 305895
rect 217152 269074 217180 372846
rect 217244 302841 217272 375022
rect 217428 371074 217456 477414
rect 218060 475380 218112 475386
rect 218060 475322 218112 475328
rect 217600 469940 217652 469946
rect 217600 469882 217652 469888
rect 217508 463616 217560 463622
rect 217508 463558 217560 463564
rect 217520 374270 217548 463558
rect 217612 406065 217640 469882
rect 217692 467356 217744 467362
rect 217692 467298 217744 467304
rect 217704 410961 217732 467298
rect 217876 457496 217928 457502
rect 217876 457438 217928 457444
rect 217784 417444 217836 417450
rect 217784 417386 217836 417392
rect 217796 411913 217824 417386
rect 217782 411904 217838 411913
rect 217782 411839 217838 411848
rect 217690 410952 217746 410961
rect 217690 410887 217746 410896
rect 217598 406056 217654 406065
rect 217598 405991 217654 406000
rect 217508 374264 217560 374270
rect 217508 374206 217560 374212
rect 217612 373994 217640 405991
rect 217704 373998 217732 410887
rect 217520 373966 217640 373994
rect 217692 373992 217744 373998
rect 217520 373930 217548 373966
rect 217692 373934 217744 373940
rect 217508 373924 217560 373930
rect 217508 373866 217560 373872
rect 217416 371068 217468 371074
rect 217416 371010 217468 371016
rect 217230 302832 217286 302841
rect 217230 302767 217286 302776
rect 217140 269068 217192 269074
rect 217140 269010 217192 269016
rect 217140 251116 217192 251122
rect 217140 251058 217192 251064
rect 217046 200968 217102 200977
rect 217046 200903 217102 200912
rect 217060 200114 217088 200903
rect 216968 200086 217088 200114
rect 216862 96928 216918 96937
rect 216862 96863 216918 96872
rect 216968 95985 216996 200086
rect 217048 173800 217100 173806
rect 217048 173742 217100 173748
rect 217060 173097 217088 173742
rect 217046 173088 217102 173097
rect 217046 173023 217102 173032
rect 217152 146266 217180 251058
rect 217244 197849 217272 302767
rect 217520 301073 217548 373866
rect 217704 372638 217732 373934
rect 217692 372632 217744 372638
rect 217692 372574 217744 372580
rect 217796 307737 217824 411839
rect 217888 407833 217916 457438
rect 217874 407824 217930 407833
rect 217874 407759 217930 407768
rect 217888 375358 217916 407759
rect 217876 375352 217928 375358
rect 217876 375294 217928 375300
rect 217876 373788 217928 373794
rect 217876 373730 217928 373736
rect 217888 372706 217916 373730
rect 217968 373040 218020 373046
rect 217968 372982 218020 372988
rect 217876 372700 217928 372706
rect 217876 372642 217928 372648
rect 217888 369238 217916 372642
rect 217876 369232 217928 369238
rect 217876 369174 217928 369180
rect 217782 307728 217838 307737
rect 217782 307663 217838 307672
rect 217796 306921 217824 307663
rect 217782 306912 217838 306921
rect 217782 306847 217838 306856
rect 217690 303784 217746 303793
rect 217690 303719 217746 303728
rect 217506 301064 217562 301073
rect 217506 300999 217562 301008
rect 217414 299976 217470 299985
rect 217414 299911 217470 299920
rect 217230 197840 217286 197849
rect 217230 197775 217286 197784
rect 217140 146260 217192 146266
rect 217140 146202 217192 146208
rect 216954 95976 217010 95985
rect 216954 95911 217010 95920
rect 216678 68368 216734 68377
rect 216678 68303 216734 68312
rect 216692 67658 216720 68303
rect 216680 67652 216732 67658
rect 216680 67594 216732 67600
rect 217152 59702 217180 146202
rect 217244 92857 217272 197775
rect 217428 194993 217456 299911
rect 217520 196081 217548 300999
rect 217598 299432 217654 299441
rect 217598 299367 217654 299376
rect 217612 298217 217640 299367
rect 217598 298208 217654 298217
rect 217598 298143 217654 298152
rect 217506 196072 217562 196081
rect 217506 196007 217562 196016
rect 217414 194984 217470 194993
rect 217414 194919 217470 194928
rect 217230 92848 217286 92857
rect 217230 92783 217286 92792
rect 217428 90001 217456 194919
rect 217612 193225 217640 298143
rect 217704 198801 217732 303719
rect 217784 269068 217836 269074
rect 217784 269010 217836 269016
rect 217796 267850 217824 269010
rect 217784 267844 217836 267850
rect 217784 267786 217836 267792
rect 217690 198792 217746 198801
rect 217690 198727 217746 198736
rect 217690 196072 217746 196081
rect 217690 196007 217746 196016
rect 217598 193216 217654 193225
rect 217598 193151 217654 193160
rect 217612 180794 217640 193151
rect 217520 180766 217640 180794
rect 217414 89992 217470 90001
rect 217414 89927 217470 89936
rect 217520 88233 217548 180766
rect 217704 91089 217732 196007
rect 217796 161090 217824 267786
rect 217888 265742 217916 369174
rect 217876 265736 217928 265742
rect 217876 265678 217928 265684
rect 217980 251122 218008 372982
rect 218072 372570 218100 475322
rect 218060 372564 218112 372570
rect 218060 372506 218112 372512
rect 218164 372337 218192 480023
rect 218440 470594 218468 480023
rect 218704 476876 218756 476882
rect 218704 476818 218756 476824
rect 218256 470566 218468 470594
rect 218716 470594 218744 476818
rect 218808 475386 218836 480023
rect 219544 475658 219572 480037
rect 219636 480023 220018 480051
rect 220096 480023 220478 480051
rect 219532 475652 219584 475658
rect 219532 475594 219584 475600
rect 219636 475538 219664 480023
rect 219452 475510 219664 475538
rect 218796 475380 218848 475386
rect 218796 475322 218848 475328
rect 218716 470566 218836 470594
rect 218256 374241 218284 470566
rect 218702 463040 218758 463049
rect 218702 462975 218758 462984
rect 218336 460896 218388 460902
rect 218336 460838 218388 460844
rect 218348 459785 218376 460838
rect 218334 459776 218390 459785
rect 218334 459711 218390 459720
rect 218242 374232 218298 374241
rect 218242 374167 218298 374176
rect 218150 372328 218206 372337
rect 218150 372263 218206 372272
rect 218428 353456 218480 353462
rect 218428 353398 218480 353404
rect 218334 270464 218390 270473
rect 218334 270399 218390 270408
rect 217968 251116 218020 251122
rect 217968 251058 218020 251064
rect 217966 198792 218022 198801
rect 217966 198727 218022 198736
rect 217784 161084 217836 161090
rect 217784 161026 217836 161032
rect 217690 91080 217746 91089
rect 217690 91015 217746 91024
rect 217506 88224 217562 88233
rect 217506 88159 217562 88168
rect 217140 59696 217192 59702
rect 217140 59638 217192 59644
rect 217796 59226 217824 161026
rect 217874 146024 217930 146033
rect 217874 145959 217930 145968
rect 217888 145926 217916 145959
rect 217876 145920 217928 145926
rect 217876 145862 217928 145868
rect 217876 145784 217928 145790
rect 217876 145726 217928 145732
rect 217784 59220 217836 59226
rect 217784 59162 217836 59168
rect 216588 57316 216640 57322
rect 216588 57258 216640 57264
rect 217888 54874 217916 145726
rect 217980 93809 218008 198727
rect 218244 162920 218296 162926
rect 218244 162862 218296 162868
rect 217966 93800 218022 93809
rect 217966 93735 218022 93744
rect 217966 68368 218022 68377
rect 217966 68303 218022 68312
rect 217980 59362 218008 68303
rect 217968 59356 218020 59362
rect 217968 59298 218020 59304
rect 218256 56302 218284 162862
rect 218348 57526 218376 270399
rect 218440 266218 218468 353398
rect 218612 353388 218664 353394
rect 218612 353330 218664 353336
rect 218520 353320 218572 353326
rect 218520 353262 218572 353268
rect 218532 269482 218560 353262
rect 218520 269476 218572 269482
rect 218520 269418 218572 269424
rect 218624 266286 218652 353330
rect 218612 266280 218664 266286
rect 218612 266222 218664 266228
rect 218428 266212 218480 266218
rect 218428 266154 218480 266160
rect 218520 265600 218572 265606
rect 218520 265542 218572 265548
rect 218532 162926 218560 265542
rect 218520 162920 218572 162926
rect 218520 162862 218572 162868
rect 218428 160132 218480 160138
rect 218428 160074 218480 160080
rect 218440 59634 218468 160074
rect 218612 145784 218664 145790
rect 218612 145726 218664 145732
rect 218520 145444 218572 145450
rect 218520 145386 218572 145392
rect 218532 59770 218560 145386
rect 218520 59764 218572 59770
rect 218520 59706 218572 59712
rect 218428 59628 218480 59634
rect 218428 59570 218480 59576
rect 218336 57520 218388 57526
rect 218336 57462 218388 57468
rect 218244 56296 218296 56302
rect 218244 56238 218296 56244
rect 218624 55962 218652 145726
rect 218716 57254 218744 462975
rect 218808 161974 218836 470566
rect 219164 466064 219216 466070
rect 219164 466006 219216 466012
rect 218886 465760 218942 465769
rect 218886 465695 218942 465704
rect 218900 162654 218928 465695
rect 218980 460284 219032 460290
rect 218980 460226 219032 460232
rect 218888 162648 218940 162654
rect 218888 162590 218940 162596
rect 218992 162314 219020 460226
rect 219072 459196 219124 459202
rect 219072 459138 219124 459144
rect 219084 266830 219112 459138
rect 219176 369238 219204 466006
rect 219348 372972 219400 372978
rect 219348 372914 219400 372920
rect 219254 372736 219310 372745
rect 219254 372671 219310 372680
rect 219268 372638 219296 372671
rect 219256 372632 219308 372638
rect 219256 372574 219308 372580
rect 219164 369232 219216 369238
rect 219164 369174 219216 369180
rect 219268 270094 219296 372574
rect 219256 270088 219308 270094
rect 219256 270030 219308 270036
rect 219360 267782 219388 372914
rect 219452 372298 219480 475510
rect 219532 475448 219584 475454
rect 220096 475402 220124 480023
rect 220176 477556 220228 477562
rect 220176 477498 220228 477504
rect 219532 475390 219584 475396
rect 219440 372292 219492 372298
rect 219440 372234 219492 372240
rect 219544 372065 219572 475390
rect 219636 475374 220124 475402
rect 219636 374105 219664 475374
rect 220188 470594 220216 477498
rect 220004 470566 220216 470594
rect 219622 374096 219678 374105
rect 219622 374031 219678 374040
rect 219898 373144 219954 373153
rect 219898 373079 219954 373088
rect 219716 372224 219768 372230
rect 219716 372166 219768 372172
rect 219624 372088 219676 372094
rect 219530 372056 219586 372065
rect 219624 372030 219676 372036
rect 219530 371991 219586 372000
rect 219532 371816 219584 371822
rect 219532 371758 219584 371764
rect 219348 267776 219400 267782
rect 219348 267718 219400 267724
rect 219072 266824 219124 266830
rect 219072 266766 219124 266772
rect 219164 266280 219216 266286
rect 219164 266222 219216 266228
rect 219072 266076 219124 266082
rect 219072 266018 219124 266024
rect 218980 162308 219032 162314
rect 218980 162250 219032 162256
rect 218796 161968 218848 161974
rect 218796 161910 218848 161916
rect 218888 159384 218940 159390
rect 218888 159326 218940 159332
rect 218796 146124 218848 146130
rect 218796 146066 218848 146072
rect 218704 57248 218756 57254
rect 218704 57190 218756 57196
rect 218808 56166 218836 146066
rect 218900 59294 218928 159326
rect 219084 145994 219112 266018
rect 219176 146130 219204 266222
rect 219256 265940 219308 265946
rect 219256 265882 219308 265888
rect 219164 146124 219216 146130
rect 219164 146066 219216 146072
rect 219072 145988 219124 145994
rect 219072 145930 219124 145936
rect 218978 60616 219034 60625
rect 218978 60551 219034 60560
rect 218888 59288 218940 59294
rect 218888 59230 218940 59236
rect 218992 57730 219020 60551
rect 218980 57724 219032 57730
rect 218980 57666 219032 57672
rect 218796 56160 218848 56166
rect 218796 56102 218848 56108
rect 219084 56098 219112 145930
rect 219268 145790 219296 265882
rect 219360 161158 219388 267718
rect 219544 265946 219572 371758
rect 219636 265985 219664 372030
rect 219728 266082 219756 372166
rect 219808 270088 219860 270094
rect 219808 270030 219860 270036
rect 219820 269618 219848 270030
rect 219808 269612 219860 269618
rect 219808 269554 219860 269560
rect 219716 266076 219768 266082
rect 219716 266018 219768 266024
rect 219622 265976 219678 265985
rect 219532 265940 219584 265946
rect 219622 265911 219678 265920
rect 219532 265882 219584 265888
rect 219716 265736 219768 265742
rect 219716 265678 219768 265684
rect 219624 250504 219676 250510
rect 219624 250446 219676 250452
rect 219636 171134 219664 250446
rect 219544 171106 219664 171134
rect 219544 161430 219572 171106
rect 219728 161474 219756 265678
rect 219636 161446 219756 161474
rect 219532 161424 219584 161430
rect 219532 161366 219584 161372
rect 219348 161152 219400 161158
rect 219348 161094 219400 161100
rect 219360 160138 219388 161094
rect 219348 160132 219400 160138
rect 219348 160074 219400 160080
rect 219256 145784 219308 145790
rect 219256 145726 219308 145732
rect 219164 145376 219216 145382
rect 219164 145318 219216 145324
rect 219176 56438 219204 145318
rect 219254 60616 219310 60625
rect 219254 60551 219310 60560
rect 219268 58682 219296 60551
rect 219256 58676 219308 58682
rect 219256 58618 219308 58624
rect 219164 56432 219216 56438
rect 219164 56374 219216 56380
rect 219072 56092 219124 56098
rect 219072 56034 219124 56040
rect 218612 55956 218664 55962
rect 218612 55898 218664 55904
rect 219544 55010 219572 161366
rect 219636 161226 219664 161446
rect 219820 161294 219848 269554
rect 219912 264858 219940 373079
rect 219900 264852 219952 264858
rect 219900 264794 219952 264800
rect 219808 161288 219860 161294
rect 219808 161230 219860 161236
rect 219624 161220 219676 161226
rect 219624 161162 219676 161168
rect 219636 59158 219664 161162
rect 219624 59152 219676 59158
rect 219624 59094 219676 59100
rect 219820 56234 219848 161230
rect 219912 146198 219940 264794
rect 219900 146192 219952 146198
rect 219900 146134 219952 146140
rect 219808 56228 219860 56234
rect 219808 56170 219860 56176
rect 219532 55004 219584 55010
rect 219532 54946 219584 54952
rect 219912 54942 219940 146134
rect 220004 55826 220032 470566
rect 220924 459610 220952 480037
rect 221016 480023 221398 480051
rect 221016 459678 221044 480023
rect 221752 478310 221780 480037
rect 221740 478304 221792 478310
rect 221740 478246 221792 478252
rect 222212 475386 222240 480037
rect 222672 477562 222700 480037
rect 223132 477601 223160 480037
rect 223118 477592 223174 477601
rect 222660 477556 222712 477562
rect 223118 477527 223174 477536
rect 222660 477498 222712 477504
rect 223592 475561 223620 480037
rect 223684 480023 223974 480051
rect 223578 475552 223634 475561
rect 223578 475487 223634 475496
rect 223684 475402 223712 480023
rect 224420 478378 224448 480037
rect 224512 480023 224894 480051
rect 224408 478372 224460 478378
rect 224408 478314 224460 478320
rect 222200 475380 222252 475386
rect 222200 475322 222252 475328
rect 223592 475374 223712 475402
rect 221004 459672 221056 459678
rect 221004 459614 221056 459620
rect 220912 459604 220964 459610
rect 220912 459546 220964 459552
rect 223592 458862 223620 475374
rect 224512 470594 224540 480023
rect 225340 478242 225368 480037
rect 225328 478236 225380 478242
rect 225328 478178 225380 478184
rect 225708 478174 225736 480037
rect 226168 478281 226196 480037
rect 226642 480023 226672 480051
rect 226644 479890 226672 480023
rect 226904 480023 227102 480051
rect 227180 480023 227562 480051
rect 227732 480023 227930 480051
rect 226644 479862 226840 479890
rect 226154 478272 226210 478281
rect 226154 478207 226210 478216
rect 225696 478168 225748 478174
rect 225696 478110 225748 478116
rect 226812 471306 226840 479862
rect 226800 471300 226852 471306
rect 226800 471242 226852 471248
rect 226904 471186 226932 480023
rect 223684 470566 224540 470594
rect 226352 471158 226932 471186
rect 223684 469849 223712 470566
rect 223670 469840 223726 469849
rect 223670 469775 223726 469784
rect 226352 465798 226380 471158
rect 227180 470594 227208 480023
rect 226444 470566 227208 470594
rect 226340 465792 226392 465798
rect 226340 465734 226392 465740
rect 226444 465730 226472 470566
rect 227732 467158 227760 480023
rect 228376 474026 228404 480037
rect 228836 474162 228864 480037
rect 229112 480023 229310 480051
rect 229480 480023 229770 480051
rect 228824 474156 228876 474162
rect 228824 474098 228876 474104
rect 228364 474020 228416 474026
rect 228364 473962 228416 473968
rect 227720 467152 227772 467158
rect 227720 467094 227772 467100
rect 229112 465769 229140 480023
rect 229480 470594 229508 480023
rect 230124 472841 230152 480037
rect 230584 478310 230612 480037
rect 230572 478304 230624 478310
rect 230572 478246 230624 478252
rect 230110 472832 230166 472841
rect 230110 472767 230166 472776
rect 231044 471209 231072 480037
rect 231504 478417 231532 480037
rect 231490 478408 231546 478417
rect 231490 478343 231546 478352
rect 231872 472569 231900 480037
rect 232332 478514 232360 480037
rect 232320 478508 232372 478514
rect 232320 478450 232372 478456
rect 232792 472705 232820 480037
rect 233252 478553 233280 480037
rect 233238 478544 233294 478553
rect 233238 478479 233294 478488
rect 233712 474065 233740 480037
rect 234080 478281 234108 480037
rect 234066 478272 234122 478281
rect 234066 478207 234122 478216
rect 234540 478145 234568 480037
rect 234632 480023 235014 480051
rect 234526 478136 234582 478145
rect 234526 478071 234582 478080
rect 233698 474056 233754 474065
rect 233698 473991 233754 474000
rect 232778 472696 232834 472705
rect 232778 472631 232834 472640
rect 231858 472560 231914 472569
rect 231858 472495 231914 472504
rect 231030 471200 231086 471209
rect 231030 471135 231086 471144
rect 229204 470566 229508 470594
rect 229204 469878 229232 470566
rect 229192 469872 229244 469878
rect 229192 469814 229244 469820
rect 234632 468489 234660 480023
rect 235460 478446 235488 480037
rect 235920 478825 235948 480037
rect 235906 478816 235962 478825
rect 235906 478751 235962 478760
rect 236288 478689 236316 480037
rect 236274 478680 236330 478689
rect 236274 478615 236330 478624
rect 235448 478440 235500 478446
rect 235448 478382 235500 478388
rect 236748 476882 236776 480037
rect 236840 480023 237222 480051
rect 237392 480023 237682 480051
rect 236736 476876 236788 476882
rect 236736 476818 236788 476824
rect 236840 470594 236868 480023
rect 236012 470566 236868 470594
rect 234618 468480 234674 468489
rect 234618 468415 234674 468424
rect 229098 465760 229154 465769
rect 226432 465724 226484 465730
rect 229098 465695 229154 465704
rect 226432 465666 226484 465672
rect 236012 458930 236040 470566
rect 237392 467226 237420 480023
rect 238128 474094 238156 480037
rect 238116 474088 238168 474094
rect 238116 474030 238168 474036
rect 238496 472734 238524 480037
rect 238956 478718 238984 480037
rect 238944 478712 238996 478718
rect 238944 478654 238996 478660
rect 238484 472728 238536 472734
rect 238484 472670 238536 472676
rect 239416 472666 239444 480037
rect 239876 478650 239904 480037
rect 239864 478644 239916 478650
rect 239864 478586 239916 478592
rect 240244 478582 240272 480037
rect 240336 480023 240718 480051
rect 240796 480023 241178 480051
rect 241532 480023 241638 480051
rect 241808 480023 242098 480051
rect 240232 478576 240284 478582
rect 240232 478518 240284 478524
rect 240336 475300 240364 480023
rect 240152 475272 240364 475300
rect 239404 472660 239456 472666
rect 239404 472602 239456 472608
rect 237380 467220 237432 467226
rect 237380 467162 237432 467168
rect 240152 463010 240180 475272
rect 240796 470594 240824 480023
rect 240244 470566 240824 470594
rect 240244 465934 240272 470566
rect 240232 465928 240284 465934
rect 240232 465870 240284 465876
rect 241532 465866 241560 480023
rect 241808 470594 241836 480023
rect 242452 474230 242480 480037
rect 242912 477018 242940 480037
rect 242900 477012 242952 477018
rect 242900 476954 242952 476960
rect 243372 475522 243400 480037
rect 243464 480023 243846 480051
rect 244306 480023 244336 480051
rect 243360 475516 243412 475522
rect 243360 475458 243412 475464
rect 242440 474224 242492 474230
rect 242440 474166 242492 474172
rect 243464 470594 243492 480023
rect 244308 479890 244336 480023
rect 244568 480023 244674 480051
rect 244752 480023 245134 480051
rect 245304 480023 245594 480051
rect 245764 480023 246054 480051
rect 246132 480023 246422 480051
rect 246592 480023 246882 480051
rect 244308 479862 244504 479890
rect 244280 475312 244332 475318
rect 244280 475254 244332 475260
rect 241624 470566 241836 470594
rect 242912 470566 243492 470594
rect 241624 468586 241652 470566
rect 242912 469946 242940 470566
rect 242900 469940 242952 469946
rect 242900 469882 242952 469888
rect 241612 468580 241664 468586
rect 241612 468522 241664 468528
rect 241520 465860 241572 465866
rect 241520 465802 241572 465808
rect 240140 463004 240192 463010
rect 240140 462946 240192 462952
rect 244292 459066 244320 475254
rect 244476 471374 244504 479862
rect 244568 475318 244596 480023
rect 244556 475312 244608 475318
rect 244556 475254 244608 475260
rect 244464 471368 244516 471374
rect 244464 471310 244516 471316
rect 244752 471186 244780 480023
rect 244384 471158 244780 471186
rect 244384 460358 244412 471158
rect 245304 470594 245332 480023
rect 245660 475312 245712 475318
rect 245660 475254 245712 475260
rect 244476 470566 245332 470594
rect 244476 467294 244504 470566
rect 244464 467288 244516 467294
rect 244464 467230 244516 467236
rect 244372 460352 244424 460358
rect 244372 460294 244424 460300
rect 244280 459060 244332 459066
rect 244280 459002 244332 459008
rect 245672 458998 245700 475254
rect 245764 468654 245792 480023
rect 246132 470594 246160 480023
rect 246592 475318 246620 480023
rect 247328 476950 247356 480037
rect 247316 476944 247368 476950
rect 247316 476886 247368 476892
rect 247788 475454 247816 480037
rect 247880 480023 248262 480051
rect 248432 480023 248630 480051
rect 248800 480023 249090 480051
rect 249168 480023 249550 480051
rect 249812 480023 250010 480051
rect 250088 480023 250470 480051
rect 250548 480023 250838 480051
rect 247776 475448 247828 475454
rect 247776 475390 247828 475396
rect 246580 475312 246632 475318
rect 246580 475254 246632 475260
rect 247880 470594 247908 480023
rect 245856 470566 246160 470594
rect 247052 470566 247908 470594
rect 245856 470014 245884 470566
rect 245844 470008 245896 470014
rect 245844 469950 245896 469956
rect 245752 468648 245804 468654
rect 245752 468590 245804 468596
rect 247052 460222 247080 470566
rect 248432 460426 248460 480023
rect 248512 475312 248564 475318
rect 248512 475254 248564 475260
rect 248420 460420 248472 460426
rect 248420 460362 248472 460368
rect 248524 460290 248552 475254
rect 248800 470594 248828 480023
rect 249168 475318 249196 480023
rect 249156 475312 249208 475318
rect 249156 475254 249208 475260
rect 248616 470566 248828 470594
rect 248616 463078 248644 470566
rect 248604 463072 248656 463078
rect 248604 463014 248656 463020
rect 249812 460494 249840 480023
rect 250088 475402 250116 480023
rect 249904 475374 250116 475402
rect 249904 460630 249932 475374
rect 250548 470594 250576 480023
rect 251180 475312 251232 475318
rect 251180 475254 251232 475260
rect 249996 470566 250576 470594
rect 249996 463146 250024 470566
rect 249984 463140 250036 463146
rect 249984 463082 250036 463088
rect 249892 460624 249944 460630
rect 249892 460566 249944 460572
rect 251192 460562 251220 475254
rect 251284 461718 251312 480037
rect 251376 480023 251758 480051
rect 251376 475318 251404 480023
rect 251364 475312 251416 475318
rect 251364 475254 251416 475260
rect 252204 474298 252232 480037
rect 252586 480023 252692 480051
rect 252560 475312 252612 475318
rect 252560 475254 252612 475260
rect 252192 474292 252244 474298
rect 252192 474234 252244 474240
rect 251272 461712 251324 461718
rect 251272 461654 251324 461660
rect 252572 461650 252600 475254
rect 252664 470082 252692 480023
rect 253032 475590 253060 480037
rect 253216 480023 253506 480051
rect 253020 475584 253072 475590
rect 253020 475526 253072 475532
rect 253216 475318 253244 480023
rect 253204 475312 253256 475318
rect 253204 475254 253256 475260
rect 253952 471442 253980 480037
rect 254136 480023 254426 480051
rect 253940 471436 253992 471442
rect 253940 471378 253992 471384
rect 254136 470594 254164 480023
rect 254780 474434 254808 480037
rect 254768 474428 254820 474434
rect 254768 474370 254820 474376
rect 255240 474366 255268 480037
rect 255700 476785 255728 480037
rect 255792 480023 256174 480051
rect 255686 476776 255742 476785
rect 255686 476711 255742 476720
rect 255228 474360 255280 474366
rect 255228 474302 255280 474308
rect 255792 470594 255820 480023
rect 256620 477086 256648 480037
rect 256712 480023 257002 480051
rect 256608 477080 256660 477086
rect 256608 477022 256660 477028
rect 253952 470566 254164 470594
rect 255332 470566 255820 470594
rect 252652 470076 252704 470082
rect 252652 470018 252704 470024
rect 253952 467430 253980 470566
rect 255332 468625 255360 470566
rect 255318 468616 255374 468625
rect 255318 468551 255374 468560
rect 253940 467424 253992 467430
rect 253940 467366 253992 467372
rect 252560 461644 252612 461650
rect 252560 461586 252612 461592
rect 251180 460556 251232 460562
rect 251180 460498 251232 460504
rect 249800 460488 249852 460494
rect 249800 460430 249852 460436
rect 248512 460284 248564 460290
rect 248512 460226 248564 460232
rect 247040 460216 247092 460222
rect 247040 460158 247092 460164
rect 256712 459134 256740 480023
rect 257448 471578 257476 480037
rect 257540 480023 257922 480051
rect 258092 480023 258382 480051
rect 257436 471572 257488 471578
rect 257436 471514 257488 471520
rect 257540 470594 257568 480023
rect 256804 470566 257568 470594
rect 256804 459270 256832 470566
rect 258092 467362 258120 480023
rect 258828 472802 258856 480037
rect 258920 480023 259210 480051
rect 258816 472796 258868 472802
rect 258816 472738 258868 472744
rect 258920 470594 258948 480023
rect 259460 475312 259512 475318
rect 259460 475254 259512 475260
rect 258184 470566 258948 470594
rect 258184 470150 258212 470566
rect 258172 470144 258224 470150
rect 258172 470086 258224 470092
rect 258080 467356 258132 467362
rect 258080 467298 258132 467304
rect 259472 460698 259500 475254
rect 259656 471510 259684 480037
rect 259840 480023 260130 480051
rect 260208 480023 260590 480051
rect 259644 471504 259696 471510
rect 259644 471446 259696 471452
rect 259840 470594 259868 480023
rect 260208 475318 260236 480023
rect 260196 475312 260248 475318
rect 260196 475254 260248 475260
rect 260944 474502 260972 480037
rect 261128 480023 261418 480051
rect 260932 474496 260984 474502
rect 260932 474438 260984 474444
rect 261128 470594 261156 480023
rect 261864 477154 261892 480037
rect 261852 477148 261904 477154
rect 261852 477090 261904 477096
rect 262220 475312 262272 475318
rect 262220 475254 262272 475260
rect 259564 470566 259868 470594
rect 260852 470566 261156 470594
rect 259564 468722 259592 470566
rect 259552 468716 259604 468722
rect 259552 468658 259604 468664
rect 260852 462058 260880 470566
rect 260840 462052 260892 462058
rect 260840 461994 260892 462000
rect 259460 460692 259512 460698
rect 259460 460634 259512 460640
rect 256792 459264 256844 459270
rect 256792 459206 256844 459212
rect 262232 459202 262260 475254
rect 262324 461786 262352 480037
rect 262416 480023 262798 480051
rect 262876 480023 263166 480051
rect 263626 480023 263732 480051
rect 262416 475318 262444 480023
rect 262404 475312 262456 475318
rect 262404 475254 262456 475260
rect 262876 470594 262904 480023
rect 262416 470566 262904 470594
rect 262416 468790 262444 470566
rect 262404 468784 262456 468790
rect 263704 468761 263732 480023
rect 263796 480023 264086 480051
rect 264256 480023 264546 480051
rect 263796 468858 263824 480023
rect 263784 468852 263836 468858
rect 263784 468794 263836 468800
rect 262404 468726 262456 468732
rect 263690 468752 263746 468761
rect 263690 468687 263746 468696
rect 264256 466454 264284 480023
rect 263612 466426 264284 466454
rect 263612 461922 263640 466426
rect 263600 461916 263652 461922
rect 263600 461858 263652 461864
rect 264992 461854 265020 480037
rect 265084 480023 265374 480051
rect 265084 467634 265112 480023
rect 265820 471646 265848 480037
rect 266280 471714 266308 480037
rect 266372 480023 266754 480051
rect 266268 471708 266320 471714
rect 266268 471650 266320 471656
rect 265808 471640 265860 471646
rect 265808 471582 265860 471588
rect 265072 467628 265124 467634
rect 265072 467570 265124 467576
rect 264980 461848 265032 461854
rect 264980 461790 265032 461796
rect 262312 461780 262364 461786
rect 262312 461722 262364 461728
rect 266372 460766 266400 480023
rect 267108 475794 267136 480037
rect 267568 475862 267596 480037
rect 267844 480023 268042 480051
rect 268120 480023 268502 480051
rect 268672 480023 268962 480051
rect 269224 480023 269330 480051
rect 269408 480023 269790 480051
rect 269960 480023 270250 480051
rect 267556 475856 267608 475862
rect 267556 475798 267608 475804
rect 267096 475788 267148 475794
rect 267096 475730 267148 475736
rect 267740 471232 267792 471238
rect 267740 471174 267792 471180
rect 267752 463214 267780 471174
rect 267844 463350 267872 480023
rect 268120 471238 268148 480023
rect 268108 471232 268160 471238
rect 268108 471174 268160 471180
rect 268672 467498 268700 480023
rect 269224 467566 269252 480023
rect 269212 467560 269264 467566
rect 269212 467502 269264 467508
rect 268660 467492 268712 467498
rect 268660 467434 268712 467440
rect 269408 466454 269436 480023
rect 269960 470218 269988 480023
rect 270696 471850 270724 480037
rect 270684 471844 270736 471850
rect 270684 471786 270736 471792
rect 271156 471345 271184 480037
rect 271248 480023 271538 480051
rect 271892 480023 271998 480051
rect 271142 471336 271198 471345
rect 271142 471271 271198 471280
rect 269948 470212 270000 470218
rect 269948 470154 270000 470160
rect 271248 468994 271276 480023
rect 271236 468988 271288 468994
rect 271236 468930 271288 468936
rect 269132 466426 269436 466454
rect 267832 463344 267884 463350
rect 267832 463286 267884 463292
rect 267740 463208 267792 463214
rect 267740 463150 267792 463156
rect 269132 461990 269160 466426
rect 269120 461984 269172 461990
rect 269120 461926 269172 461932
rect 266360 460760 266412 460766
rect 266360 460702 266412 460708
rect 271892 459338 271920 480023
rect 272444 471782 272472 480037
rect 272904 475658 272932 480037
rect 273272 475726 273300 480037
rect 273364 480023 273746 480051
rect 273824 480023 274206 480051
rect 274666 480023 274772 480051
rect 273260 475720 273312 475726
rect 273260 475662 273312 475668
rect 272892 475652 272944 475658
rect 272892 475594 272944 475600
rect 273364 475402 273392 480023
rect 273272 475374 273392 475402
rect 272432 471776 272484 471782
rect 272432 471718 272484 471724
rect 273272 463418 273300 475374
rect 273824 470594 273852 480023
rect 274744 475930 274772 480023
rect 274836 480023 275126 480051
rect 274732 475924 274784 475930
rect 274732 475866 274784 475872
rect 274836 475538 274864 480023
rect 274916 475924 274968 475930
rect 274916 475866 274968 475872
rect 273364 470566 273852 470594
rect 274652 475510 274864 475538
rect 273364 468926 273392 470566
rect 273352 468920 273404 468926
rect 273352 468862 273404 468868
rect 273260 463412 273312 463418
rect 273260 463354 273312 463360
rect 274652 463282 274680 475510
rect 274928 475266 274956 475866
rect 274744 475238 274956 475266
rect 274744 469062 274772 475238
rect 275480 473074 275508 480037
rect 275940 474570 275968 480037
rect 276216 480023 276414 480051
rect 276584 480023 276874 480051
rect 276952 480023 277334 480051
rect 277596 480023 277702 480051
rect 277872 480023 278162 480051
rect 278240 480023 278622 480051
rect 279082 480023 279112 480051
rect 276112 475312 276164 475318
rect 276112 475254 276164 475260
rect 276020 475244 276072 475250
rect 276020 475186 276072 475192
rect 275928 474564 275980 474570
rect 275928 474506 275980 474512
rect 275468 473068 275520 473074
rect 275468 473010 275520 473016
rect 274732 469056 274784 469062
rect 274732 468998 274784 469004
rect 274640 463276 274692 463282
rect 274640 463218 274692 463224
rect 276032 459406 276060 475186
rect 276124 462913 276152 475254
rect 276216 463554 276244 480023
rect 276584 475318 276612 480023
rect 276572 475312 276624 475318
rect 276572 475254 276624 475260
rect 276952 475250 276980 480023
rect 277492 475312 277544 475318
rect 277492 475254 277544 475260
rect 276940 475244 276992 475250
rect 276940 475186 276992 475192
rect 277400 475244 277452 475250
rect 277400 475186 277452 475192
rect 276204 463548 276256 463554
rect 276204 463490 276256 463496
rect 277412 463486 277440 475186
rect 277400 463480 277452 463486
rect 277400 463422 277452 463428
rect 277504 463049 277532 475254
rect 277596 463622 277624 480023
rect 277872 475318 277900 480023
rect 277860 475312 277912 475318
rect 277860 475254 277912 475260
rect 278240 475250 278268 480023
rect 279084 479890 279112 480023
rect 279344 480023 279542 480051
rect 279620 480023 279910 480051
rect 280172 480023 280370 480051
rect 279084 479862 279280 479890
rect 278228 475244 278280 475250
rect 278228 475186 278280 475192
rect 279252 472938 279280 479862
rect 279240 472932 279292 472938
rect 279240 472874 279292 472880
rect 279344 472818 279372 480023
rect 278792 472790 279372 472818
rect 277584 463616 277636 463622
rect 277584 463558 277636 463564
rect 277490 463040 277546 463049
rect 277490 462975 277546 462984
rect 276110 462904 276166 462913
rect 276110 462839 276166 462848
rect 278792 460154 278820 472790
rect 279620 470594 279648 480023
rect 278884 470566 279648 470594
rect 278884 470354 278912 470566
rect 278872 470348 278924 470354
rect 278872 470290 278924 470296
rect 280172 462126 280200 480023
rect 280816 472870 280844 480037
rect 281000 480023 281290 480051
rect 281552 480023 281658 480051
rect 280804 472864 280856 472870
rect 280804 472806 280856 472812
rect 281000 470594 281028 480023
rect 280264 470566 281028 470594
rect 280264 469985 280292 470566
rect 280250 469976 280306 469985
rect 280250 469911 280306 469920
rect 280160 462120 280212 462126
rect 280160 462062 280212 462068
rect 278780 460148 278832 460154
rect 278780 460090 278832 460096
rect 281552 459474 281580 480023
rect 282104 474638 282132 480037
rect 282564 477222 282592 480037
rect 283024 477290 283052 480037
rect 283116 480023 283498 480051
rect 283576 480023 283866 480051
rect 284326 480023 284432 480051
rect 283012 477284 283064 477290
rect 283012 477226 283064 477232
rect 282552 477216 282604 477222
rect 282552 477158 282604 477164
rect 283116 475402 283144 480023
rect 282932 475374 283144 475402
rect 282092 474632 282144 474638
rect 282092 474574 282144 474580
rect 282932 463690 282960 475374
rect 283576 470594 283604 480023
rect 284300 475312 284352 475318
rect 284300 475254 284352 475260
rect 283024 470566 283604 470594
rect 283024 464778 283052 470566
rect 283012 464772 283064 464778
rect 283012 464714 283064 464720
rect 284312 464370 284340 475254
rect 284404 464710 284432 480023
rect 284496 480023 284786 480051
rect 284864 480023 285246 480051
rect 285706 480023 285812 480051
rect 284392 464704 284444 464710
rect 284392 464646 284444 464652
rect 284496 464642 284524 480023
rect 284864 475318 284892 480023
rect 284852 475312 284904 475318
rect 284852 475254 284904 475260
rect 285680 475312 285732 475318
rect 285680 475254 285732 475260
rect 284484 464636 284536 464642
rect 284484 464578 284536 464584
rect 284300 464364 284352 464370
rect 284300 464306 284352 464312
rect 282920 463684 282972 463690
rect 282920 463626 282972 463632
rect 285692 460902 285720 475254
rect 285784 464438 285812 480023
rect 285876 480023 286074 480051
rect 286152 480023 286534 480051
rect 286704 480023 286994 480051
rect 287072 480023 287454 480051
rect 287532 480023 287822 480051
rect 287900 480023 288282 480051
rect 285876 467770 285904 480023
rect 286152 470594 286180 480023
rect 286704 475318 286732 480023
rect 286692 475312 286744 475318
rect 286692 475254 286744 475260
rect 285968 470566 286180 470594
rect 285968 470286 285996 470566
rect 285956 470280 286008 470286
rect 285956 470222 286008 470228
rect 285864 467764 285916 467770
rect 285864 467706 285916 467712
rect 285772 464432 285824 464438
rect 285772 464374 285824 464380
rect 285680 460896 285732 460902
rect 285680 460838 285732 460844
rect 287072 460834 287100 480023
rect 287532 475402 287560 480023
rect 287164 475374 287560 475402
rect 287164 462262 287192 475374
rect 287900 470594 287928 480023
rect 288728 471918 288756 480037
rect 288820 480023 289202 480051
rect 289280 480023 289662 480051
rect 289832 480023 290030 480051
rect 290200 480023 290490 480051
rect 288716 471912 288768 471918
rect 288716 471854 288768 471860
rect 288820 471730 288848 480023
rect 287256 470566 287928 470594
rect 288452 471702 288848 471730
rect 287256 465905 287284 470566
rect 287242 465896 287298 465905
rect 287242 465831 287298 465840
rect 287152 462256 287204 462262
rect 287152 462198 287204 462204
rect 287060 460828 287112 460834
rect 287060 460770 287112 460776
rect 288452 460018 288480 471702
rect 289280 470594 289308 480023
rect 288544 470566 289308 470594
rect 288544 466002 288572 470566
rect 289832 466274 289860 480023
rect 290200 470594 290228 480023
rect 290936 477358 290964 480037
rect 291304 480023 291410 480051
rect 290924 477352 290976 477358
rect 290924 477294 290976 477300
rect 291200 475312 291252 475318
rect 291200 475254 291252 475260
rect 289924 470566 290228 470594
rect 289924 469130 289952 470566
rect 289912 469124 289964 469130
rect 289912 469066 289964 469072
rect 289820 466268 289872 466274
rect 289820 466210 289872 466216
rect 288532 465996 288584 466002
rect 288532 465938 288584 465944
rect 291212 460086 291240 475254
rect 291304 464506 291332 480023
rect 291856 475930 291884 480037
rect 291948 480023 292238 480051
rect 292592 480023 292698 480051
rect 292776 480023 293158 480051
rect 291844 475924 291896 475930
rect 291844 475866 291896 475872
rect 291948 475318 291976 480023
rect 291936 475312 291988 475318
rect 291936 475254 291988 475260
rect 291292 464500 291344 464506
rect 291292 464442 291344 464448
rect 291200 460080 291252 460086
rect 291200 460022 291252 460028
rect 288440 460012 288492 460018
rect 288440 459954 288492 459960
rect 281540 459468 281592 459474
rect 281540 459410 281592 459416
rect 276020 459400 276072 459406
rect 276020 459342 276072 459348
rect 271880 459332 271932 459338
rect 271880 459274 271932 459280
rect 262220 459196 262272 459202
rect 262220 459138 262272 459144
rect 256700 459128 256752 459134
rect 256700 459070 256752 459076
rect 245660 458992 245712 458998
rect 245660 458934 245712 458940
rect 236000 458924 236052 458930
rect 236000 458866 236052 458872
rect 223580 458856 223632 458862
rect 223580 458798 223632 458804
rect 292592 458794 292620 480023
rect 292776 470594 292804 480023
rect 293604 474706 293632 480037
rect 293986 480023 294092 480051
rect 294064 475998 294092 480023
rect 294156 480023 294446 480051
rect 294524 480023 294906 480051
rect 294052 475992 294104 475998
rect 294052 475934 294104 475940
rect 294156 475538 294184 480023
rect 294236 475992 294288 475998
rect 294236 475934 294288 475940
rect 293972 475510 294184 475538
rect 293592 474700 293644 474706
rect 293592 474642 293644 474648
rect 292684 470566 292804 470594
rect 292684 464846 292712 470566
rect 292672 464840 292724 464846
rect 292672 464782 292724 464788
rect 293972 464574 294000 475510
rect 294248 475130 294276 475934
rect 294064 475102 294276 475130
rect 294064 464914 294092 475102
rect 294524 470594 294552 480023
rect 295352 473958 295380 480037
rect 295340 473952 295392 473958
rect 295340 473894 295392 473900
rect 295812 473006 295840 480037
rect 295800 473000 295852 473006
rect 295800 472942 295852 472948
rect 296180 471986 296208 480037
rect 296272 480023 296654 480051
rect 296168 471980 296220 471986
rect 296168 471922 296220 471928
rect 296272 470594 296300 480023
rect 297100 477426 297128 480037
rect 297192 480023 297574 480051
rect 297744 480023 298034 480051
rect 298402 480023 298432 480051
rect 297088 477420 297140 477426
rect 297088 477362 297140 477368
rect 296720 475312 296772 475318
rect 296720 475254 296772 475260
rect 294156 470566 294552 470594
rect 295352 470566 296300 470594
rect 294156 467702 294184 470566
rect 294144 467696 294196 467702
rect 294144 467638 294196 467644
rect 294052 464908 294104 464914
rect 294052 464850 294104 464856
rect 293960 464568 294012 464574
rect 293960 464510 294012 464516
rect 295352 459542 295380 470566
rect 296732 464409 296760 475254
rect 297192 470594 297220 480023
rect 297744 475318 297772 480023
rect 298404 479890 298432 480023
rect 298664 480023 298862 480051
rect 298940 480023 299322 480051
rect 298404 479862 298600 479890
rect 297732 475312 297784 475318
rect 297732 475254 297784 475260
rect 298572 473142 298600 479862
rect 298560 473136 298612 473142
rect 298560 473078 298612 473084
rect 298664 472954 298692 480023
rect 296824 470566 297220 470594
rect 298112 472926 298692 472954
rect 296824 466138 296852 470566
rect 296812 466132 296864 466138
rect 296812 466074 296864 466080
rect 296718 464400 296774 464409
rect 296718 464335 296774 464344
rect 298112 462194 298140 472926
rect 298940 470594 298968 480023
rect 299860 470594 299888 480134
rect 356704 478712 356756 478718
rect 356704 478654 356756 478660
rect 298204 470566 298968 470594
rect 299492 470566 299888 470594
rect 298204 466070 298232 470566
rect 299492 466206 299520 470566
rect 299480 466200 299532 466206
rect 299480 466142 299532 466148
rect 298192 466064 298244 466070
rect 298192 466006 298244 466012
rect 298100 462188 298152 462194
rect 298100 462130 298152 462136
rect 338304 461100 338356 461106
rect 338304 461042 338356 461048
rect 338316 461009 338344 461042
rect 339776 461032 339828 461038
rect 338302 461000 338358 461009
rect 338302 460935 338304 460944
rect 338356 460935 338358 460944
rect 339774 461000 339776 461009
rect 339828 461000 339830 461009
rect 339774 460935 339830 460944
rect 350998 461000 351054 461009
rect 350998 460935 351000 460944
rect 338304 460906 338356 460912
rect 351052 460935 351054 460944
rect 351000 460906 351052 460912
rect 295340 459536 295392 459542
rect 295340 459478 295392 459484
rect 292580 458788 292632 458794
rect 292580 458730 292632 458736
rect 275284 374876 275336 374882
rect 275284 374818 275336 374824
rect 235998 374504 236054 374513
rect 235998 374439 236054 374448
rect 244278 374504 244334 374513
rect 244278 374439 244334 374448
rect 250074 374504 250130 374513
rect 250074 374439 250130 374448
rect 250718 374504 250774 374513
rect 250718 374439 250774 374448
rect 251270 374504 251326 374513
rect 251270 374439 251326 374448
rect 256054 374504 256110 374513
rect 256054 374439 256110 374448
rect 270498 374504 270554 374513
rect 270498 374439 270554 374448
rect 222014 374232 222070 374241
rect 222014 374167 222070 374176
rect 221922 374096 221978 374105
rect 221922 374031 221978 374040
rect 221830 373688 221886 373697
rect 221830 373623 221886 373632
rect 220818 373280 220874 373289
rect 220818 373215 220874 373224
rect 220726 373144 220782 373153
rect 220726 373079 220728 373088
rect 220780 373079 220782 373088
rect 220728 373050 220780 373056
rect 220728 372292 220780 372298
rect 220728 372234 220780 372240
rect 220544 372224 220596 372230
rect 220544 372166 220596 372172
rect 220556 372026 220584 372166
rect 220544 372020 220596 372026
rect 220544 371962 220596 371968
rect 220740 371278 220768 372234
rect 220728 371272 220780 371278
rect 220728 371214 220780 371220
rect 220832 353326 220860 373215
rect 221096 372156 221148 372162
rect 221096 372098 221148 372104
rect 220912 371952 220964 371958
rect 220912 371894 220964 371900
rect 220924 353394 220952 371894
rect 221004 371272 221056 371278
rect 221004 371214 221056 371220
rect 221016 353433 221044 371214
rect 221108 353462 221136 372098
rect 221844 371958 221872 373623
rect 221832 371952 221884 371958
rect 221936 371929 221964 374031
rect 222028 372201 222056 374167
rect 236012 374066 236040 374439
rect 244292 374406 244320 374439
rect 244280 374400 244332 374406
rect 244280 374342 244332 374348
rect 250088 374134 250116 374439
rect 250732 374202 250760 374439
rect 250720 374196 250772 374202
rect 250720 374138 250772 374144
rect 241060 374128 241112 374134
rect 241060 374070 241112 374076
rect 250076 374128 250128 374134
rect 250076 374070 250128 374076
rect 236000 374060 236052 374066
rect 236000 374002 236052 374008
rect 224224 373516 224276 373522
rect 224224 373458 224276 373464
rect 222014 372192 222070 372201
rect 222014 372127 222070 372136
rect 222108 372156 222160 372162
rect 222108 372098 222160 372104
rect 221832 371894 221884 371900
rect 221922 371920 221978 371929
rect 221922 371855 221978 371864
rect 222120 371686 222148 372098
rect 224236 371890 224264 373458
rect 236458 373416 236514 373425
rect 236458 373351 236514 373360
rect 236472 373250 236500 373351
rect 236460 373244 236512 373250
rect 236460 373186 236512 373192
rect 238114 372600 238170 372609
rect 238114 372535 238170 372544
rect 239310 372600 239366 372609
rect 239310 372535 239366 372544
rect 240414 372600 240470 372609
rect 240414 372535 240470 372544
rect 224224 371884 224276 371890
rect 224224 371826 224276 371832
rect 222108 371680 222160 371686
rect 222108 371622 222160 371628
rect 238128 371414 238156 372535
rect 239324 371618 239352 372535
rect 239312 371612 239364 371618
rect 239312 371554 239364 371560
rect 240428 371550 240456 372535
rect 241072 372094 241100 374070
rect 242898 373416 242954 373425
rect 242898 373351 242954 373360
rect 242912 373182 242940 373351
rect 242900 373176 242952 373182
rect 242900 373118 242952 373124
rect 247130 373144 247186 373153
rect 247130 373079 247186 373088
rect 241702 372600 241758 372609
rect 241702 372535 241758 372544
rect 244278 372600 244334 372609
rect 244278 372535 244334 372544
rect 241060 372088 241112 372094
rect 241060 372030 241112 372036
rect 241716 371754 241744 372535
rect 244292 372434 244320 372535
rect 244280 372428 244332 372434
rect 244280 372370 244332 372376
rect 247144 371890 247172 373079
rect 248418 372600 248474 372609
rect 248418 372535 248474 372544
rect 251178 372600 251234 372609
rect 251178 372535 251234 372544
rect 247132 371884 247184 371890
rect 247132 371826 247184 371832
rect 248432 371822 248460 372535
rect 248420 371816 248472 371822
rect 245658 371784 245714 371793
rect 241704 371748 241756 371754
rect 241704 371690 241756 371696
rect 242808 371748 242860 371754
rect 248420 371758 248472 371764
rect 245658 371719 245714 371728
rect 242808 371690 242860 371696
rect 242820 371550 242848 371690
rect 240416 371544 240468 371550
rect 240416 371486 240468 371492
rect 241428 371544 241480 371550
rect 241428 371486 241480 371492
rect 242808 371544 242860 371550
rect 242808 371486 242860 371492
rect 241440 371414 241468 371486
rect 238116 371408 238168 371414
rect 238116 371350 238168 371356
rect 241428 371408 241480 371414
rect 241428 371350 241480 371356
rect 245672 371346 245700 371719
rect 251192 371686 251220 372535
rect 251284 372026 251312 374439
rect 256068 374270 256096 374439
rect 256056 374264 256108 374270
rect 256056 374206 256108 374212
rect 270222 374096 270278 374105
rect 270222 374031 270278 374040
rect 262770 373824 262826 373833
rect 262770 373759 262826 373768
rect 255410 373552 255466 373561
rect 255410 373487 255466 373496
rect 256698 373552 256754 373561
rect 256698 373487 256754 373496
rect 253938 373144 253994 373153
rect 253938 373079 253940 373088
rect 253992 373079 253994 373088
rect 253940 373050 253992 373056
rect 255424 373046 255452 373487
rect 256712 373454 256740 373487
rect 256700 373448 256752 373454
rect 256700 373390 256752 373396
rect 260010 373416 260066 373425
rect 260010 373351 260012 373360
rect 260064 373351 260066 373360
rect 260012 373322 260064 373328
rect 258078 373144 258134 373153
rect 258078 373079 258134 373088
rect 261298 373144 261354 373153
rect 261298 373079 261354 373088
rect 255412 373040 255464 373046
rect 255412 372982 255464 372988
rect 258092 372910 258120 373079
rect 261312 372978 261340 373079
rect 261300 372972 261352 372978
rect 261300 372914 261352 372920
rect 258080 372904 258132 372910
rect 258080 372846 258132 372852
rect 259460 372836 259512 372842
rect 259460 372778 259512 372784
rect 252558 372736 252614 372745
rect 252558 372671 252614 372680
rect 251272 372020 251324 372026
rect 251272 371962 251324 371968
rect 252572 371958 252600 372671
rect 259472 372609 259500 372778
rect 262220 372768 262272 372774
rect 262220 372710 262272 372716
rect 262232 372609 262260 372710
rect 259458 372600 259514 372609
rect 259458 372535 259514 372544
rect 262218 372600 262274 372609
rect 262218 372535 262274 372544
rect 252560 371952 252612 371958
rect 252560 371894 252612 371900
rect 251180 371680 251232 371686
rect 262784 371657 262812 373759
rect 269210 373416 269266 373425
rect 269210 373351 269266 373360
rect 269224 373318 269252 373351
rect 262864 373312 262916 373318
rect 262864 373254 262916 373260
rect 269212 373312 269264 373318
rect 269212 373254 269264 373260
rect 262876 372337 262904 373254
rect 264978 373144 265034 373153
rect 264978 373079 265034 373088
rect 264992 372706 265020 373079
rect 264980 372700 265032 372706
rect 264980 372642 265032 372648
rect 266360 372632 266412 372638
rect 266358 372600 266360 372609
rect 266412 372600 266414 372609
rect 266358 372535 266414 372544
rect 262862 372328 262918 372337
rect 262862 372263 262918 372272
rect 270236 371929 270264 374031
rect 270512 372201 270540 374439
rect 271878 372600 271934 372609
rect 275296 372570 275324 374818
rect 295340 374808 295392 374814
rect 295340 374750 295392 374756
rect 271878 372535 271880 372544
rect 271932 372535 271934 372544
rect 275284 372564 275336 372570
rect 271880 372506 271932 372512
rect 275284 372506 275336 372512
rect 295352 372502 295380 374750
rect 305000 374740 305052 374746
rect 305000 374682 305052 374688
rect 300858 373144 300914 373153
rect 300858 373079 300914 373088
rect 295340 372496 295392 372502
rect 278686 372464 278742 372473
rect 295340 372438 295392 372444
rect 278686 372399 278742 372408
rect 276938 372328 276994 372337
rect 276938 372263 276994 372272
rect 270498 372192 270554 372201
rect 270498 372127 270554 372136
rect 270222 371920 270278 371929
rect 270222 371855 270278 371864
rect 273442 371784 273498 371793
rect 276952 371754 276980 372263
rect 278700 371822 278728 372399
rect 278688 371816 278740 371822
rect 278688 371758 278740 371764
rect 273442 371719 273498 371728
rect 276020 371748 276072 371754
rect 273352 371680 273404 371686
rect 251180 371622 251232 371628
rect 262770 371648 262826 371657
rect 273352 371622 273404 371628
rect 262770 371583 262826 371592
rect 247038 371376 247094 371385
rect 245660 371340 245712 371346
rect 247038 371311 247094 371320
rect 252558 371376 252614 371385
rect 252558 371311 252614 371320
rect 258170 371376 258226 371385
rect 258170 371311 258226 371320
rect 260838 371376 260894 371385
rect 260838 371311 260894 371320
rect 263598 371376 263654 371385
rect 263598 371311 263654 371320
rect 264978 371376 265034 371385
rect 264978 371311 265034 371320
rect 266358 371376 266414 371385
rect 266358 371311 266414 371320
rect 267738 371376 267794 371385
rect 267738 371311 267794 371320
rect 270498 371376 270554 371385
rect 270498 371311 270554 371320
rect 273258 371376 273314 371385
rect 273258 371311 273314 371320
rect 245660 371282 245712 371288
rect 247052 369102 247080 371311
rect 252572 369374 252600 371311
rect 252560 369368 252612 369374
rect 252560 369310 252612 369316
rect 258184 369170 258212 371311
rect 260852 369306 260880 371311
rect 260840 369300 260892 369306
rect 260840 369242 260892 369248
rect 263612 369238 263640 371311
rect 264992 369578 265020 371311
rect 264980 369572 265032 369578
rect 264980 369514 265032 369520
rect 263600 369232 263652 369238
rect 263600 369174 263652 369180
rect 258172 369164 258224 369170
rect 258172 369106 258224 369112
rect 247040 369096 247092 369102
rect 247040 369038 247092 369044
rect 266372 368393 266400 371311
rect 267752 369442 267780 371311
rect 270512 369782 270540 371311
rect 273272 371278 273300 371311
rect 273260 371272 273312 371278
rect 273260 371214 273312 371220
rect 273364 370394 273392 371622
rect 273352 370388 273404 370394
rect 273352 370330 273404 370336
rect 270500 369776 270552 369782
rect 270500 369718 270552 369724
rect 273456 369510 273484 371719
rect 276020 371690 276072 371696
rect 276940 371748 276992 371754
rect 276940 371690 276992 371696
rect 276032 371521 276060 371690
rect 276018 371512 276074 371521
rect 276018 371447 276074 371456
rect 277674 371512 277730 371521
rect 277674 371447 277730 371456
rect 276018 371376 276074 371385
rect 276018 371311 276074 371320
rect 276032 369646 276060 371311
rect 277688 370462 277716 371447
rect 280158 371376 280214 371385
rect 280158 371311 280214 371320
rect 282918 371376 282974 371385
rect 282918 371311 282974 371320
rect 285678 371376 285734 371385
rect 285678 371311 285734 371320
rect 287334 371376 287390 371385
rect 287334 371311 287390 371320
rect 289818 371376 289874 371385
rect 289818 371311 289874 371320
rect 292578 371376 292634 371385
rect 292578 371311 292634 371320
rect 295338 371376 295394 371385
rect 295338 371311 295394 371320
rect 298098 371376 298154 371385
rect 298098 371311 298154 371320
rect 277676 370456 277728 370462
rect 277676 370398 277728 370404
rect 280172 369714 280200 371311
rect 282932 370530 282960 371311
rect 285692 370598 285720 371311
rect 287348 370666 287376 371311
rect 289832 370734 289860 371311
rect 292592 370802 292620 371311
rect 295352 370938 295380 371311
rect 298112 371006 298140 371311
rect 300872 371142 300900 373079
rect 305012 372434 305040 374682
rect 312820 374672 312872 374678
rect 312820 374614 312872 374620
rect 310518 372600 310574 372609
rect 310518 372535 310574 372544
rect 310532 372502 310560 372535
rect 312832 372502 312860 374614
rect 320914 374504 320970 374513
rect 320914 374439 320916 374448
rect 320968 374439 320970 374448
rect 320916 374410 320968 374416
rect 314658 372600 314714 372609
rect 314658 372535 314660 372544
rect 314712 372535 314714 372544
rect 322938 372600 322994 372609
rect 322938 372535 322994 372544
rect 314660 372506 314712 372512
rect 322952 372502 322980 372535
rect 310520 372496 310572 372502
rect 310520 372438 310572 372444
rect 312820 372496 312872 372502
rect 322940 372496 322992 372502
rect 312820 372438 312872 372444
rect 313278 372464 313334 372473
rect 305000 372428 305052 372434
rect 322940 372438 322992 372444
rect 313278 372399 313280 372408
rect 305000 372370 305052 372376
rect 313332 372399 313334 372408
rect 313280 372370 313332 372376
rect 304998 372328 305054 372337
rect 304998 372263 305054 372272
rect 305012 371686 305040 372263
rect 356612 371816 356664 371822
rect 317418 371784 317474 371793
rect 356612 371758 356664 371764
rect 317418 371719 317474 371728
rect 305000 371680 305052 371686
rect 305000 371622 305052 371628
rect 302238 371376 302294 371385
rect 302238 371311 302294 371320
rect 307758 371376 307814 371385
rect 307758 371311 307814 371320
rect 302252 371210 302280 371311
rect 302240 371204 302292 371210
rect 302240 371146 302292 371152
rect 300860 371136 300912 371142
rect 300860 371078 300912 371084
rect 298100 371000 298152 371006
rect 298100 370942 298152 370948
rect 295340 370932 295392 370938
rect 295340 370874 295392 370880
rect 307772 370870 307800 371311
rect 317432 371074 317460 371719
rect 326158 371376 326214 371385
rect 342902 371376 342958 371385
rect 326158 371311 326214 371320
rect 342260 371340 342312 371346
rect 317420 371068 317472 371074
rect 317420 371010 317472 371016
rect 307760 370864 307812 370870
rect 307760 370806 307812 370812
rect 292580 370796 292632 370802
rect 292580 370738 292632 370744
rect 289820 370728 289872 370734
rect 289820 370670 289872 370676
rect 287336 370660 287388 370666
rect 287336 370602 287388 370608
rect 285680 370592 285732 370598
rect 285680 370534 285732 370540
rect 282920 370524 282972 370530
rect 282920 370466 282972 370472
rect 326172 369850 326200 371311
rect 342902 371311 342958 371320
rect 343362 371376 343418 371385
rect 343362 371311 343364 371320
rect 342260 371282 342312 371288
rect 326160 369844 326212 369850
rect 326160 369786 326212 369792
rect 280160 369708 280212 369714
rect 280160 369650 280212 369656
rect 276020 369640 276072 369646
rect 276020 369582 276072 369588
rect 273444 369504 273496 369510
rect 273444 369446 273496 369452
rect 267740 369436 267792 369442
rect 267740 369378 267792 369384
rect 342272 368490 342300 371282
rect 342916 371278 342944 371311
rect 343416 371311 343418 371320
rect 343364 371282 343416 371288
rect 342904 371272 342956 371278
rect 342904 371214 342956 371220
rect 342260 368484 342312 368490
rect 342260 368426 342312 368432
rect 266358 368384 266414 368393
rect 266358 368319 266414 368328
rect 342916 360874 342944 371214
rect 342904 360868 342956 360874
rect 342904 360810 342956 360816
rect 338488 355428 338540 355434
rect 338488 355370 338540 355376
rect 338500 355065 338528 355370
rect 351736 355360 351788 355366
rect 351736 355302 351788 355308
rect 351748 355065 351776 355302
rect 338486 355056 338542 355065
rect 338486 354991 338542 355000
rect 351734 355056 351790 355065
rect 351734 354991 351790 355000
rect 339774 354784 339830 354793
rect 339774 354719 339776 354728
rect 339828 354719 339830 354728
rect 339776 354690 339828 354696
rect 221096 353456 221148 353462
rect 221002 353424 221058 353433
rect 220912 353388 220964 353394
rect 221096 353398 221148 353404
rect 221002 353359 221058 353368
rect 220912 353330 220964 353336
rect 220820 353320 220872 353326
rect 220820 353262 220872 353268
rect 250718 269920 250774 269929
rect 250718 269855 250774 269864
rect 263506 269920 263562 269929
rect 263506 269855 263562 269864
rect 250732 269550 250760 269855
rect 263520 269618 263548 269855
rect 275742 269784 275798 269793
rect 275742 269719 275798 269728
rect 280894 269784 280950 269793
rect 280894 269719 280950 269728
rect 315854 269784 315910 269793
rect 315854 269719 315910 269728
rect 263508 269612 263560 269618
rect 263508 269554 263560 269560
rect 250720 269544 250772 269550
rect 250720 269486 250772 269492
rect 275756 269414 275784 269719
rect 279146 269648 279202 269657
rect 279146 269583 279202 269592
rect 279160 269482 279188 269583
rect 279148 269476 279200 269482
rect 279148 269418 279200 269424
rect 275744 269408 275796 269414
rect 275744 269350 275796 269356
rect 280908 269346 280936 269719
rect 283470 269648 283526 269657
rect 283470 269583 283526 269592
rect 285954 269648 286010 269657
rect 285954 269583 286010 269592
rect 288254 269648 288310 269657
rect 288254 269583 288310 269592
rect 293406 269648 293462 269657
rect 293406 269583 293462 269592
rect 308494 269648 308550 269657
rect 308494 269583 308550 269592
rect 280896 269340 280948 269346
rect 280896 269282 280948 269288
rect 283484 269278 283512 269583
rect 283472 269272 283524 269278
rect 283472 269214 283524 269220
rect 285968 269142 285996 269583
rect 288268 269210 288296 269583
rect 288256 269204 288308 269210
rect 288256 269146 288308 269152
rect 285956 269136 286008 269142
rect 285956 269078 286008 269084
rect 290922 268968 290978 268977
rect 290922 268903 290978 268912
rect 290936 268870 290964 268903
rect 290924 268864 290976 268870
rect 243082 268832 243138 268841
rect 243082 268767 243138 268776
rect 258078 268832 258134 268841
rect 258078 268767 258134 268776
rect 261666 268832 261722 268841
rect 290924 268806 290976 268812
rect 261666 268767 261722 268776
rect 236644 267980 236696 267986
rect 236644 267922 236696 267928
rect 220728 266008 220780 266014
rect 220726 265976 220728 265985
rect 220780 265976 220782 265985
rect 220726 265911 220782 265920
rect 230388 265124 230440 265130
rect 230388 265066 230440 265072
rect 230400 264790 230428 265066
rect 233148 265056 233200 265062
rect 233148 264998 233200 265004
rect 231768 264988 231820 264994
rect 231768 264930 231820 264936
rect 230388 264784 230440 264790
rect 230388 264726 230440 264732
rect 231780 264654 231808 264930
rect 233160 264722 233188 264998
rect 233148 264716 233200 264722
rect 233148 264658 233200 264664
rect 231768 264648 231820 264654
rect 231768 264590 231820 264596
rect 236656 251122 236684 267922
rect 243096 267918 243124 268767
rect 255780 267980 255832 267986
rect 255780 267922 255832 267928
rect 243084 267912 243136 267918
rect 243084 267854 243136 267860
rect 255792 267753 255820 267922
rect 258092 267850 258120 268767
rect 258080 267844 258132 267850
rect 258080 267786 258132 267792
rect 261680 267782 261708 268767
rect 293420 268734 293448 269583
rect 298466 269104 298522 269113
rect 298466 269039 298522 269048
rect 300858 269104 300914 269113
rect 300858 269039 300914 269048
rect 295890 268968 295946 268977
rect 295890 268903 295946 268912
rect 295904 268802 295932 268903
rect 295892 268796 295944 268802
rect 295892 268738 295944 268744
rect 293408 268728 293460 268734
rect 293408 268670 293460 268676
rect 298480 268598 298508 269039
rect 298468 268592 298520 268598
rect 298468 268534 298520 268540
rect 300872 268530 300900 269039
rect 308508 268666 308536 269583
rect 308496 268660 308548 268666
rect 308496 268602 308548 268608
rect 300860 268524 300912 268530
rect 300860 268466 300912 268472
rect 315868 268394 315896 269719
rect 318430 269648 318486 269657
rect 318430 269583 318486 269592
rect 318444 268462 318472 269583
rect 318432 268456 318484 268462
rect 318432 268398 318484 268404
rect 315856 268388 315908 268394
rect 315856 268330 315908 268336
rect 265162 268152 265218 268161
rect 265162 268087 265218 268096
rect 272154 268152 272210 268161
rect 272154 268087 272210 268096
rect 261668 267776 261720 267782
rect 255778 267744 255834 267753
rect 255778 267679 255834 267688
rect 260838 267744 260894 267753
rect 261668 267718 261720 267724
rect 263598 267744 263654 267753
rect 260838 267679 260894 267688
rect 263598 267679 263654 267688
rect 260852 267238 260880 267679
rect 263612 267306 263640 267679
rect 263600 267300 263652 267306
rect 263600 267242 263652 267248
rect 260840 267232 260892 267238
rect 258262 267200 258318 267209
rect 260840 267174 260892 267180
rect 258262 267135 258318 267144
rect 258276 267102 258304 267135
rect 258264 267096 258316 267102
rect 255318 267064 255374 267073
rect 258264 267038 258316 267044
rect 255318 266999 255374 267008
rect 255332 266966 255360 266999
rect 255320 266960 255372 266966
rect 247038 266928 247094 266937
rect 247038 266863 247094 266872
rect 252558 266928 252614 266937
rect 255320 266902 255372 266908
rect 263598 266928 263654 266937
rect 252558 266863 252560 266872
rect 247052 266830 247080 266863
rect 252612 266863 252614 266872
rect 263598 266863 263654 266872
rect 252560 266834 252612 266840
rect 247040 266824 247092 266830
rect 247040 266766 247092 266772
rect 244370 266520 244426 266529
rect 244370 266455 244426 266464
rect 251270 266520 251326 266529
rect 251270 266455 251326 266464
rect 259550 266520 259606 266529
rect 259550 266455 259606 266464
rect 244278 266384 244334 266393
rect 244278 266319 244334 266328
rect 244292 265878 244320 266319
rect 244280 265872 244332 265878
rect 244280 265814 244332 265820
rect 244384 264382 244412 266455
rect 245658 266384 245714 266393
rect 245658 266319 245714 266328
rect 247038 266384 247094 266393
rect 247038 266319 247094 266328
rect 248510 266384 248566 266393
rect 248510 266319 248566 266328
rect 249798 266384 249854 266393
rect 249798 266319 249854 266328
rect 251178 266384 251234 266393
rect 251178 266319 251234 266328
rect 245672 266150 245700 266319
rect 245660 266144 245712 266150
rect 245660 266086 245712 266092
rect 247052 265810 247080 266319
rect 248524 265946 248552 266319
rect 249812 266014 249840 266319
rect 251192 266082 251220 266319
rect 251284 266218 251312 266455
rect 252558 266384 252614 266393
rect 252558 266319 252614 266328
rect 253938 266384 253994 266393
rect 253938 266319 253994 266328
rect 256698 266384 256754 266393
rect 256698 266319 256754 266328
rect 259458 266384 259514 266393
rect 259458 266319 259514 266328
rect 252572 266286 252600 266319
rect 252560 266280 252612 266286
rect 252560 266222 252612 266228
rect 251272 266212 251324 266218
rect 251272 266154 251324 266160
rect 251180 266076 251232 266082
rect 251180 266018 251232 266024
rect 249800 266008 249852 266014
rect 249800 265950 249852 265956
rect 248512 265940 248564 265946
rect 248512 265882 248564 265888
rect 247040 265804 247092 265810
rect 247040 265746 247092 265752
rect 253952 264858 253980 266319
rect 253940 264852 253992 264858
rect 253940 264794 253992 264800
rect 256712 264654 256740 266319
rect 259472 264722 259500 266319
rect 259564 264790 259592 266455
rect 262218 266384 262274 266393
rect 262218 266319 262220 266328
rect 262272 266319 262274 266328
rect 262220 266290 262272 266296
rect 259552 264784 259604 264790
rect 259552 264726 259604 264732
rect 259460 264716 259512 264722
rect 259460 264658 259512 264664
rect 256700 264648 256752 264654
rect 256700 264590 256752 264596
rect 244372 264376 244424 264382
rect 244372 264318 244424 264324
rect 263612 251190 263640 266863
rect 265176 265742 265204 268087
rect 265806 267744 265862 267753
rect 265806 267679 265862 267688
rect 267094 267744 267150 267753
rect 267094 267679 267150 267688
rect 268198 267744 268254 267753
rect 268198 267679 268254 267688
rect 270866 267744 270922 267753
rect 270866 267679 270922 267688
rect 265820 267170 265848 267679
rect 265808 267164 265860 267170
rect 265808 267106 265860 267112
rect 265164 265736 265216 265742
rect 265164 265678 265216 265684
rect 267108 265674 267136 267679
rect 268212 267442 268240 267679
rect 270880 267510 270908 267679
rect 270868 267504 270920 267510
rect 270868 267446 270920 267452
rect 268200 267436 268252 267442
rect 268200 267378 268252 267384
rect 269762 267200 269818 267209
rect 269762 267135 269818 267144
rect 271234 267200 271290 267209
rect 271234 267135 271290 267144
rect 267738 266928 267794 266937
rect 267738 266863 267794 266872
rect 267096 265668 267148 265674
rect 267096 265610 267148 265616
rect 263600 251184 263652 251190
rect 263600 251126 263652 251132
rect 236644 251116 236696 251122
rect 236644 251058 236696 251064
rect 267752 250510 267780 266863
rect 269776 264314 269804 267135
rect 269764 264308 269816 264314
rect 269764 264250 269816 264256
rect 271248 264246 271276 267135
rect 272168 264926 272196 268087
rect 356520 267980 356572 267986
rect 356520 267922 356572 267928
rect 273258 267744 273314 267753
rect 273258 267679 273314 267688
rect 276018 267744 276074 267753
rect 276018 267679 276074 267688
rect 302238 267744 302294 267753
rect 302238 267679 302294 267688
rect 273272 267374 273300 267679
rect 276032 267578 276060 267679
rect 302252 267646 302280 267679
rect 302240 267640 302292 267646
rect 302240 267582 302292 267588
rect 276020 267572 276072 267578
rect 276020 267514 276072 267520
rect 343454 267472 343510 267481
rect 343454 267407 343510 267416
rect 273260 267368 273312 267374
rect 273260 267310 273312 267316
rect 343468 267238 343496 267407
rect 356532 267374 356560 267922
rect 356520 267368 356572 267374
rect 343546 267336 343602 267345
rect 356520 267310 356572 267316
rect 343546 267271 343602 267280
rect 343456 267232 343508 267238
rect 277122 267200 277178 267209
rect 277122 267135 277178 267144
rect 278134 267200 278190 267209
rect 343456 267174 343508 267180
rect 278134 267135 278136 267144
rect 273258 267064 273314 267073
rect 277136 267034 277164 267135
rect 278188 267135 278190 267144
rect 278136 267106 278188 267112
rect 343560 267102 343588 267271
rect 356520 267232 356572 267238
rect 356520 267174 356572 267180
rect 343548 267096 343600 267102
rect 343548 267038 343600 267044
rect 356532 267034 356560 267174
rect 356624 267170 356652 371758
rect 356612 267164 356664 267170
rect 356612 267106 356664 267112
rect 273258 266999 273260 267008
rect 273312 266999 273314 267008
rect 277124 267028 277176 267034
rect 273260 266970 273312 266976
rect 277124 266970 277176 266976
rect 356520 267028 356572 267034
rect 356520 266970 356572 266976
rect 310518 266928 310574 266937
rect 310518 266863 310574 266872
rect 310532 266762 310560 266863
rect 310520 266756 310572 266762
rect 310520 266698 310572 266704
rect 279974 266384 280030 266393
rect 279974 266319 280030 266328
rect 272156 264920 272208 264926
rect 272156 264862 272208 264868
rect 271236 264240 271288 264246
rect 271236 264182 271288 264188
rect 279988 250510 280016 266319
rect 356532 258074 356560 266970
rect 356624 266422 356652 267106
rect 356612 266416 356664 266422
rect 356612 266358 356664 266364
rect 356532 258046 356652 258074
rect 340236 251184 340288 251190
rect 340236 251126 340288 251132
rect 338488 250572 338540 250578
rect 338488 250514 338540 250520
rect 267740 250504 267792 250510
rect 267740 250446 267792 250452
rect 279976 250504 280028 250510
rect 279976 250446 280028 250452
rect 338500 249937 338528 250514
rect 340248 249937 340276 251126
rect 338486 249928 338542 249937
rect 338486 249863 338542 249872
rect 340234 249928 340290 249937
rect 340234 249863 340290 249872
rect 350998 249928 351054 249937
rect 350998 249863 351054 249872
rect 351012 249830 351040 249863
rect 351000 249824 351052 249830
rect 351000 249766 351052 249772
rect 258446 164792 258502 164801
rect 258446 164727 258502 164736
rect 282182 164792 282238 164801
rect 282182 164727 282238 164736
rect 249154 164520 249210 164529
rect 249154 164455 249210 164464
rect 249168 164257 249196 164455
rect 258460 164354 258488 164727
rect 261022 164656 261078 164665
rect 261022 164591 261078 164600
rect 276110 164656 276166 164665
rect 276110 164591 276166 164600
rect 258448 164348 258500 164354
rect 258448 164290 258500 164296
rect 249154 164248 249210 164257
rect 249154 164183 249210 164192
rect 261036 163742 261064 164591
rect 262862 164520 262918 164529
rect 262862 164455 262918 164464
rect 262876 164257 262904 164455
rect 262862 164248 262918 164257
rect 262862 164183 262918 164192
rect 261024 163736 261076 163742
rect 261024 163678 261076 163684
rect 235998 163160 236054 163169
rect 235998 163095 236054 163104
rect 264978 163160 265034 163169
rect 264978 163095 265034 163104
rect 224144 145858 224356 145874
rect 224144 145852 224368 145858
rect 224144 145846 224316 145852
rect 224144 145722 224172 145846
rect 224316 145794 224368 145800
rect 224132 145716 224184 145722
rect 224132 145658 224184 145664
rect 224224 145716 224276 145722
rect 224224 145658 224276 145664
rect 224236 145246 224264 145658
rect 236012 145382 236040 163095
rect 236090 162752 236146 162761
rect 236090 162687 236146 162696
rect 237378 162752 237434 162761
rect 237378 162687 237434 162696
rect 240138 162752 240194 162761
rect 240138 162687 240194 162696
rect 241518 162752 241574 162761
rect 241518 162687 241574 162696
rect 242898 162752 242954 162761
rect 242898 162687 242954 162696
rect 244278 162752 244334 162761
rect 244278 162687 244334 162696
rect 245658 162752 245714 162761
rect 245658 162687 245714 162696
rect 247130 162752 247186 162761
rect 247130 162687 247186 162696
rect 247866 162752 247922 162761
rect 247866 162687 247922 162696
rect 248418 162752 248474 162761
rect 248418 162687 248474 162696
rect 249798 162752 249854 162761
rect 249798 162687 249854 162696
rect 251270 162752 251326 162761
rect 251270 162687 251326 162696
rect 252558 162752 252614 162761
rect 252558 162687 252614 162696
rect 253938 162752 253994 162761
rect 253938 162687 253994 162696
rect 255410 162752 255466 162761
rect 255410 162687 255466 162696
rect 255962 162752 256018 162761
rect 255962 162687 256018 162696
rect 256698 162752 256754 162761
rect 256698 162687 256754 162696
rect 259550 162752 259606 162761
rect 259550 162687 259606 162696
rect 260838 162752 260894 162761
rect 260838 162687 260894 162696
rect 262218 162752 262274 162761
rect 262218 162687 262274 162696
rect 263598 162752 263654 162761
rect 263598 162687 263654 162696
rect 236104 145450 236132 162687
rect 237392 145897 237420 162687
rect 238758 161528 238814 161537
rect 238758 161463 238814 161472
rect 238772 148374 238800 161463
rect 240152 148850 240180 162687
rect 241532 148918 241560 162687
rect 241520 148912 241572 148918
rect 241520 148854 241572 148860
rect 240140 148844 240192 148850
rect 240140 148786 240192 148792
rect 238760 148368 238812 148374
rect 238760 148310 238812 148316
rect 237378 145888 237434 145897
rect 237378 145823 237434 145832
rect 242912 145518 242940 162687
rect 244292 145722 244320 162687
rect 244370 162208 244426 162217
rect 244370 162143 244426 162152
rect 244280 145716 244332 145722
rect 244280 145658 244332 145664
rect 244384 145654 244412 162143
rect 244372 145648 244424 145654
rect 244372 145590 244424 145596
rect 245672 145586 245700 162687
rect 247144 145858 247172 162687
rect 247880 161974 247908 162687
rect 247868 161968 247920 161974
rect 247868 161910 247920 161916
rect 247132 145852 247184 145858
rect 247132 145794 247184 145800
rect 248432 145790 248460 162687
rect 249812 145926 249840 162687
rect 251178 162480 251234 162489
rect 251178 162415 251234 162424
rect 251192 146062 251220 162415
rect 251180 146056 251232 146062
rect 251180 145998 251232 146004
rect 251284 145994 251312 162687
rect 252572 146130 252600 162687
rect 253952 146198 253980 162687
rect 255424 146266 255452 162687
rect 255976 162110 256004 162687
rect 255964 162104 256016 162110
rect 255964 162046 256016 162052
rect 256712 159390 256740 162687
rect 259458 162616 259514 162625
rect 259458 162551 259514 162560
rect 258078 162208 258134 162217
rect 258078 162143 258134 162152
rect 258092 161090 258120 162143
rect 258080 161084 258132 161090
rect 258080 161026 258132 161032
rect 259472 160070 259500 162551
rect 259460 160064 259512 160070
rect 259460 160006 259512 160012
rect 259564 160002 259592 162687
rect 260852 161158 260880 162687
rect 260840 161152 260892 161158
rect 260840 161094 260892 161100
rect 262232 160818 262260 162687
rect 263612 161362 263640 162687
rect 263690 162616 263746 162625
rect 263690 162551 263746 162560
rect 263704 162042 263732 162551
rect 263692 162036 263744 162042
rect 263692 161978 263744 161984
rect 263600 161356 263652 161362
rect 263600 161298 263652 161304
rect 264992 161226 265020 163095
rect 267556 162920 267608 162926
rect 267556 162862 267608 162868
rect 267568 162761 267596 162862
rect 265438 162752 265494 162761
rect 265438 162687 265494 162696
rect 266358 162752 266414 162761
rect 266358 162687 266414 162696
rect 267554 162752 267610 162761
rect 267554 162687 267610 162696
rect 267738 162752 267794 162761
rect 267738 162687 267794 162696
rect 269118 162752 269174 162761
rect 269118 162687 269174 162696
rect 270498 162752 270554 162761
rect 270498 162687 270554 162696
rect 271878 162752 271934 162761
rect 271878 162687 271934 162696
rect 273258 162752 273314 162761
rect 273258 162687 273314 162696
rect 276018 162752 276074 162761
rect 276018 162687 276074 162696
rect 265452 162178 265480 162687
rect 265440 162172 265492 162178
rect 265440 162114 265492 162120
rect 266372 161294 266400 162687
rect 267752 161430 267780 162687
rect 268290 162616 268346 162625
rect 268290 162551 268346 162560
rect 268304 162382 268332 162551
rect 268292 162376 268344 162382
rect 268292 162318 268344 162324
rect 267740 161424 267792 161430
rect 267740 161366 267792 161372
rect 266360 161288 266412 161294
rect 266360 161230 266412 161236
rect 264980 161220 265032 161226
rect 264980 161162 265032 161168
rect 262220 160812 262272 160818
rect 262220 160754 262272 160760
rect 259552 159996 259604 160002
rect 259552 159938 259604 159944
rect 256700 159384 256752 159390
rect 256700 159326 256752 159332
rect 269132 146305 269160 162687
rect 269118 146296 269174 146305
rect 255412 146260 255464 146266
rect 269118 146231 269174 146240
rect 255412 146202 255464 146208
rect 253940 146192 253992 146198
rect 253940 146134 253992 146140
rect 252560 146124 252612 146130
rect 252560 146066 252612 146072
rect 251272 145988 251324 145994
rect 251272 145930 251324 145936
rect 249800 145920 249852 145926
rect 249800 145862 249852 145868
rect 248420 145784 248472 145790
rect 270512 145761 270540 162687
rect 248420 145726 248472 145732
rect 270498 145752 270554 145761
rect 270498 145687 270554 145696
rect 271892 145625 271920 162687
rect 273272 160750 273300 162687
rect 274546 162616 274602 162625
rect 274546 162551 274602 162560
rect 273442 162344 273498 162353
rect 273442 162279 273498 162288
rect 273456 162246 273484 162279
rect 273444 162240 273496 162246
rect 273444 162182 273496 162188
rect 274560 161474 274588 162551
rect 274560 161446 274772 161474
rect 273260 160744 273312 160750
rect 273260 160686 273312 160692
rect 274744 148986 274772 161446
rect 274732 148980 274784 148986
rect 274732 148922 274784 148928
rect 276032 146441 276060 162687
rect 276124 149054 276152 164591
rect 282196 164257 282224 164727
rect 305918 164656 305974 164665
rect 305918 164591 305974 164600
rect 318430 164656 318486 164665
rect 318430 164591 318486 164600
rect 282182 164248 282238 164257
rect 282182 164183 282238 164192
rect 298466 164248 298522 164257
rect 298466 164183 298522 164192
rect 300858 164248 300914 164257
rect 300858 164183 300914 164192
rect 298480 163674 298508 164183
rect 298468 163668 298520 163674
rect 298468 163610 298520 163616
rect 300872 163538 300900 164183
rect 305932 163606 305960 164591
rect 318444 164286 318472 164591
rect 318432 164280 318484 164286
rect 318432 164222 318484 164228
rect 305920 163600 305972 163606
rect 305920 163542 305972 163548
rect 300860 163532 300912 163538
rect 300860 163474 300912 163480
rect 320916 162852 320968 162858
rect 320916 162794 320968 162800
rect 308588 162784 308640 162790
rect 278410 162752 278466 162761
rect 278410 162687 278466 162696
rect 280066 162752 280122 162761
rect 280066 162687 280122 162696
rect 280802 162752 280858 162761
rect 280802 162687 280858 162696
rect 283746 162752 283802 162761
rect 283746 162687 283802 162696
rect 285954 162752 286010 162761
rect 285954 162687 286010 162696
rect 293314 162752 293370 162761
rect 293314 162687 293370 162696
rect 303434 162752 303490 162761
rect 303434 162687 303436 162696
rect 278424 162450 278452 162687
rect 278412 162444 278464 162450
rect 278412 162386 278464 162392
rect 278042 161528 278098 161537
rect 278042 161463 278098 161472
rect 278056 151814 278084 161463
rect 278056 151786 278268 151814
rect 276112 149048 276164 149054
rect 278240 149025 278268 151786
rect 276112 148990 276164 148996
rect 278226 149016 278282 149025
rect 278226 148951 278282 148960
rect 278240 148345 278268 148951
rect 278226 148336 278282 148345
rect 278226 148271 278282 148280
rect 276018 146432 276074 146441
rect 276018 146367 276074 146376
rect 276032 146266 276060 146367
rect 276020 146260 276072 146266
rect 276020 146202 276072 146208
rect 280080 145654 280108 162687
rect 280816 162314 280844 162687
rect 283760 162586 283788 162687
rect 283748 162580 283800 162586
rect 283748 162522 283800 162528
rect 285968 162518 285996 162687
rect 293328 162654 293356 162687
rect 303488 162687 303490 162696
rect 308586 162752 308588 162761
rect 308640 162752 308642 162761
rect 308586 162687 308642 162696
rect 303436 162658 303488 162664
rect 293316 162648 293368 162654
rect 320928 162625 320956 162794
rect 343454 162752 343510 162761
rect 343454 162687 343510 162696
rect 293316 162590 293368 162596
rect 320914 162616 320970 162625
rect 320914 162551 320970 162560
rect 343362 162616 343418 162625
rect 343362 162551 343418 162560
rect 285956 162512 286008 162518
rect 285956 162454 286008 162460
rect 280804 162308 280856 162314
rect 280804 162250 280856 162256
rect 343376 162178 343404 162551
rect 343468 162314 343496 162687
rect 343456 162308 343508 162314
rect 343456 162250 343508 162256
rect 343364 162172 343416 162178
rect 343364 162114 343416 162120
rect 356624 146266 356652 258046
rect 356716 163946 356744 478654
rect 362316 478644 362368 478650
rect 362316 478586 362368 478592
rect 360844 478508 360896 478514
rect 360844 478450 360896 478456
rect 358176 478372 358228 478378
rect 358176 478314 358228 478320
rect 356888 473068 356940 473074
rect 356888 473010 356940 473016
rect 356796 471708 356848 471714
rect 356796 471650 356848 471656
rect 356808 269113 356836 471650
rect 356900 374746 356928 473010
rect 358084 472728 358136 472734
rect 358084 472670 358136 472676
rect 356980 470348 357032 470354
rect 356980 470290 357032 470296
rect 356888 374740 356940 374746
rect 356888 374682 356940 374688
rect 356888 371748 356940 371754
rect 356888 371690 356940 371696
rect 356794 269104 356850 269113
rect 356794 269039 356850 269048
rect 356900 267238 356928 371690
rect 356992 371210 357020 470290
rect 357072 467764 357124 467770
rect 357072 467706 357124 467712
rect 356980 371204 357032 371210
rect 356980 371146 357032 371152
rect 357084 370530 357112 467706
rect 357992 464772 358044 464778
rect 357992 464714 358044 464720
rect 357440 461100 357492 461106
rect 357440 461042 357492 461048
rect 357164 460012 357216 460018
rect 357164 459954 357216 459960
rect 357176 372094 357204 459954
rect 357164 372088 357216 372094
rect 357164 372030 357216 372036
rect 357256 371272 357308 371278
rect 357256 371214 357308 371220
rect 357072 370524 357124 370530
rect 357072 370466 357124 370472
rect 357268 267714 357296 371214
rect 357348 356040 357400 356046
rect 357348 355982 357400 355988
rect 357360 354754 357388 355982
rect 357452 355434 357480 461042
rect 358004 406434 358032 464714
rect 357992 406428 358044 406434
rect 357992 406370 358044 406376
rect 357440 355428 357492 355434
rect 357440 355370 357492 355376
rect 357348 354748 357400 354754
rect 357348 354690 357400 354696
rect 357256 267708 357308 267714
rect 357256 267650 357308 267656
rect 356980 267368 357032 267374
rect 356980 267310 357032 267316
rect 356888 267232 356940 267238
rect 356888 267174 356940 267180
rect 356796 266416 356848 266422
rect 356796 266358 356848 266364
rect 356704 163940 356756 163946
rect 356704 163882 356756 163888
rect 356704 162852 356756 162858
rect 356704 162794 356756 162800
rect 356716 162314 356744 162794
rect 356704 162308 356756 162314
rect 356704 162250 356756 162256
rect 356612 146260 356664 146266
rect 356612 146202 356664 146208
rect 338488 146192 338540 146198
rect 338488 146134 338540 146140
rect 280068 145648 280120 145654
rect 271878 145616 271934 145625
rect 245660 145580 245712 145586
rect 280068 145590 280120 145596
rect 271878 145551 271934 145560
rect 245660 145522 245712 145528
rect 242900 145512 242952 145518
rect 242900 145454 242952 145460
rect 236092 145444 236144 145450
rect 236092 145386 236144 145392
rect 236000 145376 236052 145382
rect 236000 145318 236052 145324
rect 224224 145240 224276 145246
rect 224224 145182 224276 145188
rect 338500 144945 338528 146134
rect 340236 146124 340288 146130
rect 340236 146066 340288 146072
rect 340248 144945 340276 146066
rect 356612 145648 356664 145654
rect 356612 145590 356664 145596
rect 351644 145580 351696 145586
rect 351644 145522 351696 145528
rect 351656 144945 351684 145522
rect 338486 144936 338542 144945
rect 338486 144871 338542 144880
rect 340234 144936 340290 144945
rect 340234 144871 340290 144880
rect 351642 144936 351698 144945
rect 351642 144871 351698 144880
rect 237102 59800 237158 59809
rect 237102 59735 237104 59744
rect 237156 59735 237158 59744
rect 255870 59800 255926 59809
rect 255870 59735 255926 59744
rect 259458 59800 259514 59809
rect 259458 59735 259514 59744
rect 260654 59800 260710 59809
rect 260654 59735 260710 59744
rect 261758 59800 261814 59809
rect 261758 59735 261814 59744
rect 263874 59800 263930 59809
rect 263874 59735 263930 59744
rect 237104 59706 237156 59712
rect 255884 59702 255912 59735
rect 255872 59696 255924 59702
rect 255872 59638 255924 59644
rect 256974 59664 257030 59673
rect 256974 59599 257030 59608
rect 258078 59664 258134 59673
rect 258078 59599 258134 59608
rect 256988 59294 257016 59599
rect 256976 59288 257028 59294
rect 256976 59230 257028 59236
rect 258092 59226 258120 59599
rect 259472 59498 259500 59735
rect 260668 59566 260696 59735
rect 261772 59634 261800 59735
rect 261760 59628 261812 59634
rect 261760 59570 261812 59576
rect 260656 59560 260708 59566
rect 260656 59502 260708 59508
rect 262770 59528 262826 59537
rect 259460 59492 259512 59498
rect 262770 59463 262826 59472
rect 259460 59434 259512 59440
rect 258080 59220 258132 59226
rect 258080 59162 258132 59168
rect 262784 59090 262812 59463
rect 263888 59430 263916 59735
rect 265254 59664 265310 59673
rect 265254 59599 265310 59608
rect 315854 59664 315910 59673
rect 315854 59599 315910 59608
rect 263876 59424 263928 59430
rect 263876 59366 263928 59372
rect 265268 59158 265296 59599
rect 295890 59256 295946 59265
rect 295890 59191 295946 59200
rect 298466 59256 298522 59265
rect 298466 59191 298522 59200
rect 303434 59256 303490 59265
rect 303434 59191 303490 59200
rect 265256 59152 265308 59158
rect 265256 59094 265308 59100
rect 262772 59084 262824 59090
rect 262772 59026 262824 59032
rect 295904 59022 295932 59191
rect 295892 59016 295944 59022
rect 295892 58958 295944 58964
rect 298480 58886 298508 59191
rect 303448 58954 303476 59191
rect 303436 58948 303488 58954
rect 303436 58890 303488 58896
rect 298468 58880 298520 58886
rect 298468 58822 298520 58828
rect 315868 58818 315896 59599
rect 323306 59256 323362 59265
rect 323306 59191 323362 59200
rect 315856 58812 315908 58818
rect 315856 58754 315908 58760
rect 323320 58750 323348 59191
rect 323308 58744 323360 58750
rect 323308 58686 323360 58692
rect 325882 58168 325938 58177
rect 325882 58103 325938 58112
rect 325896 57934 325924 58103
rect 325884 57928 325936 57934
rect 235998 57896 236054 57905
rect 235998 57831 236054 57840
rect 237378 57896 237434 57905
rect 237378 57831 237434 57840
rect 239218 57896 239274 57905
rect 239218 57831 239274 57840
rect 242898 57896 242954 57905
rect 242898 57831 242954 57840
rect 244370 57896 244426 57905
rect 244370 57831 244426 57840
rect 246394 57896 246450 57905
rect 246394 57831 246450 57840
rect 248602 57896 248658 57905
rect 248602 57831 248658 57840
rect 251178 57896 251234 57905
rect 251178 57831 251234 57840
rect 253386 57896 253442 57905
rect 253386 57831 253442 57840
rect 265346 57896 265402 57905
rect 265346 57831 265402 57840
rect 266358 57896 266414 57905
rect 266358 57831 266414 57840
rect 267002 57896 267058 57905
rect 267002 57831 267058 57840
rect 269762 57896 269818 57905
rect 269762 57831 269818 57840
rect 272154 57896 272210 57905
rect 272154 57831 272210 57840
rect 273626 57896 273682 57905
rect 273626 57831 273682 57840
rect 274638 57896 274694 57905
rect 274638 57831 274694 57840
rect 279054 57896 279110 57905
rect 279054 57831 279110 57840
rect 283654 57896 283710 57905
rect 283654 57831 283710 57840
rect 287610 57896 287666 57905
rect 287610 57831 287666 57840
rect 293314 57896 293370 57905
rect 293314 57831 293370 57840
rect 300858 57896 300914 57905
rect 300858 57831 300914 57840
rect 305826 57896 305882 57905
rect 305826 57831 305882 57840
rect 310978 57896 311034 57905
rect 310978 57831 311034 57840
rect 313370 57896 313426 57905
rect 313370 57831 313426 57840
rect 318338 57896 318394 57905
rect 318338 57831 318340 57840
rect 236012 56438 236040 57831
rect 236000 56432 236052 56438
rect 236000 56374 236052 56380
rect 219992 55820 220044 55826
rect 219992 55762 220044 55768
rect 219900 54936 219952 54942
rect 219900 54878 219952 54884
rect 217876 54868 217928 54874
rect 217876 54810 217928 54816
rect 216312 54596 216364 54602
rect 216312 54538 216364 54544
rect 237392 54466 237420 57831
rect 239232 56506 239260 57831
rect 240138 57488 240194 57497
rect 240138 57423 240194 57432
rect 241518 57488 241574 57497
rect 241518 57423 241574 57432
rect 239862 57352 239918 57361
rect 239862 57287 239918 57296
rect 239876 56953 239904 57287
rect 239862 56944 239918 56953
rect 239862 56879 239918 56888
rect 239220 56500 239272 56506
rect 239220 56442 239272 56448
rect 240152 54534 240180 57423
rect 241532 54738 241560 57423
rect 242912 56574 242940 57831
rect 244278 57488 244334 57497
rect 244278 57423 244334 57432
rect 242900 56568 242952 56574
rect 242900 56510 242952 56516
rect 241520 54732 241572 54738
rect 241520 54674 241572 54680
rect 244292 54670 244320 57423
rect 244280 54664 244332 54670
rect 244280 54606 244332 54612
rect 244384 54602 244412 57831
rect 246408 56030 246436 57831
rect 247038 57488 247094 57497
rect 247038 57423 247094 57432
rect 246396 56024 246448 56030
rect 246396 55966 246448 55972
rect 247052 54806 247080 57423
rect 248616 55962 248644 57831
rect 249798 57488 249854 57497
rect 249798 57423 249854 57432
rect 248604 55956 248656 55962
rect 248604 55898 248656 55904
rect 249812 54913 249840 57423
rect 251192 56098 251220 57831
rect 251362 57488 251418 57497
rect 251362 57423 251418 57432
rect 251180 56092 251232 56098
rect 251180 56034 251232 56040
rect 249798 54904 249854 54913
rect 251376 54874 251404 57423
rect 253400 56166 253428 57831
rect 253938 57488 253994 57497
rect 253938 57423 253994 57432
rect 253388 56160 253440 56166
rect 253388 56102 253440 56108
rect 253952 54942 253980 57423
rect 265360 57254 265388 57831
rect 265348 57248 265400 57254
rect 265348 57190 265400 57196
rect 266372 56234 266400 57831
rect 267016 56302 267044 57831
rect 267738 57624 267794 57633
rect 267738 57559 267794 57568
rect 267004 56296 267056 56302
rect 267004 56238 267056 56244
rect 266360 56228 266412 56234
rect 266360 56170 266412 56176
rect 267752 55010 267780 57559
rect 269776 56370 269804 57831
rect 270498 57624 270554 57633
rect 270498 57559 270554 57568
rect 269764 56364 269816 56370
rect 269764 56306 269816 56312
rect 270512 55078 270540 57559
rect 272168 55758 272196 57831
rect 273350 57624 273406 57633
rect 273350 57559 273406 57568
rect 272156 55752 272208 55758
rect 272156 55694 272208 55700
rect 273364 55146 273392 57559
rect 273640 55894 273668 57831
rect 273628 55888 273680 55894
rect 273628 55830 273680 55836
rect 274652 55214 274680 57831
rect 277398 57624 277454 57633
rect 277398 57559 277454 57568
rect 274640 55208 274692 55214
rect 274640 55150 274692 55156
rect 273352 55140 273404 55146
rect 273352 55082 273404 55088
rect 270500 55072 270552 55078
rect 277412 55049 277440 57559
rect 279068 57458 279096 57831
rect 279056 57452 279108 57458
rect 279056 57394 279108 57400
rect 283668 57186 283696 57831
rect 287624 57322 287652 57831
rect 293328 57390 293356 57831
rect 300872 57526 300900 57831
rect 305840 57594 305868 57831
rect 310992 57798 311020 57831
rect 310980 57792 311032 57798
rect 310980 57734 311032 57740
rect 313384 57662 313412 57831
rect 318392 57831 318394 57840
rect 320914 57896 320970 57905
rect 343180 57928 343232 57934
rect 325884 57870 325936 57876
rect 343178 57896 343180 57905
rect 343232 57896 343234 57905
rect 320914 57831 320970 57840
rect 343178 57831 343234 57840
rect 343454 57896 343510 57905
rect 343454 57831 343456 57840
rect 318340 57802 318392 57808
rect 320928 57730 320956 57831
rect 343508 57831 343510 57840
rect 343456 57802 343508 57808
rect 320916 57724 320968 57730
rect 320916 57666 320968 57672
rect 313372 57656 313424 57662
rect 307758 57624 307814 57633
rect 305828 57588 305880 57594
rect 313372 57598 313424 57604
rect 307758 57559 307814 57568
rect 305828 57530 305880 57536
rect 300860 57520 300912 57526
rect 300860 57462 300912 57468
rect 293316 57384 293368 57390
rect 293316 57326 293368 57332
rect 287612 57316 287664 57322
rect 287612 57258 287664 57264
rect 283656 57180 283708 57186
rect 283656 57122 283708 57128
rect 307772 55185 307800 57559
rect 356624 57458 356652 145590
rect 356716 57866 356744 162250
rect 356808 149025 356836 266358
rect 356888 252544 356940 252550
rect 356888 252486 356940 252492
rect 356900 250578 356928 252486
rect 356888 250572 356940 250578
rect 356888 250514 356940 250520
rect 356794 149016 356850 149025
rect 356794 148951 356850 148960
rect 356900 146198 356928 250514
rect 356992 162858 357020 267310
rect 357360 252498 357388 354690
rect 357452 252618 357480 355370
rect 357532 267708 357584 267714
rect 357532 267650 357584 267656
rect 357544 267102 357572 267650
rect 357532 267096 357584 267102
rect 357532 267038 357584 267044
rect 357440 252612 357492 252618
rect 357440 252554 357492 252560
rect 357360 252470 357480 252498
rect 357452 251258 357480 252470
rect 357440 251252 357492 251258
rect 357440 251194 357492 251200
rect 356980 162852 357032 162858
rect 356980 162794 357032 162800
rect 356888 146192 356940 146198
rect 356888 146134 356940 146140
rect 357452 146130 357480 251194
rect 357544 162178 357572 267038
rect 357624 250504 357676 250510
rect 357624 250446 357676 250452
rect 357532 162172 357584 162178
rect 357532 162114 357584 162120
rect 357440 146124 357492 146130
rect 357440 146066 357492 146072
rect 357544 57934 357572 162114
rect 357636 145654 357664 250446
rect 358096 162178 358124 472670
rect 358084 162172 358136 162178
rect 358084 162114 358136 162120
rect 357624 145648 357676 145654
rect 357624 145590 357676 145596
rect 358084 68196 358136 68202
rect 358084 68138 358136 68144
rect 358096 59362 358124 68138
rect 358188 59430 358216 478314
rect 359740 477284 359792 477290
rect 359740 477226 359792 477232
rect 359464 475856 359516 475862
rect 359464 475798 359516 475804
rect 358452 471844 358504 471850
rect 358452 471786 358504 471792
rect 358360 471572 358412 471578
rect 358360 471514 358412 471520
rect 358268 467220 358320 467226
rect 358268 467162 358320 467168
rect 358280 162110 358308 467162
rect 358372 267374 358400 471514
rect 358464 369646 358492 471786
rect 358544 464908 358596 464914
rect 358544 464850 358596 464856
rect 358452 369640 358504 369646
rect 358452 369582 358504 369588
rect 358556 369374 358584 464850
rect 358820 461032 358872 461038
rect 358820 460974 358872 460980
rect 358636 459400 358688 459406
rect 358636 459342 358688 459348
rect 358648 373318 358676 459342
rect 358728 459332 358780 459338
rect 358728 459274 358780 459280
rect 358740 374202 358768 459274
rect 358728 374196 358780 374202
rect 358728 374138 358780 374144
rect 358636 373312 358688 373318
rect 358636 373254 358688 373260
rect 358544 369368 358596 369374
rect 358544 369310 358596 369316
rect 358832 356046 358860 460974
rect 358912 458312 358964 458318
rect 358912 458254 358964 458260
rect 358924 454753 358952 458254
rect 358910 454744 358966 454753
rect 358910 454679 358966 454688
rect 358820 356040 358872 356046
rect 358820 355982 358872 355988
rect 358924 349625 358952 454679
rect 359002 393816 359058 393825
rect 359002 393751 359058 393760
rect 359016 362234 359044 393751
rect 359094 392184 359150 392193
rect 359094 392119 359150 392128
rect 359108 362386 359136 392119
rect 359186 389328 359242 389337
rect 359186 389263 359242 389272
rect 359200 365022 359228 389263
rect 359476 374474 359504 475798
rect 359556 475788 359608 475794
rect 359556 475730 359608 475736
rect 359568 383654 359596 475730
rect 359648 459468 359700 459474
rect 359648 459410 359700 459416
rect 359660 385014 359688 459410
rect 359752 403646 359780 477226
rect 360752 471776 360804 471782
rect 360752 471718 360804 471724
rect 359924 464704 359976 464710
rect 359924 464646 359976 464652
rect 359832 463684 359884 463690
rect 359832 463626 359884 463632
rect 359844 405006 359872 463626
rect 359936 407794 359964 464646
rect 360568 464636 360620 464642
rect 360568 464578 360620 464584
rect 360580 409154 360608 464578
rect 360660 463616 360712 463622
rect 360660 463558 360712 463564
rect 360568 409148 360620 409154
rect 360568 409090 360620 409096
rect 359924 407788 359976 407794
rect 359924 407730 359976 407736
rect 359832 405000 359884 405006
rect 359832 404942 359884 404948
rect 359740 403640 359792 403646
rect 359740 403582 359792 403588
rect 359738 390824 359794 390833
rect 359738 390759 359794 390768
rect 359648 385008 359700 385014
rect 359648 384950 359700 384956
rect 359556 383648 359608 383654
rect 359556 383590 359608 383596
rect 359464 374468 359516 374474
rect 359464 374410 359516 374416
rect 359752 365022 359780 390759
rect 359830 388104 359886 388113
rect 359830 388039 359886 388048
rect 359188 365016 359240 365022
rect 359188 364958 359240 364964
rect 359740 365016 359792 365022
rect 359740 364958 359792 364964
rect 359200 364334 359228 364958
rect 359200 364306 359504 364334
rect 359108 362358 359320 362386
rect 359004 362228 359056 362234
rect 359004 362170 359056 362176
rect 359188 362228 359240 362234
rect 359188 362170 359240 362176
rect 359004 359508 359056 359514
rect 359004 359450 359056 359456
rect 358910 349616 358966 349625
rect 358910 349551 358966 349560
rect 358924 335354 358952 349551
rect 358832 335326 358952 335354
rect 358360 267368 358412 267374
rect 358360 267310 358412 267316
rect 358832 243817 358860 335326
rect 358910 288416 358966 288425
rect 358910 288351 358966 288360
rect 358924 287745 358952 288351
rect 358910 287736 358966 287745
rect 358910 287671 358966 287680
rect 358818 243808 358874 243817
rect 358818 243743 358874 243752
rect 358924 182753 358952 287671
rect 359016 286385 359044 359450
rect 359096 357400 359148 357406
rect 359096 357342 359148 357348
rect 359108 356726 359136 357342
rect 359096 356720 359148 356726
rect 359096 356662 359148 356668
rect 359002 286376 359058 286385
rect 359002 286311 359058 286320
rect 359016 277394 359044 286311
rect 359108 283121 359136 356662
rect 359200 289785 359228 362170
rect 359292 358057 359320 362358
rect 359476 359582 359504 364306
rect 359464 359576 359516 359582
rect 359464 359518 359516 359524
rect 359278 358048 359334 358057
rect 359278 357983 359334 357992
rect 359186 289776 359242 289785
rect 359186 289711 359242 289720
rect 359292 288425 359320 357983
rect 359278 288416 359334 288425
rect 359278 288351 359334 288360
rect 359476 284889 359504 359518
rect 359752 359514 359780 364958
rect 359844 363662 359872 388039
rect 360200 371340 360252 371346
rect 360200 371282 360252 371288
rect 359832 363656 359884 363662
rect 359832 363598 359884 363604
rect 359740 359508 359792 359514
rect 359740 359450 359792 359456
rect 359844 357406 359872 363598
rect 359832 357400 359884 357406
rect 359832 357342 359884 357348
rect 359554 289776 359610 289785
rect 359554 289711 359610 289720
rect 359462 284880 359518 284889
rect 359462 284815 359518 284824
rect 359094 283112 359150 283121
rect 359094 283047 359150 283056
rect 359370 283112 359426 283121
rect 359370 283047 359426 283056
rect 359016 277366 359228 277394
rect 359002 184920 359058 184929
rect 359002 184855 359058 184864
rect 358910 182744 358966 182753
rect 358910 182679 358966 182688
rect 358924 180794 358952 182679
rect 358832 180766 358952 180794
rect 358728 173188 358780 173194
rect 358728 173130 358780 173136
rect 358268 162104 358320 162110
rect 358268 162046 358320 162052
rect 358740 146266 358768 173130
rect 358728 146260 358780 146266
rect 358728 146202 358780 146208
rect 358740 145586 358768 146202
rect 358728 145580 358780 145586
rect 358728 145522 358780 145528
rect 358740 68338 358768 145522
rect 358832 78305 358860 180766
rect 358910 179480 358966 179489
rect 358910 179415 358966 179424
rect 358818 78296 358874 78305
rect 358818 78231 358874 78240
rect 358924 75449 358952 179415
rect 359016 79937 359044 184855
rect 359200 181393 359228 277366
rect 359278 243808 359334 243817
rect 359278 243743 359334 243752
rect 359186 181384 359242 181393
rect 359186 181319 359242 181328
rect 359094 178120 359150 178129
rect 359094 178055 359150 178064
rect 359002 79928 359058 79937
rect 359002 79863 359058 79872
rect 358910 75440 358966 75449
rect 358910 75375 358966 75384
rect 359108 74089 359136 178055
rect 359200 76945 359228 181319
rect 359292 139369 359320 243743
rect 359384 178129 359412 283047
rect 359476 179489 359504 284815
rect 359568 184929 359596 289711
rect 360212 267986 360240 371282
rect 360672 371006 360700 463558
rect 360764 374270 360792 471718
rect 360752 374264 360804 374270
rect 360752 374206 360804 374212
rect 360660 371000 360712 371006
rect 360660 370942 360712 370948
rect 360200 267980 360252 267986
rect 360200 267922 360252 267928
rect 359554 184920 359610 184929
rect 359554 184855 359610 184864
rect 359462 179480 359518 179489
rect 359462 179415 359518 179424
rect 359370 178120 359426 178129
rect 359370 178055 359426 178064
rect 359278 139360 359334 139369
rect 359278 139295 359334 139304
rect 359186 76936 359242 76945
rect 359186 76871 359242 76880
rect 359094 74080 359150 74089
rect 359094 74015 359150 74024
rect 358728 68332 358780 68338
rect 358728 68274 358780 68280
rect 358740 68202 358768 68274
rect 358728 68196 358780 68202
rect 358728 68138 358780 68144
rect 358176 59424 358228 59430
rect 358176 59366 358228 59372
rect 358084 59356 358136 59362
rect 358084 59298 358136 59304
rect 360856 58886 360884 478450
rect 362224 478236 362276 478242
rect 362224 478178 362276 478184
rect 361028 471640 361080 471646
rect 361028 471582 361080 471588
rect 360936 467288 360988 467294
rect 360936 467230 360988 467236
rect 360948 161906 360976 467230
rect 361040 268394 361068 471582
rect 361304 468988 361356 468994
rect 361304 468930 361356 468936
rect 361120 462052 361172 462058
rect 361120 461994 361172 462000
rect 361028 268388 361080 268394
rect 361028 268330 361080 268336
rect 361132 267714 361160 461994
rect 361212 459264 361264 459270
rect 361212 459206 361264 459212
rect 361120 267708 361172 267714
rect 361120 267650 361172 267656
rect 361224 267306 361252 459206
rect 361316 369714 361344 468930
rect 361396 466268 361448 466274
rect 361396 466210 361448 466216
rect 361304 369708 361356 369714
rect 361304 369650 361356 369656
rect 361408 367946 361436 466210
rect 362132 460148 362184 460154
rect 362132 460090 362184 460096
rect 361486 408640 361542 408649
rect 361486 408575 361542 408584
rect 361396 367940 361448 367946
rect 361396 367882 361448 367888
rect 361212 267300 361264 267306
rect 361212 267242 361264 267248
rect 360936 161900 360988 161906
rect 360936 161842 360988 161848
rect 360844 58880 360896 58886
rect 360844 58822 360896 58828
rect 361500 58750 361528 408575
rect 362144 371142 362172 460090
rect 362132 371136 362184 371142
rect 362132 371078 362184 371084
rect 362236 59022 362264 478178
rect 362328 164014 362356 478586
rect 365168 478576 365220 478582
rect 365168 478518 365220 478524
rect 363512 477216 363564 477222
rect 363512 477158 363564 477164
rect 362500 474496 362552 474502
rect 362500 474438 362552 474444
rect 362408 460624 362460 460630
rect 362408 460566 362460 460572
rect 362420 164286 362448 460566
rect 362512 267646 362540 474438
rect 362684 469124 362736 469130
rect 362684 469066 362736 469072
rect 362592 468852 362644 468858
rect 362592 468794 362644 468800
rect 362604 268530 362632 468794
rect 362696 370598 362724 469066
rect 363420 469056 363472 469062
rect 363420 468998 363472 469004
rect 362868 463344 362920 463350
rect 362868 463286 362920 463292
rect 362776 462256 362828 462262
rect 362776 462198 362828 462204
rect 362788 371890 362816 462198
rect 362880 374542 362908 463286
rect 363328 462120 363380 462126
rect 363328 462062 363380 462068
rect 362868 374536 362920 374542
rect 362868 374478 362920 374484
rect 362868 372632 362920 372638
rect 362868 372574 362920 372580
rect 362776 371884 362828 371890
rect 362776 371826 362828 371832
rect 362684 370592 362736 370598
rect 362684 370534 362736 370540
rect 362592 268524 362644 268530
rect 362592 268466 362644 268472
rect 362500 267640 362552 267646
rect 362500 267582 362552 267588
rect 362880 250578 362908 372574
rect 363340 369850 363368 462062
rect 363432 373386 363460 468998
rect 363420 373380 363472 373386
rect 363420 373322 363472 373328
rect 363524 370666 363552 477158
rect 364984 476876 365036 476882
rect 364984 476818 365036 476824
rect 363604 474156 363656 474162
rect 363604 474098 363656 474104
rect 363512 370660 363564 370666
rect 363512 370602 363564 370608
rect 363328 369844 363380 369850
rect 363328 369786 363380 369792
rect 362868 250572 362920 250578
rect 362868 250514 362920 250520
rect 362408 164280 362460 164286
rect 362408 164222 362460 164228
rect 362316 164008 362368 164014
rect 362316 163950 362368 163956
rect 362224 59016 362276 59022
rect 362224 58958 362276 58964
rect 361488 58744 361540 58750
rect 361488 58686 361540 58692
rect 357532 57928 357584 57934
rect 357532 57870 357584 57876
rect 356704 57860 356756 57866
rect 356704 57802 356756 57808
rect 363616 57798 363644 474098
rect 364892 472932 364944 472938
rect 364892 472874 364944 472880
rect 364064 470144 364116 470150
rect 364064 470086 364116 470092
rect 363696 465792 363748 465798
rect 363696 465734 363748 465740
rect 363604 57792 363656 57798
rect 363604 57734 363656 57740
rect 363708 57594 363736 465734
rect 363788 463004 363840 463010
rect 363788 462946 363840 462952
rect 363800 164422 363828 462946
rect 363972 460556 364024 460562
rect 363972 460498 364024 460504
rect 363880 459060 363932 459066
rect 363880 459002 363932 459008
rect 363788 164416 363840 164422
rect 363788 164358 363840 164364
rect 363892 162654 363920 459002
rect 363984 175234 364012 460498
rect 364076 267578 364104 470086
rect 364156 467424 364208 467430
rect 364156 467366 364208 467372
rect 364168 269346 364196 467366
rect 364800 463548 364852 463554
rect 364800 463490 364852 463496
rect 364246 372736 364302 372745
rect 364246 372671 364302 372680
rect 364156 269340 364208 269346
rect 364156 269282 364208 269288
rect 364064 267572 364116 267578
rect 364064 267514 364116 267520
rect 363972 175228 364024 175234
rect 363972 175170 364024 175176
rect 363880 162648 363932 162654
rect 363880 162590 363932 162596
rect 364260 57934 364288 372671
rect 364812 370870 364840 463490
rect 364904 371074 364932 472874
rect 364892 371068 364944 371074
rect 364892 371010 364944 371016
rect 364800 370864 364852 370870
rect 364800 370806 364852 370812
rect 364996 70378 365024 476818
rect 365076 458856 365128 458862
rect 365076 458798 365128 458804
rect 364984 70372 365036 70378
rect 364984 70314 365036 70320
rect 364248 57928 364300 57934
rect 364248 57870 364300 57876
rect 363696 57588 363748 57594
rect 363696 57530 363748 57536
rect 356612 57452 356664 57458
rect 356612 57394 356664 57400
rect 365088 57322 365116 458798
rect 365180 164082 365208 478518
rect 366456 478440 366508 478446
rect 366456 478382 366508 478388
rect 366364 478304 366416 478310
rect 366364 478246 366416 478252
rect 365628 477352 365680 477358
rect 365628 477294 365680 477300
rect 365444 475584 365496 475590
rect 365444 475526 365496 475532
rect 365260 468648 365312 468654
rect 365260 468590 365312 468596
rect 365168 164076 365220 164082
rect 365168 164018 365220 164024
rect 365272 162790 365300 468590
rect 365352 461712 365404 461718
rect 365352 461654 365404 461660
rect 365364 164121 365392 461654
rect 365456 267034 365484 475526
rect 365536 467628 365588 467634
rect 365536 467570 365588 467576
rect 365548 268462 365576 467570
rect 365640 370802 365668 477294
rect 366180 463412 366232 463418
rect 366180 463354 366232 463360
rect 366192 374134 366220 463354
rect 366272 458788 366324 458794
rect 366272 458730 366324 458736
rect 366180 374128 366232 374134
rect 366180 374070 366232 374076
rect 365628 370796 365680 370802
rect 365628 370738 365680 370744
rect 366284 369238 366312 458730
rect 366272 369232 366324 369238
rect 366272 369174 366324 369180
rect 365536 268456 365588 268462
rect 365536 268398 365588 268404
rect 365444 267028 365496 267034
rect 365444 266970 365496 266976
rect 365350 164112 365406 164121
rect 365350 164047 365406 164056
rect 365260 162784 365312 162790
rect 365260 162726 365312 162732
rect 366376 58954 366404 478246
rect 366364 58948 366416 58954
rect 366364 58890 366416 58896
rect 366468 58818 366496 478382
rect 373264 478168 373316 478174
rect 373264 478110 373316 478116
rect 372528 477420 372580 477426
rect 372528 477362 372580 477368
rect 368020 477012 368072 477018
rect 368020 476954 368072 476960
rect 366824 474428 366876 474434
rect 366824 474370 366876 474376
rect 366548 468580 366600 468586
rect 366548 468522 366600 468528
rect 366560 162314 366588 468522
rect 366640 465928 366692 465934
rect 366640 465870 366692 465876
rect 366652 163878 366680 465870
rect 366732 460352 366784 460358
rect 366732 460294 366784 460300
rect 366744 164354 366772 460294
rect 366836 268802 366864 474370
rect 366916 474292 366968 474298
rect 366916 474234 366968 474240
rect 366928 278730 366956 474234
rect 367836 474020 367888 474026
rect 367836 473962 367888 473968
rect 367652 464840 367704 464846
rect 367652 464782 367704 464788
rect 367560 463480 367612 463486
rect 367560 463422 367612 463428
rect 367008 463208 367060 463214
rect 367008 463150 367060 463156
rect 367020 370734 367048 463150
rect 367572 370938 367600 463422
rect 367560 370932 367612 370938
rect 367560 370874 367612 370880
rect 367008 370728 367060 370734
rect 367008 370670 367060 370676
rect 367664 369102 367692 464782
rect 367744 460964 367796 460970
rect 367744 460906 367796 460912
rect 367756 382226 367784 460906
rect 367744 382220 367796 382226
rect 367744 382162 367796 382168
rect 367744 371612 367796 371618
rect 367744 371554 367796 371560
rect 367652 369096 367704 369102
rect 367652 369038 367704 369044
rect 366916 278724 366968 278730
rect 366916 278666 366968 278672
rect 366824 268796 366876 268802
rect 366824 268738 366876 268744
rect 367756 265810 367784 371554
rect 367744 265804 367796 265810
rect 367744 265746 367796 265752
rect 366732 164348 366784 164354
rect 366732 164290 366784 164296
rect 366640 163872 366692 163878
rect 366640 163814 366692 163820
rect 366548 162308 366600 162314
rect 366548 162250 366600 162256
rect 366456 58812 366508 58818
rect 366456 58754 366508 58760
rect 367848 57662 367876 473962
rect 367928 469872 367980 469878
rect 367928 469814 367980 469820
rect 367940 57730 367968 469814
rect 368032 162450 368060 476954
rect 369768 475720 369820 475726
rect 369768 475662 369820 475668
rect 369216 475516 369268 475522
rect 369216 475458 369268 475464
rect 369124 474360 369176 474366
rect 369124 474302 369176 474308
rect 368388 468920 368440 468926
rect 368388 468862 368440 468868
rect 368204 468784 368256 468790
rect 368204 468726 368256 468732
rect 368112 460488 368164 460494
rect 368112 460430 368164 460436
rect 368124 163538 368152 460430
rect 368216 269142 368244 468726
rect 368296 460760 368348 460766
rect 368296 460702 368348 460708
rect 368308 280158 368336 460702
rect 368400 373590 368428 468862
rect 369032 466132 369084 466138
rect 369032 466074 369084 466080
rect 368388 373584 368440 373590
rect 368388 373526 368440 373532
rect 368388 371680 368440 371686
rect 368388 371622 368440 371628
rect 368296 280152 368348 280158
rect 368296 280094 368348 280100
rect 368204 269136 368256 269142
rect 368204 269078 368256 269084
rect 368400 251190 368428 371622
rect 369044 367810 369072 466074
rect 369032 367804 369084 367810
rect 369032 367746 369084 367752
rect 369136 268870 369164 474302
rect 369124 268864 369176 268870
rect 369124 268806 369176 268812
rect 368388 251184 368440 251190
rect 368388 251126 368440 251132
rect 369124 249824 369176 249830
rect 369124 249766 369176 249772
rect 369136 173874 369164 249766
rect 369124 173868 369176 173874
rect 369124 173810 369176 173816
rect 369136 173194 369164 173810
rect 369124 173188 369176 173194
rect 369124 173130 369176 173136
rect 368112 163532 368164 163538
rect 368112 163474 368164 163480
rect 369228 162518 369256 475458
rect 369676 472864 369728 472870
rect 369676 472806 369728 472812
rect 369492 471504 369544 471510
rect 369492 471446 369544 471452
rect 369308 465860 369360 465866
rect 369308 465802 369360 465808
rect 369320 163810 369348 465802
rect 369400 460420 369452 460426
rect 369400 460362 369452 460368
rect 369308 163804 369360 163810
rect 369308 163746 369360 163752
rect 369412 163742 369440 460362
rect 369504 267442 369532 471446
rect 369584 471436 369636 471442
rect 369584 471378 369636 471384
rect 369492 267436 369544 267442
rect 369492 267378 369544 267384
rect 369596 267102 369624 471378
rect 369688 369782 369716 472806
rect 369780 374338 369808 475662
rect 372436 475652 372488 475658
rect 372436 475594 372488 475600
rect 370596 474224 370648 474230
rect 370596 474166 370648 474172
rect 370504 467152 370556 467158
rect 370504 467094 370556 467100
rect 370412 463276 370464 463282
rect 370412 463218 370464 463224
rect 370320 461984 370372 461990
rect 370320 461926 370372 461932
rect 370228 459536 370280 459542
rect 370228 459478 370280 459484
rect 369768 374332 369820 374338
rect 369768 374274 369820 374280
rect 369768 373652 369820 373658
rect 369768 373594 369820 373600
rect 369676 369776 369728 369782
rect 369676 369718 369728 369724
rect 369584 267096 369636 267102
rect 369584 267038 369636 267044
rect 369780 264790 369808 373594
rect 369860 372020 369912 372026
rect 369860 371962 369912 371968
rect 369872 371482 369900 371962
rect 369860 371476 369912 371482
rect 369860 371418 369912 371424
rect 370240 369034 370268 459478
rect 370332 369442 370360 461926
rect 370424 373522 370452 463218
rect 370412 373516 370464 373522
rect 370412 373458 370464 373464
rect 370412 372020 370464 372026
rect 370412 371962 370464 371968
rect 370320 369436 370372 369442
rect 370320 369378 370372 369384
rect 370228 369028 370280 369034
rect 370228 368970 370280 368976
rect 370424 265878 370452 371962
rect 370412 265872 370464 265878
rect 370412 265814 370464 265820
rect 369768 264784 369820 264790
rect 369768 264726 369820 264732
rect 369400 163736 369452 163742
rect 369400 163678 369452 163684
rect 369216 162512 369268 162518
rect 369216 162454 369268 162460
rect 368020 162444 368072 162450
rect 368020 162386 368072 162392
rect 367928 57724 367980 57730
rect 367928 57666 367980 57672
rect 367836 57656 367888 57662
rect 367836 57598 367888 57604
rect 370516 57526 370544 467094
rect 370608 162246 370636 474166
rect 372252 472796 372304 472802
rect 372252 472738 372304 472744
rect 371976 471368 372028 471374
rect 371976 471310 372028 471316
rect 371792 470212 371844 470218
rect 371792 470154 371844 470160
rect 370688 470008 370740 470014
rect 370688 469950 370740 469956
rect 370700 162722 370728 469950
rect 370872 468716 370924 468722
rect 370872 468658 370924 468664
rect 370780 463140 370832 463146
rect 370780 463082 370832 463088
rect 370792 163985 370820 463082
rect 370884 267510 370912 468658
rect 371240 466200 371292 466206
rect 371240 466142 371292 466148
rect 371056 465996 371108 466002
rect 371056 465938 371108 465944
rect 370964 460692 371016 460698
rect 370964 460634 371016 460640
rect 370976 269210 371004 460634
rect 371068 372162 371096 465938
rect 371146 372736 371202 372745
rect 371146 372671 371202 372680
rect 371056 372156 371108 372162
rect 371056 372098 371108 372104
rect 371056 369028 371108 369034
rect 371056 368970 371108 368976
rect 370964 269204 371016 269210
rect 370964 269146 371016 269152
rect 370872 267504 370924 267510
rect 370872 267446 370924 267452
rect 370964 265804 371016 265810
rect 370964 265746 371016 265752
rect 370778 163976 370834 163985
rect 370778 163911 370834 163920
rect 370688 162716 370740 162722
rect 370688 162658 370740 162664
rect 370596 162240 370648 162246
rect 370596 162182 370648 162188
rect 370976 147626 371004 265746
rect 371068 250714 371096 368970
rect 371160 250782 371188 372671
rect 371252 372638 371280 466142
rect 371804 373726 371832 470154
rect 371884 465724 371936 465730
rect 371884 465666 371936 465672
rect 371792 373720 371844 373726
rect 371792 373662 371844 373668
rect 371240 372632 371292 372638
rect 371240 372574 371292 372580
rect 371252 372337 371280 372574
rect 371238 372328 371294 372337
rect 371238 372263 371294 372272
rect 371240 371748 371292 371754
rect 371240 371690 371292 371696
rect 371608 371748 371660 371754
rect 371608 371690 371660 371696
rect 371252 371550 371280 371690
rect 371240 371544 371292 371550
rect 371240 371486 371292 371492
rect 371620 266150 371648 371690
rect 371792 369096 371844 369102
rect 371792 369038 371844 369044
rect 371700 354000 371752 354006
rect 371700 353942 371752 353948
rect 371608 266144 371660 266150
rect 371608 266086 371660 266092
rect 371712 265674 371740 353942
rect 371700 265668 371752 265674
rect 371700 265610 371752 265616
rect 371804 265305 371832 369038
rect 371790 265296 371846 265305
rect 371790 265231 371846 265240
rect 371792 251184 371844 251190
rect 371792 251126 371844 251132
rect 371148 250776 371200 250782
rect 371148 250718 371200 250724
rect 371056 250708 371108 250714
rect 371056 250650 371108 250656
rect 371804 250646 371832 251126
rect 371792 250640 371844 250646
rect 371792 250582 371844 250588
rect 371804 148374 371832 250582
rect 371792 148368 371844 148374
rect 371792 148310 371844 148316
rect 370964 147620 371016 147626
rect 370964 147562 371016 147568
rect 370504 57520 370556 57526
rect 370504 57462 370556 57468
rect 371896 57458 371924 465666
rect 371988 162586 372016 471310
rect 372068 463072 372120 463078
rect 372068 463014 372120 463020
rect 372080 163674 372108 463014
rect 372160 458924 372212 458930
rect 372160 458866 372212 458872
rect 372172 173806 372200 458866
rect 372264 267238 372292 472738
rect 372344 461916 372396 461922
rect 372344 461858 372396 461864
rect 372356 268598 372384 461858
rect 372448 374406 372476 475594
rect 372436 374400 372488 374406
rect 372436 374342 372488 374348
rect 372436 369572 372488 369578
rect 372436 369514 372488 369520
rect 372344 268592 372396 268598
rect 372344 268534 372396 268540
rect 372252 267232 372304 267238
rect 372252 267174 372304 267180
rect 372344 266144 372396 266150
rect 372344 266086 372396 266092
rect 372252 251116 372304 251122
rect 372252 251058 372304 251064
rect 372160 173800 372212 173806
rect 372160 173742 372212 173748
rect 372068 163668 372120 163674
rect 372068 163610 372120 163616
rect 371976 162580 372028 162586
rect 371976 162522 372028 162528
rect 372264 161430 372292 251058
rect 372252 161424 372304 161430
rect 372252 161366 372304 161372
rect 372160 148912 372212 148918
rect 372160 148854 372212 148860
rect 371884 57452 371936 57458
rect 371884 57394 371936 57400
rect 365076 57316 365128 57322
rect 365076 57258 365128 57264
rect 307758 55176 307814 55185
rect 307758 55111 307814 55120
rect 270500 55014 270552 55020
rect 277398 55040 277454 55049
rect 267740 55004 267792 55010
rect 277398 54975 277454 54984
rect 267740 54946 267792 54952
rect 253940 54936 253992 54942
rect 253940 54878 253992 54884
rect 249798 54839 249854 54848
rect 251364 54868 251416 54874
rect 251364 54810 251416 54816
rect 247040 54800 247092 54806
rect 247040 54742 247092 54748
rect 244372 54596 244424 54602
rect 244372 54538 244424 54544
rect 240140 54528 240192 54534
rect 240140 54470 240192 54476
rect 372172 54466 372200 148854
rect 372264 56506 372292 161366
rect 372356 148986 372384 266086
rect 372448 251122 372476 369514
rect 372540 368490 372568 477362
rect 373172 466064 373224 466070
rect 373172 466006 373224 466012
rect 373184 372570 373212 466006
rect 373172 372564 373224 372570
rect 373172 372506 373224 372512
rect 372896 372360 372948 372366
rect 372896 372302 372948 372308
rect 372908 371414 372936 372302
rect 372896 371408 372948 371414
rect 372896 371350 372948 371356
rect 373080 370524 373132 370530
rect 373080 370466 373132 370472
rect 372528 368484 372580 368490
rect 372528 368426 372580 368432
rect 373092 267986 373120 370466
rect 373172 367804 373224 367810
rect 373172 367746 373224 367752
rect 373184 268122 373212 367746
rect 373172 268116 373224 268122
rect 373172 268058 373224 268064
rect 373080 267980 373132 267986
rect 373080 267922 373132 267928
rect 372528 265872 372580 265878
rect 372528 265814 372580 265820
rect 372436 251116 372488 251122
rect 372436 251058 372488 251064
rect 372436 250572 372488 250578
rect 372436 250514 372488 250520
rect 372344 148980 372396 148986
rect 372344 148922 372396 148928
rect 372252 56500 372304 56506
rect 372252 56442 372304 56448
rect 372356 55894 372384 148922
rect 372448 144129 372476 250514
rect 372540 148510 372568 265814
rect 373172 265668 373224 265674
rect 373172 265610 373224 265616
rect 372528 148504 372580 148510
rect 372528 148446 372580 148452
rect 373184 144906 373212 265610
rect 373172 144900 373224 144906
rect 373172 144842 373224 144848
rect 372434 144120 372490 144129
rect 372434 144055 372490 144064
rect 373276 59090 373304 478110
rect 374184 477148 374236 477154
rect 374184 477090 374236 477096
rect 373908 475924 373960 475930
rect 373908 475866 373960 475872
rect 373724 474564 373776 474570
rect 373724 474506 373776 474512
rect 373448 467356 373500 467362
rect 373448 467298 373500 467304
rect 373356 460284 373408 460290
rect 373356 460226 373408 460232
rect 373368 163606 373396 460226
rect 373460 267170 373488 467298
rect 373540 461780 373592 461786
rect 373540 461722 373592 461728
rect 373448 267164 373500 267170
rect 373448 267106 373500 267112
rect 373552 266937 373580 461722
rect 373632 459128 373684 459134
rect 373632 459070 373684 459076
rect 373644 269278 373672 459070
rect 373736 373454 373764 474506
rect 373816 471980 373868 471986
rect 373816 471922 373868 471928
rect 373724 373448 373776 373454
rect 373724 373390 373776 373396
rect 373724 371408 373776 371414
rect 373724 371350 373776 371356
rect 373632 269272 373684 269278
rect 373632 269214 373684 269220
rect 373736 267734 373764 371350
rect 373828 369510 373856 471922
rect 373816 369504 373868 369510
rect 373816 369446 373868 369452
rect 373644 267706 373764 267734
rect 373538 266928 373594 266937
rect 373538 266863 373594 266872
rect 373644 266014 373672 267706
rect 373632 266008 373684 266014
rect 373632 265950 373684 265956
rect 373448 251184 373500 251190
rect 373448 251126 373500 251132
rect 373356 163600 373408 163606
rect 373356 163542 373408 163548
rect 373460 160818 373488 251126
rect 373540 250708 373592 250714
rect 373540 250650 373592 250656
rect 373448 160812 373500 160818
rect 373448 160754 373500 160760
rect 373552 160750 373580 250650
rect 373540 160744 373592 160750
rect 373540 160686 373592 160692
rect 373644 148918 373672 265950
rect 373724 265736 373776 265742
rect 373724 265678 373776 265684
rect 373632 148912 373684 148918
rect 373632 148854 373684 148860
rect 373736 144770 373764 265678
rect 373828 251190 373856 369446
rect 373920 369306 373948 475866
rect 374000 473136 374052 473142
rect 374000 473078 374052 473084
rect 374012 378826 374040 473078
rect 374000 378820 374052 378826
rect 374000 378762 374052 378768
rect 373908 369300 373960 369306
rect 373908 369242 373960 369248
rect 373906 269376 373962 269385
rect 373906 269311 373962 269320
rect 373816 251184 373868 251190
rect 373816 251126 373868 251132
rect 373920 146305 373948 269311
rect 374196 267481 374224 477090
rect 376392 477080 376444 477086
rect 376392 477022 376444 477028
rect 374736 476944 374788 476950
rect 374736 476886 374788 476892
rect 374644 475380 374696 475386
rect 374644 475322 374696 475328
rect 374460 460080 374512 460086
rect 374460 460022 374512 460028
rect 374368 378820 374420 378826
rect 374368 378762 374420 378768
rect 374380 369578 374408 378762
rect 374368 369572 374420 369578
rect 374368 369514 374420 369520
rect 374380 368422 374408 369514
rect 374472 369102 374500 460022
rect 374552 370796 374604 370802
rect 374552 370738 374604 370744
rect 374460 369096 374512 369102
rect 374460 369038 374512 369044
rect 374460 368484 374512 368490
rect 374460 368426 374512 368432
rect 374368 368416 374420 368422
rect 374368 368358 374420 368364
rect 374472 269074 374500 368426
rect 374460 269068 374512 269074
rect 374460 269010 374512 269016
rect 374564 268938 374592 370738
rect 374552 268932 374604 268938
rect 374552 268874 374604 268880
rect 374276 268116 374328 268122
rect 374276 268058 374328 268064
rect 374182 267472 374238 267481
rect 374182 267407 374238 267416
rect 374288 149054 374316 268058
rect 374366 266384 374422 266393
rect 374366 266319 374422 266328
rect 374276 149048 374328 149054
rect 374276 148990 374328 148996
rect 374288 148238 374316 148990
rect 374276 148232 374328 148238
rect 374276 148174 374328 148180
rect 373906 146296 373962 146305
rect 373906 146231 373962 146240
rect 374380 145994 374408 266319
rect 374552 264988 374604 264994
rect 374552 264930 374604 264936
rect 374460 250776 374512 250782
rect 374460 250718 374512 250724
rect 374472 165578 374500 250718
rect 374460 165572 374512 165578
rect 374460 165514 374512 165520
rect 374564 164150 374592 264930
rect 374552 164144 374604 164150
rect 374552 164086 374604 164092
rect 374552 146192 374604 146198
rect 374552 146134 374604 146140
rect 374460 146124 374512 146130
rect 374460 146066 374512 146072
rect 374368 145988 374420 145994
rect 374368 145930 374420 145936
rect 373724 144764 373776 144770
rect 373724 144706 373776 144712
rect 373264 59084 373316 59090
rect 373264 59026 373316 59032
rect 374472 58614 374500 146066
rect 374564 59294 374592 146134
rect 374656 69018 374684 475322
rect 374748 162489 374776 476886
rect 376208 475448 376260 475454
rect 376208 475390 376260 475396
rect 375472 473952 375524 473958
rect 375472 473894 375524 473900
rect 375196 471912 375248 471918
rect 375196 471854 375248 471860
rect 374828 469940 374880 469946
rect 374828 469882 374880 469888
rect 374734 162480 374790 162489
rect 374734 162415 374790 162424
rect 374840 162382 374868 469882
rect 375104 461848 375156 461854
rect 375104 461790 375156 461796
rect 375012 461644 375064 461650
rect 375012 461586 375064 461592
rect 374920 370660 374972 370666
rect 374920 370602 374972 370608
rect 374932 367606 374960 370602
rect 374920 367600 374972 367606
rect 374920 367542 374972 367548
rect 374920 269068 374972 269074
rect 374920 269010 374972 269016
rect 374932 267850 374960 269010
rect 374920 267844 374972 267850
rect 374920 267786 374972 267792
rect 374932 163062 374960 267786
rect 375024 266898 375052 461586
rect 375116 268666 375144 461790
rect 375208 372230 375236 471854
rect 375288 467492 375340 467498
rect 375288 467434 375340 467440
rect 375300 373862 375328 467434
rect 375380 382220 375432 382226
rect 375380 382162 375432 382168
rect 375288 373856 375340 373862
rect 375288 373798 375340 373804
rect 375196 372224 375248 372230
rect 375196 372166 375248 372172
rect 375196 370796 375248 370802
rect 375196 370738 375248 370744
rect 375208 370530 375236 370738
rect 375288 370660 375340 370666
rect 375288 370602 375340 370608
rect 375196 370524 375248 370530
rect 375196 370466 375248 370472
rect 375300 370394 375328 370602
rect 375288 370388 375340 370394
rect 375288 370330 375340 370336
rect 375196 369300 375248 369306
rect 375196 369242 375248 369248
rect 375208 367690 375236 369242
rect 375288 368484 375340 368490
rect 375288 368426 375340 368432
rect 375300 367878 375328 368426
rect 375288 367872 375340 367878
rect 375288 367814 375340 367820
rect 375208 367662 375328 367690
rect 375196 367600 375248 367606
rect 375196 367542 375248 367548
rect 375104 268660 375156 268666
rect 375104 268602 375156 268608
rect 375208 267209 375236 367542
rect 375194 267200 375250 267209
rect 375194 267135 375250 267144
rect 375012 266892 375064 266898
rect 375012 266834 375064 266840
rect 375208 266393 375236 267135
rect 375194 266384 375250 266393
rect 375194 266319 375250 266328
rect 375300 265402 375328 367662
rect 375392 355366 375420 382162
rect 375484 373658 375512 473894
rect 376116 471300 376168 471306
rect 376116 471242 376168 471248
rect 375932 467560 375984 467566
rect 375932 467502 375984 467508
rect 375748 462188 375800 462194
rect 375748 462130 375800 462136
rect 375472 373652 375524 373658
rect 375472 373594 375524 373600
rect 375760 368490 375788 462130
rect 375944 373794 375972 467502
rect 375932 373788 375984 373794
rect 375932 373730 375984 373736
rect 375840 369232 375892 369238
rect 375840 369174 375892 369180
rect 375748 368484 375800 368490
rect 375748 368426 375800 368432
rect 375380 355360 375432 355366
rect 375380 355302 375432 355308
rect 375392 355162 375420 355302
rect 375380 355156 375432 355162
rect 375380 355098 375432 355104
rect 375656 267980 375708 267986
rect 375656 267922 375708 267928
rect 375288 265396 375340 265402
rect 375288 265338 375340 265344
rect 375104 265328 375156 265334
rect 375104 265270 375156 265276
rect 374920 163056 374972 163062
rect 374920 162998 374972 163004
rect 374828 162376 374880 162382
rect 374828 162318 374880 162324
rect 374828 160744 374880 160750
rect 374828 160686 374880 160692
rect 374736 148504 374788 148510
rect 374736 148446 374788 148452
rect 374644 69012 374696 69018
rect 374644 68954 374696 68960
rect 374552 59288 374604 59294
rect 374552 59230 374604 59236
rect 374460 58608 374512 58614
rect 374460 58550 374512 58556
rect 372344 55888 372396 55894
rect 372344 55830 372396 55836
rect 214564 54460 214616 54466
rect 214564 54402 214616 54408
rect 237380 54460 237432 54466
rect 237380 54402 237432 54408
rect 372160 54460 372212 54466
rect 372160 54402 372212 54408
rect 374748 54398 374776 148446
rect 374840 55010 374868 160686
rect 374932 56370 374960 162998
rect 375012 148232 375064 148238
rect 375012 148174 375064 148180
rect 374920 56364 374972 56370
rect 374920 56306 374972 56312
rect 375024 55146 375052 148174
rect 375116 146130 375144 265270
rect 375196 265260 375248 265266
rect 375196 265202 375248 265208
rect 375104 146124 375156 146130
rect 375104 146066 375156 146072
rect 375116 145858 375144 146066
rect 375104 145852 375156 145858
rect 375104 145794 375156 145800
rect 375208 145738 375236 265202
rect 375300 264994 375328 265338
rect 375378 265160 375434 265169
rect 375378 265095 375434 265104
rect 375288 264988 375340 264994
rect 375288 264930 375340 264936
rect 375392 160002 375420 265095
rect 375470 265024 375526 265033
rect 375470 264959 375526 264968
rect 375380 159996 375432 160002
rect 375380 159938 375432 159944
rect 375392 158794 375420 159938
rect 375484 158817 375512 264959
rect 375564 165572 375616 165578
rect 375564 165514 375616 165520
rect 375576 164490 375604 165514
rect 375564 164484 375616 164490
rect 375564 164426 375616 164432
rect 375116 145710 375236 145738
rect 375300 158766 375420 158794
rect 375470 158808 375526 158817
rect 375116 144838 375144 145710
rect 375196 145580 375248 145586
rect 375196 145522 375248 145528
rect 375208 144906 375236 145522
rect 375196 144900 375248 144906
rect 375196 144842 375248 144848
rect 375104 144832 375156 144838
rect 375104 144774 375156 144780
rect 375208 142154 375236 144842
rect 375116 142126 375236 142154
rect 375012 55140 375064 55146
rect 375012 55082 375064 55088
rect 374828 55004 374880 55010
rect 374828 54946 374880 54952
rect 375116 54670 375144 142126
rect 375300 59158 375328 158766
rect 375470 158743 375526 158752
rect 375288 59152 375340 59158
rect 375288 59094 375340 59100
rect 375576 55078 375604 164426
rect 375668 146198 375696 267922
rect 375852 265169 375880 369174
rect 375932 369096 375984 369102
rect 375932 369038 375984 369044
rect 375838 265160 375894 265169
rect 375748 265124 375800 265130
rect 375838 265095 375894 265104
rect 375748 265066 375800 265072
rect 375656 146192 375708 146198
rect 375656 146134 375708 146140
rect 375668 145722 375696 146134
rect 375760 145926 375788 265066
rect 375944 265033 375972 369038
rect 376024 355156 376076 355162
rect 376024 355098 376076 355104
rect 376036 278322 376064 355098
rect 376024 278316 376076 278322
rect 376024 278258 376076 278264
rect 375930 265024 375986 265033
rect 375930 264959 375986 264968
rect 375840 263152 375892 263158
rect 375840 263094 375892 263100
rect 375852 164218 375880 263094
rect 376036 249830 376064 278258
rect 376024 249824 376076 249830
rect 376024 249766 376076 249772
rect 375840 164212 375892 164218
rect 375840 164154 375892 164160
rect 376024 147620 376076 147626
rect 376024 147562 376076 147568
rect 375748 145920 375800 145926
rect 375748 145862 375800 145868
rect 375656 145716 375708 145722
rect 375656 145658 375708 145664
rect 375760 145518 375788 145862
rect 375930 145616 375986 145625
rect 375930 145551 375986 145560
rect 375748 145512 375800 145518
rect 375748 145454 375800 145460
rect 375944 59498 375972 145551
rect 375932 59492 375984 59498
rect 375932 59434 375984 59440
rect 376036 56574 376064 147562
rect 376128 57390 376156 471242
rect 376220 162625 376248 475390
rect 376300 474088 376352 474094
rect 376300 474030 376352 474036
rect 376206 162616 376262 162625
rect 376206 162551 376262 162560
rect 376312 161974 376340 474030
rect 376404 268734 376432 477022
rect 377772 473000 377824 473006
rect 377772 472942 377824 472948
rect 376484 470076 376536 470082
rect 376484 470018 376536 470024
rect 376392 268728 376444 268734
rect 376392 268670 376444 268676
rect 376496 266830 376524 470018
rect 376576 467696 376628 467702
rect 376576 467638 376628 467644
rect 376588 371482 376616 467638
rect 377496 464432 377548 464438
rect 377496 464374 377548 464380
rect 377404 464364 377456 464370
rect 377404 464306 377456 464312
rect 377128 460896 377180 460902
rect 377128 460838 377180 460844
rect 377036 409148 377088 409154
rect 377036 409090 377088 409096
rect 377048 408785 377076 409090
rect 377034 408776 377090 408785
rect 377034 408711 377090 408720
rect 376942 407824 376998 407833
rect 376760 407788 376812 407794
rect 376942 407759 376944 407768
rect 376760 407730 376812 407736
rect 376996 407759 376998 407768
rect 376944 407730 376996 407736
rect 376666 383344 376722 383353
rect 376666 383279 376722 383288
rect 376680 382226 376708 383279
rect 376668 382220 376720 382226
rect 376668 382162 376720 382168
rect 376666 373280 376722 373289
rect 376666 373215 376722 373224
rect 376576 371476 376628 371482
rect 376576 371418 376628 371424
rect 376576 368484 376628 368490
rect 376576 368426 376628 368432
rect 376484 266824 376536 266830
rect 376484 266766 376536 266772
rect 376588 266098 376616 368426
rect 376404 266070 376616 266098
rect 376404 263566 376432 266070
rect 376576 265940 376628 265946
rect 376576 265882 376628 265888
rect 376588 265742 376616 265882
rect 376680 265742 376708 373215
rect 376772 302841 376800 407730
rect 376944 385008 376996 385014
rect 376942 384976 376944 384985
rect 376996 384976 376998 384985
rect 376942 384911 376998 384920
rect 376944 383648 376996 383654
rect 376944 383590 376996 383596
rect 376956 383081 376984 383590
rect 376942 383072 376998 383081
rect 376942 383007 376998 383016
rect 377140 373994 377168 460838
rect 377416 412634 377444 464306
rect 377508 422294 377536 464374
rect 377508 422266 377628 422294
rect 377416 412606 377536 412634
rect 377508 410961 377536 412606
rect 377600 411913 377628 422266
rect 377586 411904 377642 411913
rect 377586 411839 377642 411848
rect 377494 410952 377550 410961
rect 377494 410887 377550 410896
rect 377310 408776 377366 408785
rect 377310 408711 377366 408720
rect 377220 406428 377272 406434
rect 377220 406370 377272 406376
rect 377232 406065 377260 406370
rect 377218 406056 377274 406065
rect 377218 405991 377274 406000
rect 377324 405906 377352 408711
rect 377048 373966 377168 373994
rect 377232 405878 377352 405906
rect 377048 371414 377076 373966
rect 377036 371408 377088 371414
rect 377036 371350 377088 371356
rect 376944 369368 376996 369374
rect 376944 369310 376996 369316
rect 376956 368529 376984 369310
rect 376942 368520 376998 368529
rect 376942 368455 376998 368464
rect 376850 307728 376906 307737
rect 376850 307663 376906 307672
rect 376864 306921 376892 307663
rect 376850 306912 376906 306921
rect 376850 306847 376906 306856
rect 376758 302832 376814 302841
rect 376758 302767 376814 302776
rect 376758 301064 376814 301073
rect 376758 300999 376814 301008
rect 376576 265736 376628 265742
rect 376576 265678 376628 265684
rect 376668 265736 376720 265742
rect 376668 265678 376720 265684
rect 376482 265296 376538 265305
rect 376482 265231 376538 265240
rect 376392 263560 376444 263566
rect 376392 263502 376444 263508
rect 376404 263158 376432 263502
rect 376392 263152 376444 263158
rect 376392 263094 376444 263100
rect 376496 171134 376524 265231
rect 376772 196081 376800 300999
rect 376864 202881 376892 306847
rect 376942 305008 376998 305017
rect 376942 304943 376998 304952
rect 376850 202872 376906 202881
rect 376850 202807 376906 202816
rect 376956 200977 376984 304943
rect 377232 303793 377260 405878
rect 377312 405000 377364 405006
rect 377310 404968 377312 404977
rect 377364 404968 377366 404977
rect 377310 404903 377366 404912
rect 377218 303784 377274 303793
rect 377218 303719 377274 303728
rect 377036 280152 377088 280158
rect 377036 280094 377088 280100
rect 377048 279993 377076 280094
rect 377034 279984 377090 279993
rect 377034 279919 377090 279928
rect 377036 278724 377088 278730
rect 377036 278666 377088 278672
rect 377048 278089 377076 278666
rect 377034 278080 377090 278089
rect 377034 278015 377090 278024
rect 377036 265192 377088 265198
rect 377036 265134 377088 265140
rect 376942 200968 376998 200977
rect 376942 200903 376998 200912
rect 376758 196072 376814 196081
rect 376758 196007 376814 196016
rect 376852 175228 376904 175234
rect 376852 175170 376904 175176
rect 376864 175001 376892 175170
rect 376850 174992 376906 175001
rect 376850 174927 376906 174936
rect 376852 173868 376904 173874
rect 376852 173810 376904 173816
rect 376760 173800 376812 173806
rect 376760 173742 376812 173748
rect 376772 173097 376800 173742
rect 376864 173369 376892 173810
rect 376850 173360 376906 173369
rect 376850 173295 376906 173304
rect 376758 173088 376814 173097
rect 376758 173023 376814 173032
rect 376496 171106 376708 171134
rect 376392 164212 376444 164218
rect 376392 164154 376444 164160
rect 376404 162926 376432 164154
rect 376392 162920 376444 162926
rect 376392 162862 376444 162868
rect 376300 161968 376352 161974
rect 376300 161910 376352 161916
rect 376300 160812 376352 160818
rect 376300 160754 376352 160760
rect 376208 144764 376260 144770
rect 376208 144706 376260 144712
rect 376116 57384 376168 57390
rect 376116 57326 376168 57332
rect 376024 56568 376076 56574
rect 376024 56510 376076 56516
rect 375564 55072 375616 55078
rect 375564 55014 375616 55020
rect 375104 54664 375156 54670
rect 375104 54606 375156 54612
rect 376220 54534 376248 144706
rect 376312 54942 376340 160754
rect 376404 55214 376432 162862
rect 376680 160070 376708 171106
rect 376668 160064 376720 160070
rect 376668 160006 376720 160012
rect 376576 148436 376628 148442
rect 376576 148378 376628 148384
rect 376588 147626 376616 148378
rect 376576 147620 376628 147626
rect 376576 147562 376628 147568
rect 376482 146296 376538 146305
rect 376482 146231 376538 146240
rect 376496 145625 376524 146231
rect 376576 145648 376628 145654
rect 376482 145616 376538 145625
rect 376576 145590 376628 145596
rect 376482 145551 376538 145560
rect 376484 145512 376536 145518
rect 376484 145454 376536 145460
rect 376496 142154 376524 145454
rect 376588 144770 376616 145590
rect 376576 144764 376628 144770
rect 376576 144706 376628 144712
rect 376496 142126 376616 142154
rect 376392 55208 376444 55214
rect 376392 55150 376444 55156
rect 376300 54936 376352 54942
rect 376300 54878 376352 54884
rect 376588 54602 376616 142126
rect 376680 59226 376708 160006
rect 376956 95985 376984 200903
rect 377048 145314 377076 265134
rect 377128 263628 377180 263634
rect 377128 263570 377180 263576
rect 377140 163198 377168 263570
rect 377232 198801 377260 303719
rect 377324 299985 377352 404903
rect 377404 372564 377456 372570
rect 377404 372506 377456 372512
rect 377416 371929 377444 372506
rect 377402 371920 377458 371929
rect 377402 371855 377458 371864
rect 377508 305969 377536 410887
rect 377600 307737 377628 411839
rect 377678 406056 377734 406065
rect 377678 405991 377734 406000
rect 377586 307728 377642 307737
rect 377586 307663 377642 307672
rect 377494 305960 377550 305969
rect 377494 305895 377550 305904
rect 377508 305017 377536 305895
rect 377494 305008 377550 305017
rect 377494 304943 377550 304952
rect 377586 302832 377642 302841
rect 377586 302767 377642 302776
rect 377310 299976 377366 299985
rect 377310 299911 377366 299920
rect 377218 198792 377274 198801
rect 377218 198727 377274 198736
rect 377324 194993 377352 299911
rect 377402 278352 377458 278361
rect 377402 278287 377404 278296
rect 377456 278287 377458 278296
rect 377404 278258 377456 278264
rect 377494 202872 377550 202881
rect 377494 202807 377550 202816
rect 377508 201929 377536 202807
rect 377494 201920 377550 201929
rect 377494 201855 377550 201864
rect 377310 194984 377366 194993
rect 377310 194919 377366 194928
rect 377128 163192 377180 163198
rect 377128 163134 377180 163140
rect 377140 156670 377168 163134
rect 377128 156664 377180 156670
rect 377128 156606 377180 156612
rect 377220 146192 377272 146198
rect 377220 146134 377272 146140
rect 377036 145308 377088 145314
rect 377036 145250 377088 145256
rect 376942 95976 376998 95985
rect 376942 95911 376998 95920
rect 376944 70372 376996 70378
rect 376944 70314 376996 70320
rect 376956 70009 376984 70314
rect 376942 70000 376998 70009
rect 376942 69935 376998 69944
rect 376942 68368 376998 68377
rect 376942 68303 376944 68312
rect 376996 68303 376998 68312
rect 376944 68274 376996 68280
rect 376668 59220 376720 59226
rect 376668 59162 376720 59168
rect 377048 54806 377076 145250
rect 377036 54800 377088 54806
rect 377036 54742 377088 54748
rect 377232 54738 377260 146134
rect 377324 90001 377352 194919
rect 377508 96937 377536 201855
rect 377600 197849 377628 302767
rect 377692 301073 377720 405991
rect 377784 405686 377812 472942
rect 378152 468518 378180 520118
rect 383672 518430 383700 520118
rect 387904 518498 387932 520118
rect 387892 518492 387944 518498
rect 387892 518434 387944 518440
rect 383660 518424 383712 518430
rect 383660 518366 383712 518372
rect 391952 485081 391980 520118
rect 396920 519110 396948 520118
rect 396908 519104 396960 519110
rect 396908 519046 396960 519052
rect 401612 518634 401640 520118
rect 401600 518628 401652 518634
rect 401600 518570 401652 518576
rect 406028 518566 406056 520118
rect 406016 518560 406068 518566
rect 406016 518502 406068 518508
rect 410536 518022 410564 520118
rect 414952 519042 414980 520118
rect 414940 519036 414992 519042
rect 414940 518978 414992 518984
rect 419552 518090 419580 520118
rect 423968 518702 423996 520118
rect 423956 518696 424008 518702
rect 423956 518638 424008 518644
rect 419540 518084 419592 518090
rect 419540 518026 419592 518032
rect 410524 518016 410576 518022
rect 410524 517958 410576 517964
rect 427832 514690 427860 520231
rect 428384 514758 428412 558175
rect 429212 518974 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 430948 641028 431000 641034
rect 430948 640970 431000 640976
rect 429292 638240 429344 638246
rect 429292 638182 429344 638188
rect 429304 530301 429332 638182
rect 430580 634976 430632 634982
rect 430580 634918 430632 634924
rect 429844 631236 429896 631242
rect 429844 631178 429896 631184
rect 429856 621722 429884 631178
rect 429844 621716 429896 621722
rect 429844 621658 429896 621664
rect 430592 607209 430620 634918
rect 430856 634908 430908 634914
rect 430856 634850 430908 634856
rect 430764 633616 430816 633622
rect 430764 633558 430816 633564
rect 430672 631304 430724 631310
rect 430672 631246 430724 631252
rect 430684 612513 430712 631246
rect 430776 616865 430804 633558
rect 430868 622033 430896 634850
rect 430960 626521 430988 640970
rect 457444 634840 457496 634846
rect 457444 634782 457496 634788
rect 432604 632800 432656 632806
rect 432604 632742 432656 632748
rect 430946 626512 431002 626521
rect 430946 626447 431002 626456
rect 430854 622024 430910 622033
rect 430854 621959 430910 621968
rect 432616 619614 432644 632742
rect 435364 631168 435416 631174
rect 435364 631110 435416 631116
rect 432696 631100 432748 631106
rect 432696 631042 432748 631048
rect 432708 621790 432736 631042
rect 435376 621858 435404 631110
rect 435364 621852 435416 621858
rect 435364 621794 435416 621800
rect 432696 621784 432748 621790
rect 432696 621726 432748 621732
rect 432604 619608 432656 619614
rect 432604 619550 432656 619556
rect 456800 619608 456852 619614
rect 456800 619550 456852 619556
rect 456812 619041 456840 619550
rect 456798 619032 456854 619041
rect 456798 618967 456854 618976
rect 430762 616856 430818 616865
rect 430762 616791 430818 616800
rect 430670 612504 430726 612513
rect 430670 612439 430726 612448
rect 456800 611312 456852 611318
rect 456800 611254 456852 611260
rect 456812 610881 456840 611254
rect 456798 610872 456854 610881
rect 456798 610807 456854 610816
rect 430578 607200 430634 607209
rect 430578 607135 430634 607144
rect 457456 602721 457484 634782
rect 494072 634098 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 494060 634092 494112 634098
rect 494060 634034 494112 634040
rect 489920 633548 489972 633554
rect 489920 633490 489972 633496
rect 466736 630964 466788 630970
rect 466736 630906 466788 630912
rect 466748 619970 466776 630906
rect 474832 621852 474884 621858
rect 474832 621794 474884 621800
rect 466748 619942 467130 619970
rect 474844 619956 474872 621794
rect 482560 621036 482612 621042
rect 482560 620978 482612 620984
rect 482572 619956 482600 620978
rect 489932 619970 489960 633490
rect 512000 633480 512052 633486
rect 512000 633422 512052 633428
rect 510620 630896 510672 630902
rect 510620 630838 510672 630844
rect 498016 621784 498068 621790
rect 498016 621726 498068 621732
rect 489932 619942 490314 619970
rect 498028 619956 498056 621726
rect 505744 621716 505796 621722
rect 505744 621658 505796 621664
rect 505756 619956 505784 621658
rect 509884 621036 509936 621042
rect 509884 620978 509936 620984
rect 457442 602712 457498 602721
rect 457442 602647 457498 602656
rect 431222 601760 431278 601769
rect 431222 601695 431278 601704
rect 429474 588024 429530 588033
rect 429474 587959 429530 587968
rect 429382 582720 429438 582729
rect 429382 582655 429438 582664
rect 429290 530292 429346 530301
rect 429290 530227 429346 530236
rect 429200 518968 429252 518974
rect 429200 518910 429252 518916
rect 428372 514752 428424 514758
rect 428372 514694 428424 514700
rect 427820 514684 427872 514690
rect 427820 514626 427872 514632
rect 391938 485072 391994 485081
rect 391938 485007 391994 485016
rect 429396 476814 429424 582655
rect 429488 515710 429516 587959
rect 430670 578368 430726 578377
rect 430670 578303 430726 578312
rect 429566 549400 429622 549409
rect 429566 549335 429622 549344
rect 429580 515778 429608 549335
rect 430578 539608 430634 539617
rect 430578 539543 430634 539552
rect 430592 525026 430620 539543
rect 430580 525020 430632 525026
rect 430580 524962 430632 524968
rect 430578 524920 430634 524929
rect 430578 524855 430634 524864
rect 430592 519790 430620 524855
rect 430684 520169 430712 578303
rect 430762 572792 430818 572801
rect 430762 572727 430818 572736
rect 430670 520160 430726 520169
rect 430670 520095 430726 520104
rect 430580 519784 430632 519790
rect 430580 519726 430632 519732
rect 430776 517206 430804 572727
rect 430854 567760 430910 567769
rect 430854 567695 430910 567704
rect 430868 525178 430896 567695
rect 430946 563136 431002 563145
rect 430946 563071 431002 563080
rect 430960 525298 430988 563071
rect 431038 553480 431094 553489
rect 431038 553415 431094 553424
rect 430948 525292 431000 525298
rect 430948 525234 431000 525240
rect 430868 525150 430988 525178
rect 430856 525020 430908 525026
rect 430856 524962 430908 524968
rect 430868 519994 430896 524962
rect 430960 520062 430988 525150
rect 430948 520056 431000 520062
rect 430948 519998 431000 520004
rect 430856 519988 430908 519994
rect 430856 519930 430908 519936
rect 430764 517200 430816 517206
rect 430764 517142 430816 517148
rect 431052 517138 431080 553415
rect 431130 543960 431186 543969
rect 431130 543895 431186 543904
rect 431144 518158 431172 543895
rect 431236 525434 431264 601695
rect 457442 594552 457498 594561
rect 457442 594487 457498 594496
rect 431314 534440 431370 534449
rect 431314 534375 431370 534384
rect 431224 525428 431276 525434
rect 431224 525370 431276 525376
rect 431224 525292 431276 525298
rect 431224 525234 431276 525240
rect 431236 519858 431264 525234
rect 431328 519926 431356 534375
rect 431408 525428 431460 525434
rect 431408 525370 431460 525376
rect 431316 519920 431368 519926
rect 431316 519862 431368 519868
rect 431224 519852 431276 519858
rect 431224 519794 431276 519800
rect 431420 519722 431448 525370
rect 431408 519716 431460 519722
rect 431408 519658 431460 519664
rect 431132 518152 431184 518158
rect 431132 518094 431184 518100
rect 457456 517274 457484 594487
rect 457534 586392 457590 586401
rect 457534 586327 457590 586336
rect 457548 520130 457576 586327
rect 457626 578232 457682 578241
rect 509896 578202 509924 620978
rect 510632 615641 510660 630838
rect 510618 615632 510674 615641
rect 510618 615567 510674 615576
rect 512012 607481 512040 633422
rect 580170 630864 580226 630873
rect 580170 630799 580172 630808
rect 580224 630799 580226 630808
rect 580172 630770 580224 630776
rect 511998 607472 512054 607481
rect 511998 607407 512054 607416
rect 511998 599312 512054 599321
rect 511998 599247 512054 599256
rect 511262 582992 511318 583001
rect 511262 582927 511318 582936
rect 457626 578167 457682 578176
rect 509884 578196 509936 578202
rect 457640 520198 457668 578167
rect 509884 578138 509936 578144
rect 459572 570030 460046 570058
rect 466472 570030 467774 570058
rect 474752 570030 475502 570058
rect 483032 570030 483230 570058
rect 489932 570030 490958 570058
rect 498212 570030 498686 570058
rect 505112 570030 506414 570058
rect 457628 520192 457680 520198
rect 457628 520134 457680 520140
rect 457536 520124 457588 520130
rect 457536 520066 457588 520072
rect 457444 517268 457496 517274
rect 457444 517210 457496 517216
rect 431040 517132 431092 517138
rect 431040 517074 431092 517080
rect 459572 515846 459600 570030
rect 466472 515914 466500 570030
rect 474752 515982 474780 570030
rect 483032 517342 483060 570030
rect 483020 517336 483072 517342
rect 483020 517278 483072 517284
rect 489932 516050 489960 570030
rect 489920 516044 489972 516050
rect 489920 515986 489972 515992
rect 474740 515976 474792 515982
rect 474740 515918 474792 515924
rect 466460 515908 466512 515914
rect 466460 515850 466512 515856
rect 459560 515840 459612 515846
rect 459560 515782 459612 515788
rect 429568 515772 429620 515778
rect 429568 515714 429620 515720
rect 429476 515704 429528 515710
rect 429476 515646 429528 515652
rect 498212 511970 498240 570030
rect 505112 517478 505140 570030
rect 505100 517472 505152 517478
rect 505100 517414 505152 517420
rect 498200 511964 498252 511970
rect 498200 511906 498252 511912
rect 429384 476808 429436 476814
rect 429384 476750 429436 476756
rect 379336 474700 379388 474706
rect 379336 474642 379388 474648
rect 378784 472660 378836 472666
rect 378784 472602 378836 472608
rect 378140 468512 378192 468518
rect 378140 468454 378192 468460
rect 377864 464568 377916 464574
rect 377864 464510 377916 464516
rect 377772 405680 377824 405686
rect 377772 405622 377824 405628
rect 377772 403640 377824 403646
rect 377772 403582 377824 403588
rect 377784 403209 377812 403582
rect 377770 403200 377826 403209
rect 377770 403135 377826 403144
rect 377678 301064 377734 301073
rect 377678 300999 377734 301008
rect 377784 298217 377812 403135
rect 377876 375358 377904 464510
rect 378048 464500 378100 464506
rect 378048 464442 378100 464448
rect 377864 375352 377916 375358
rect 377864 375294 377916 375300
rect 377956 372156 378008 372162
rect 377956 372098 378008 372104
rect 377864 371952 377916 371958
rect 377864 371894 377916 371900
rect 377876 371414 377904 371894
rect 377968 371550 377996 372098
rect 377956 371544 378008 371550
rect 377956 371486 378008 371492
rect 377864 371408 377916 371414
rect 377864 371350 377916 371356
rect 377770 298208 377826 298217
rect 377770 298143 377826 298152
rect 377784 296714 377812 298143
rect 377692 296686 377812 296714
rect 377586 197840 377642 197849
rect 377586 197775 377642 197784
rect 377494 96928 377550 96937
rect 377494 96863 377550 96872
rect 377600 92857 377628 197775
rect 377692 193225 377720 296686
rect 377772 282260 377824 282266
rect 377772 282202 377824 282208
rect 377784 274174 377812 282202
rect 377772 274168 377824 274174
rect 377772 274110 377824 274116
rect 377876 265946 377904 371350
rect 377968 282266 377996 371486
rect 378060 370666 378088 464442
rect 378140 405680 378192 405686
rect 378140 405622 378192 405628
rect 378152 371686 378180 405622
rect 378140 371680 378192 371686
rect 378140 371622 378192 371628
rect 378152 370802 378180 371622
rect 378140 370796 378192 370802
rect 378140 370738 378192 370744
rect 378048 370660 378100 370666
rect 378048 370602 378100 370608
rect 377956 282260 378008 282266
rect 377956 282202 378008 282208
rect 377956 274168 378008 274174
rect 377956 274110 378008 274116
rect 377864 265940 377916 265946
rect 377864 265882 377916 265888
rect 377968 265538 377996 274110
rect 377956 265532 378008 265538
rect 377956 265474 378008 265480
rect 377968 265198 377996 265474
rect 377956 265192 378008 265198
rect 377956 265134 378008 265140
rect 377956 265056 378008 265062
rect 377956 264998 378008 265004
rect 377862 198792 377918 198801
rect 377862 198727 377918 198736
rect 377770 196072 377826 196081
rect 377770 196007 377826 196016
rect 377678 193216 377734 193225
rect 377678 193151 377734 193160
rect 377586 92848 377642 92857
rect 377586 92783 377642 92792
rect 377310 89992 377366 90001
rect 377310 89927 377366 89936
rect 377692 88233 377720 193151
rect 377784 91089 377812 196007
rect 377876 93809 377904 198727
rect 377968 146198 377996 264998
rect 378060 264926 378088 370602
rect 378692 369572 378744 369578
rect 378692 369514 378744 369520
rect 378704 369034 378732 369514
rect 378692 369028 378744 369034
rect 378692 368970 378744 368976
rect 378692 353388 378744 353394
rect 378692 353330 378744 353336
rect 378600 353320 378652 353326
rect 378600 353262 378652 353268
rect 378612 270502 378640 353262
rect 378600 270496 378652 270502
rect 378506 270464 378562 270473
rect 378600 270438 378652 270444
rect 378506 270399 378562 270408
rect 378048 264920 378100 264926
rect 378048 264862 378100 264868
rect 378060 263634 378088 264862
rect 378048 263628 378100 263634
rect 378048 263570 378100 263576
rect 378046 263528 378102 263537
rect 378046 263463 378048 263472
rect 378100 263463 378102 263472
rect 378048 263434 378100 263440
rect 378414 164248 378470 164257
rect 378414 164183 378470 164192
rect 378428 162994 378456 164183
rect 378416 162988 378468 162994
rect 378416 162930 378468 162936
rect 378048 159928 378100 159934
rect 378048 159870 378100 159876
rect 378060 158817 378088 159870
rect 378046 158808 378102 158817
rect 378046 158743 378102 158752
rect 378048 156664 378100 156670
rect 378048 156606 378100 156612
rect 377956 146192 378008 146198
rect 377956 146134 378008 146140
rect 377956 144900 378008 144906
rect 377956 144842 378008 144848
rect 377968 144129 377996 144842
rect 377954 144120 378010 144129
rect 377954 144055 378010 144064
rect 377968 143721 377996 144055
rect 377954 143712 378010 143721
rect 377954 143647 378010 143656
rect 377862 93800 377918 93809
rect 377862 93735 377918 93744
rect 377770 91080 377826 91089
rect 377770 91015 377826 91024
rect 377678 88224 377734 88233
rect 377678 88159 377734 88168
rect 377312 69012 377364 69018
rect 377312 68954 377364 68960
rect 377324 68105 377352 68954
rect 377310 68096 377366 68105
rect 377310 68031 377366 68040
rect 378060 59702 378088 156606
rect 378048 59696 378100 59702
rect 378048 59638 378100 59644
rect 378428 56438 378456 162930
rect 378520 57866 378548 270399
rect 378704 266286 378732 353330
rect 378692 266280 378744 266286
rect 378692 266222 378744 266228
rect 378600 265736 378652 265742
rect 378600 265678 378652 265684
rect 378612 146198 378640 265678
rect 378704 264994 378732 266222
rect 378692 264988 378744 264994
rect 378692 264930 378744 264936
rect 378692 263628 378744 263634
rect 378692 263570 378744 263576
rect 378704 161474 378732 263570
rect 378796 162042 378824 472602
rect 379152 470280 379204 470286
rect 379152 470222 379204 470228
rect 378876 460216 378928 460222
rect 378876 460158 378928 460164
rect 378784 162036 378836 162042
rect 378784 161978 378836 161984
rect 378888 161945 378916 460158
rect 378968 459196 379020 459202
rect 378968 459138 379020 459144
rect 378980 267617 379008 459138
rect 379060 458992 379112 458998
rect 379060 458934 379112 458940
rect 378966 267608 379022 267617
rect 378966 267543 379022 267552
rect 378966 265568 379022 265577
rect 378966 265503 379022 265512
rect 378980 264790 379008 265503
rect 378968 264784 379020 264790
rect 378968 264726 379020 264732
rect 378874 161936 378930 161945
rect 378874 161871 378930 161880
rect 378704 161446 378916 161474
rect 378600 146192 378652 146198
rect 378600 146134 378652 146140
rect 378888 146033 378916 161446
rect 378980 147626 379008 264726
rect 379072 162353 379100 458934
rect 379164 372774 379192 470222
rect 379244 375352 379296 375358
rect 379244 375294 379296 375300
rect 379256 374610 379284 375294
rect 379244 374604 379296 374610
rect 379244 374546 379296 374552
rect 379152 372768 379204 372774
rect 379152 372710 379204 372716
rect 379152 371816 379204 371822
rect 379152 371758 379204 371764
rect 379164 266082 379192 371758
rect 379256 270337 379284 374546
rect 379348 371890 379376 474642
rect 379980 474632 380032 474638
rect 379980 474574 380032 474580
rect 379428 460828 379480 460834
rect 379428 460770 379480 460776
rect 379440 375018 379468 460770
rect 379428 375012 379480 375018
rect 379428 374954 379480 374960
rect 379796 372768 379848 372774
rect 379796 372710 379848 372716
rect 379808 372638 379836 372710
rect 379796 372632 379848 372638
rect 379796 372574 379848 372580
rect 379520 372224 379572 372230
rect 379520 372166 379572 372172
rect 379336 371884 379388 371890
rect 379336 371826 379388 371832
rect 379348 370002 379376 371826
rect 379532 371686 379560 372166
rect 379520 371680 379572 371686
rect 379520 371622 379572 371628
rect 379704 371680 379756 371686
rect 379704 371622 379756 371628
rect 379348 369974 379468 370002
rect 379336 367940 379388 367946
rect 379336 367882 379388 367888
rect 379242 270328 379298 270337
rect 379242 270263 379298 270272
rect 379256 269482 379284 270263
rect 379244 269476 379296 269482
rect 379244 269418 379296 269424
rect 379152 266076 379204 266082
rect 379152 266018 379204 266024
rect 379164 265130 379192 266018
rect 379152 265124 379204 265130
rect 379152 265066 379204 265072
rect 379244 264988 379296 264994
rect 379244 264930 379296 264936
rect 379058 162344 379114 162353
rect 379058 162279 379114 162288
rect 378968 147620 379020 147626
rect 378968 147562 379020 147568
rect 378968 146192 379020 146198
rect 378968 146134 379020 146140
rect 378874 146024 378930 146033
rect 378692 145988 378744 145994
rect 378874 145959 378930 145968
rect 378692 145930 378744 145936
rect 378600 145512 378652 145518
rect 378600 145454 378652 145460
rect 378612 144838 378640 145454
rect 378704 145450 378732 145930
rect 378692 145444 378744 145450
rect 378692 145386 378744 145392
rect 378600 144832 378652 144838
rect 378600 144774 378652 144780
rect 378612 59770 378640 144774
rect 378704 59838 378732 145386
rect 378784 145376 378836 145382
rect 378784 145318 378836 145324
rect 378692 59832 378744 59838
rect 378692 59774 378744 59780
rect 378600 59764 378652 59770
rect 378600 59706 378652 59712
rect 378796 59634 378824 145318
rect 378784 59628 378836 59634
rect 378784 59570 378836 59576
rect 378508 57860 378560 57866
rect 378508 57802 378560 57808
rect 378416 56432 378468 56438
rect 378416 56374 378468 56380
rect 378888 56098 378916 145959
rect 378980 145858 379008 146134
rect 379256 145994 379284 264930
rect 379348 264858 379376 367882
rect 379440 266966 379468 369974
rect 379520 270496 379572 270502
rect 379520 270438 379572 270444
rect 379532 269414 379560 270438
rect 379520 269408 379572 269414
rect 379520 269350 379572 269356
rect 379428 266960 379480 266966
rect 379428 266902 379480 266908
rect 379336 264852 379388 264858
rect 379336 264794 379388 264800
rect 379348 263634 379376 264794
rect 379336 263628 379388 263634
rect 379336 263570 379388 263576
rect 379440 161474 379468 266902
rect 379348 161446 379468 161474
rect 379348 161294 379376 161446
rect 379532 161362 379560 269350
rect 379716 266218 379744 371622
rect 379808 266354 379836 372574
rect 379992 372162 380020 474574
rect 511276 462233 511304 582927
rect 512012 520266 512040 599247
rect 512090 591152 512146 591161
rect 512090 591087 512146 591096
rect 512000 520260 512052 520266
rect 512000 520202 512052 520208
rect 512104 516118 512132 591087
rect 580172 578196 580224 578202
rect 580172 578138 580224 578144
rect 580184 577697 580212 578138
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 512182 574832 512238 574841
rect 512182 574767 512238 574776
rect 512196 517410 512224 574767
rect 512184 517404 512236 517410
rect 512184 517346 512236 517352
rect 519544 516180 519596 516186
rect 519544 516122 519596 516128
rect 512092 516112 512144 516118
rect 512092 516054 512144 516060
rect 511262 462224 511318 462233
rect 511262 462159 511318 462168
rect 511276 461922 511304 462159
rect 511264 461916 511316 461922
rect 511264 461858 511316 461864
rect 517520 461916 517572 461922
rect 517520 461858 517572 461864
rect 498384 461100 498436 461106
rect 498384 461042 498436 461048
rect 498396 461009 498424 461042
rect 499856 461032 499908 461038
rect 498382 461000 498438 461009
rect 498382 460935 498384 460944
rect 498436 460935 498438 460944
rect 499854 461000 499856 461009
rect 499908 461000 499910 461009
rect 499854 460935 499910 460944
rect 498384 460906 498436 460912
rect 516600 458312 516652 458318
rect 516600 458254 516652 458260
rect 516612 454753 516640 458254
rect 516598 454744 516654 454753
rect 516598 454679 516654 454688
rect 405922 375048 405978 375057
rect 380900 375012 380952 375018
rect 405922 374983 405978 374992
rect 407762 375048 407818 375057
rect 407762 374983 407818 374992
rect 425058 375048 425114 375057
rect 425058 374983 425114 374992
rect 440330 375048 440386 375057
rect 440330 374983 440386 374992
rect 443090 375048 443146 375057
rect 443090 374983 443146 374992
rect 452842 375048 452898 375057
rect 452842 374983 452898 374992
rect 380900 374954 380952 374960
rect 380912 374066 380940 374954
rect 405936 374066 405964 374983
rect 407776 374474 407804 374983
rect 410706 374640 410762 374649
rect 425072 374610 425100 374983
rect 410706 374575 410762 374584
rect 425060 374604 425112 374610
rect 410720 374542 410748 374575
rect 425060 374546 425112 374552
rect 410708 374536 410760 374542
rect 410708 374478 410760 374484
rect 433614 374504 433670 374513
rect 407764 374468 407816 374474
rect 433614 374439 433670 374448
rect 436006 374504 436062 374513
rect 436006 374439 436062 374448
rect 438490 374504 438546 374513
rect 438490 374439 438546 374448
rect 407764 374410 407816 374416
rect 433628 374202 433656 374439
rect 436020 374270 436048 374439
rect 438504 374406 438532 374439
rect 438492 374400 438544 374406
rect 438492 374342 438544 374348
rect 440344 374338 440372 374983
rect 440332 374332 440384 374338
rect 440332 374274 440384 374280
rect 436008 374264 436060 374270
rect 436008 374206 436060 374212
rect 433616 374196 433668 374202
rect 433616 374138 433668 374144
rect 443104 374134 443132 374983
rect 452856 374746 452884 374983
rect 452844 374740 452896 374746
rect 452844 374682 452896 374688
rect 443092 374128 443144 374134
rect 416042 374096 416098 374105
rect 380900 374060 380952 374066
rect 380900 374002 380952 374008
rect 405924 374060 405976 374066
rect 443092 374070 443144 374076
rect 416042 374031 416098 374040
rect 405924 374002 405976 374008
rect 379980 372156 380032 372162
rect 379980 372098 380032 372104
rect 379888 370592 379940 370598
rect 379888 370534 379940 370540
rect 379900 267918 379928 370534
rect 379888 267912 379940 267918
rect 379888 267854 379940 267860
rect 379796 266348 379848 266354
rect 379796 266290 379848 266296
rect 379704 266212 379756 266218
rect 379704 266154 379756 266160
rect 379716 265062 379744 266154
rect 379808 265334 379836 266290
rect 379796 265328 379848 265334
rect 379796 265270 379848 265276
rect 379704 265056 379756 265062
rect 379704 264998 379756 265004
rect 379900 258074 379928 267854
rect 379992 267073 380020 372098
rect 380912 354006 380940 374002
rect 416056 373862 416084 374031
rect 416044 373856 416096 373862
rect 416044 373798 416096 373804
rect 418252 373788 418304 373794
rect 418252 373730 418304 373736
rect 418264 373697 418292 373730
rect 423036 373720 423088 373726
rect 418250 373688 418306 373697
rect 418250 373623 418306 373632
rect 423034 373688 423036 373697
rect 423088 373688 423090 373697
rect 423034 373623 423090 373632
rect 426898 373688 426954 373697
rect 426898 373623 426900 373632
rect 426952 373623 426954 373632
rect 445850 373688 445906 373697
rect 445850 373623 445906 373632
rect 426900 373594 426952 373600
rect 445864 373590 445892 373623
rect 445852 373584 445904 373590
rect 445852 373526 445904 373532
rect 450266 373552 450322 373561
rect 450266 373487 450268 373496
rect 450320 373487 450322 373496
rect 455418 373552 455474 373561
rect 455418 373487 455474 373496
rect 450268 373458 450320 373464
rect 455432 373454 455460 373487
rect 455420 373448 455472 373454
rect 447690 373416 447746 373425
rect 455420 373390 455472 373396
rect 462778 373416 462834 373425
rect 447690 373351 447692 373360
rect 447744 373351 447746 373360
rect 462778 373351 462834 373360
rect 447692 373322 447744 373328
rect 462792 373318 462820 373351
rect 462780 373312 462832 373318
rect 462780 373254 462832 373260
rect 402888 372632 402940 372638
rect 400218 372600 400274 372609
rect 400218 372535 400274 372544
rect 402886 372600 402888 372609
rect 402940 372600 402942 372609
rect 402886 372535 402942 372544
rect 400232 372366 400260 372535
rect 400220 372360 400272 372366
rect 400220 372302 400272 372308
rect 470598 372328 470654 372337
rect 470598 372263 470654 372272
rect 396078 372192 396134 372201
rect 396078 372127 396080 372136
rect 396132 372127 396134 372136
rect 396080 372098 396132 372104
rect 380992 372088 381044 372094
rect 380992 372030 381044 372036
rect 397458 372056 397514 372065
rect 381004 371550 381032 372030
rect 397458 371991 397460 372000
rect 397512 371991 397514 372000
rect 404358 372056 404414 372065
rect 404358 371991 404414 372000
rect 407118 372056 407174 372065
rect 407118 371991 407174 372000
rect 422298 372056 422354 372065
rect 422298 371991 422354 372000
rect 397460 371962 397512 371968
rect 404372 371958 404400 371991
rect 404360 371952 404412 371958
rect 404360 371894 404412 371900
rect 407132 371822 407160 371991
rect 422312 371890 422340 371991
rect 422300 371884 422352 371890
rect 422300 371826 422352 371832
rect 407120 371816 407172 371822
rect 401598 371784 401654 371793
rect 407120 371758 407172 371764
rect 409878 371784 409934 371793
rect 401598 371719 401600 371728
rect 401652 371719 401654 371728
rect 409878 371719 409934 371728
rect 401600 371690 401652 371696
rect 409892 371686 409920 371719
rect 409880 371680 409932 371686
rect 398838 371648 398894 371657
rect 409880 371622 409932 371628
rect 411258 371648 411314 371657
rect 398838 371583 398840 371592
rect 398892 371583 398894 371592
rect 411258 371583 411314 371592
rect 465078 371648 465134 371657
rect 465078 371583 465134 371592
rect 398840 371554 398892 371560
rect 411272 371550 411300 371583
rect 380992 371544 381044 371550
rect 411260 371544 411312 371550
rect 381044 371492 381124 371498
rect 380992 371486 381124 371492
rect 411260 371486 411312 371492
rect 411350 371512 411406 371521
rect 381004 371470 381124 371486
rect 380992 371408 381044 371414
rect 380992 371350 381044 371356
rect 380900 354000 380952 354006
rect 380900 353942 380952 353948
rect 381004 353326 381032 371350
rect 381096 353394 381124 371470
rect 411350 371447 411352 371456
rect 411404 371447 411406 371456
rect 418250 371512 418306 371521
rect 418250 371447 418306 371456
rect 421010 371512 421066 371521
rect 421010 371447 421066 371456
rect 423678 371512 423734 371521
rect 423678 371447 423734 371456
rect 426438 371512 426494 371521
rect 426438 371447 426494 371456
rect 430670 371512 430726 371521
rect 430670 371447 430726 371456
rect 411352 371418 411404 371424
rect 396078 371376 396134 371385
rect 396078 371311 396134 371320
rect 402978 371376 403034 371385
rect 402978 371311 403034 371320
rect 412638 371376 412694 371385
rect 412638 371311 412694 371320
rect 413190 371376 413246 371385
rect 413190 371311 413246 371320
rect 414018 371376 414074 371385
rect 414018 371311 414074 371320
rect 415398 371376 415454 371385
rect 415398 371311 415454 371320
rect 416778 371376 416834 371385
rect 416778 371311 416834 371320
rect 418158 371376 418214 371385
rect 418158 371311 418214 371320
rect 396092 370394 396120 371311
rect 402992 370462 403020 371311
rect 402980 370456 403032 370462
rect 402980 370398 403032 370404
rect 396080 370388 396132 370394
rect 396080 370330 396132 370336
rect 412652 367946 412680 371311
rect 413204 370734 413232 371311
rect 413192 370728 413244 370734
rect 413192 370670 413244 370676
rect 414032 370598 414060 371311
rect 414020 370592 414072 370598
rect 414020 370534 414072 370540
rect 415412 370530 415440 371311
rect 416792 370666 416820 371311
rect 416780 370660 416832 370666
rect 416780 370602 416832 370608
rect 415400 370524 415452 370530
rect 415400 370466 415452 370472
rect 418172 369306 418200 371311
rect 418160 369300 418212 369306
rect 418160 369242 418212 369248
rect 418264 369102 418292 371447
rect 419538 371376 419594 371385
rect 419538 371311 419594 371320
rect 420918 371376 420974 371385
rect 420918 371311 420974 371320
rect 419552 369238 419580 371311
rect 420932 369442 420960 371311
rect 420920 369436 420972 369442
rect 420920 369378 420972 369384
rect 419540 369232 419592 369238
rect 419540 369174 419592 369180
rect 421024 369170 421052 371447
rect 423692 369374 423720 371447
rect 426452 371414 426480 371447
rect 426440 371408 426492 371414
rect 425058 371376 425114 371385
rect 426440 371350 426492 371356
rect 427818 371376 427874 371385
rect 425058 371311 425114 371320
rect 427818 371311 427874 371320
rect 429198 371376 429254 371385
rect 429198 371311 429254 371320
rect 430578 371376 430634 371385
rect 430578 371311 430634 371320
rect 425072 369646 425100 371311
rect 427832 370802 427860 371311
rect 427820 370796 427872 370802
rect 427820 370738 427872 370744
rect 425060 369640 425112 369646
rect 425060 369582 425112 369588
rect 429212 369510 429240 371311
rect 430592 369714 430620 371311
rect 430580 369708 430632 369714
rect 430580 369650 430632 369656
rect 430684 369578 430712 371447
rect 431958 371376 432014 371385
rect 431958 371311 432014 371320
rect 433338 371376 433394 371385
rect 433338 371311 433394 371320
rect 434718 371376 434774 371385
rect 434718 371311 434774 371320
rect 436098 371376 436154 371385
rect 436098 371311 436154 371320
rect 458178 371376 458234 371385
rect 458178 371311 458234 371320
rect 430672 369572 430724 369578
rect 430672 369514 430724 369520
rect 429200 369504 429252 369510
rect 429200 369446 429252 369452
rect 423680 369368 423732 369374
rect 423680 369310 423732 369316
rect 421012 369164 421064 369170
rect 421012 369106 421064 369112
rect 418252 369096 418304 369102
rect 418252 369038 418304 369044
rect 412640 367940 412692 367946
rect 412640 367882 412692 367888
rect 431972 367878 432000 371311
rect 431960 367872 432012 367878
rect 431960 367814 432012 367820
rect 433352 367810 433380 371311
rect 434732 368422 434760 371311
rect 436112 368490 436140 371311
rect 458192 370870 458220 371311
rect 465092 371006 465120 371583
rect 465080 371000 465132 371006
rect 465080 370942 465132 370948
rect 470612 370938 470640 372263
rect 503166 372192 503222 372201
rect 503166 372127 503222 372136
rect 503534 372192 503590 372201
rect 503534 372127 503590 372136
rect 483018 371920 483074 371929
rect 483018 371855 483074 371864
rect 473358 371376 473414 371385
rect 473358 371311 473414 371320
rect 474738 371376 474794 371385
rect 474738 371311 474794 371320
rect 477498 371376 477554 371385
rect 477498 371311 477554 371320
rect 480258 371376 480314 371385
rect 480258 371311 480314 371320
rect 473372 371074 473400 371311
rect 474752 371142 474780 371311
rect 477512 371210 477540 371311
rect 477500 371204 477552 371210
rect 477500 371146 477552 371152
rect 474740 371136 474792 371142
rect 474740 371078 474792 371084
rect 473360 371068 473412 371074
rect 473360 371010 473412 371016
rect 470600 370932 470652 370938
rect 470600 370874 470652 370880
rect 458180 370864 458232 370870
rect 458180 370806 458232 370812
rect 480272 369850 480300 371311
rect 480260 369844 480312 369850
rect 480260 369786 480312 369792
rect 483032 369782 483060 371855
rect 503180 371278 503208 372127
rect 503548 371346 503576 372127
rect 503536 371340 503588 371346
rect 503536 371282 503588 371288
rect 503168 371272 503220 371278
rect 503168 371214 503220 371220
rect 483020 369776 483072 369782
rect 483020 369718 483072 369724
rect 436100 368484 436152 368490
rect 436100 368426 436152 368432
rect 434720 368416 434772 368422
rect 434720 368358 434772 368364
rect 433340 367804 433392 367810
rect 433340 367746 433392 367752
rect 500868 355496 500920 355502
rect 500868 355438 500920 355444
rect 498844 355428 498896 355434
rect 498844 355370 498896 355376
rect 498856 355065 498884 355370
rect 498842 355056 498898 355065
rect 498842 354991 498898 355000
rect 500880 354929 500908 355438
rect 500866 354920 500922 354929
rect 500866 354855 500922 354864
rect 510894 354784 510950 354793
rect 517532 354754 517560 461858
rect 517612 461032 517664 461038
rect 517612 460974 517664 460980
rect 517624 355502 517652 460974
rect 517704 460964 517756 460970
rect 517704 460906 517756 460912
rect 517612 355496 517664 355502
rect 517612 355438 517664 355444
rect 510894 354719 510896 354728
rect 510948 354719 510950 354728
rect 517520 354748 517572 354754
rect 510896 354690 510948 354696
rect 517520 354690 517572 354696
rect 381084 353388 381136 353394
rect 381084 353330 381136 353336
rect 380992 353320 381044 353326
rect 380992 353262 381044 353268
rect 418434 269784 418490 269793
rect 418434 269719 418490 269728
rect 425242 269784 425298 269793
rect 425242 269719 425298 269728
rect 418448 269346 418476 269719
rect 423494 269648 423550 269657
rect 423494 269583 423550 269592
rect 418436 269340 418488 269346
rect 418436 269282 418488 269288
rect 396080 268932 396132 268938
rect 396080 268874 396132 268880
rect 396092 268054 396120 268874
rect 423508 268870 423536 269583
rect 425256 269482 425284 269719
rect 426438 269648 426494 269657
rect 426438 269583 426494 269592
rect 433614 269648 433670 269657
rect 433614 269583 433670 269592
rect 453394 269648 453450 269657
rect 453394 269583 453450 269592
rect 468482 269648 468538 269657
rect 468482 269583 468538 269592
rect 480902 269648 480958 269657
rect 480902 269583 480958 269592
rect 425244 269476 425296 269482
rect 425244 269418 425296 269424
rect 426452 269414 426480 269583
rect 426440 269408 426492 269414
rect 426440 269350 426492 269356
rect 433628 269278 433656 269583
rect 433616 269272 433668 269278
rect 433616 269214 433668 269220
rect 453408 269210 453436 269583
rect 453396 269204 453448 269210
rect 453396 269146 453448 269152
rect 468496 269142 468524 269583
rect 468484 269136 468536 269142
rect 468484 269078 468536 269084
rect 430946 268968 431002 268977
rect 430946 268903 431002 268912
rect 433338 268968 433394 268977
rect 433338 268903 433394 268912
rect 475842 268968 475898 268977
rect 475842 268903 475898 268912
rect 478418 268968 478474 268977
rect 478418 268903 478474 268912
rect 423496 268864 423548 268870
rect 415858 268832 415914 268841
rect 415858 268767 415914 268776
rect 421010 268832 421066 268841
rect 423496 268806 423548 268812
rect 421010 268767 421012 268776
rect 398194 268152 398250 268161
rect 398194 268087 398250 268096
rect 401690 268152 401746 268161
rect 401690 268087 401746 268096
rect 396080 268048 396132 268054
rect 396080 267990 396132 267996
rect 379978 267064 380034 267073
rect 379978 266999 380034 267008
rect 379992 265266 380020 266999
rect 388166 265296 388222 265305
rect 379980 265260 380032 265266
rect 388166 265231 388222 265240
rect 379980 265202 380032 265208
rect 388180 264790 388208 265231
rect 389178 265160 389234 265169
rect 389178 265095 389234 265104
rect 388168 264784 388220 264790
rect 388168 264726 388220 264732
rect 389192 264722 389220 265095
rect 390558 265024 390614 265033
rect 390558 264959 390614 264968
rect 391940 264988 391992 264994
rect 389180 264716 389232 264722
rect 389180 264658 389232 264664
rect 390572 264654 390600 264959
rect 391940 264930 391992 264936
rect 390560 264648 390612 264654
rect 390560 264590 390612 264596
rect 391952 264586 391980 264930
rect 391940 264580 391992 264586
rect 391940 264522 391992 264528
rect 379624 258046 379928 258074
rect 379520 161356 379572 161362
rect 379520 161298 379572 161304
rect 379336 161288 379388 161294
rect 379336 161230 379388 161236
rect 379244 145988 379296 145994
rect 379244 145930 379296 145936
rect 378968 145852 379020 145858
rect 378968 145794 379020 145800
rect 378876 56092 378928 56098
rect 378876 56034 378928 56040
rect 378980 55962 379008 145794
rect 379256 142154 379284 145930
rect 379164 142126 379284 142154
rect 379164 56030 379192 142126
rect 379348 59566 379376 161230
rect 379532 160138 379560 161298
rect 379520 160132 379572 160138
rect 379520 160074 379572 160080
rect 379428 147620 379480 147626
rect 379428 147562 379480 147568
rect 379336 59560 379388 59566
rect 379336 59502 379388 59508
rect 379440 56302 379468 147562
rect 379624 146198 379652 258046
rect 396092 250510 396120 267990
rect 398208 265878 398236 268087
rect 398838 266384 398894 266393
rect 398838 266319 398894 266328
rect 400218 266384 400274 266393
rect 400218 266319 400274 266328
rect 398196 265872 398248 265878
rect 398196 265814 398248 265820
rect 398852 265810 398880 266319
rect 400232 266014 400260 266319
rect 401704 266150 401732 268087
rect 415872 268054 415900 268767
rect 421064 268767 421066 268776
rect 421012 268738 421064 268744
rect 430960 268734 430988 268903
rect 430948 268728 431000 268734
rect 430948 268670 431000 268676
rect 416042 268152 416098 268161
rect 433352 268122 433380 268903
rect 475856 268598 475884 268903
rect 478432 268666 478460 268903
rect 478420 268660 478472 268666
rect 478420 268602 478472 268608
rect 475844 268592 475896 268598
rect 475844 268534 475896 268540
rect 473360 268524 473412 268530
rect 473360 268466 473412 268472
rect 434258 268152 434314 268161
rect 416042 268087 416098 268096
rect 433340 268116 433392 268122
rect 415860 268048 415912 268054
rect 415860 267990 415912 267996
rect 402980 267980 403032 267986
rect 402980 267922 403032 267928
rect 402992 267753 403020 267922
rect 414388 267912 414440 267918
rect 414388 267854 414440 267860
rect 414400 267753 414428 267854
rect 402978 267744 403034 267753
rect 402978 267679 403034 267688
rect 414386 267744 414442 267753
rect 414386 267679 414442 267688
rect 416056 267102 416084 268087
rect 434258 268087 434314 268096
rect 455786 268152 455842 268161
rect 455786 268087 455842 268096
rect 433340 268058 433392 268064
rect 421564 267912 421616 267918
rect 421564 267854 421616 267860
rect 416044 267096 416096 267102
rect 407118 267064 407174 267073
rect 407118 266999 407174 267008
rect 409878 267064 409934 267073
rect 409878 266999 409880 267008
rect 407132 266830 407160 266999
rect 409932 266999 409934 267008
rect 412914 267064 412970 267073
rect 416044 267038 416096 267044
rect 412914 266999 412970 267008
rect 409880 266970 409932 266976
rect 412928 266898 412956 266999
rect 412916 266892 412968 266898
rect 412916 266834 412968 266840
rect 407120 266824 407172 266830
rect 407120 266766 407172 266772
rect 411350 266520 411406 266529
rect 411350 266455 411406 266464
rect 418250 266520 418306 266529
rect 418250 266455 418306 266464
rect 403162 266384 403218 266393
rect 403162 266319 403164 266328
rect 403216 266319 403218 266328
rect 404358 266384 404414 266393
rect 404358 266319 404414 266328
rect 405738 266384 405794 266393
rect 405738 266319 405794 266328
rect 407118 266384 407174 266393
rect 407118 266319 407174 266328
rect 408498 266384 408554 266393
rect 408498 266319 408554 266328
rect 409878 266384 409934 266393
rect 409878 266319 409934 266328
rect 411258 266384 411314 266393
rect 411258 266319 411314 266328
rect 403164 266290 403216 266296
rect 401692 266144 401744 266150
rect 401692 266086 401744 266092
rect 400220 266008 400272 266014
rect 400220 265950 400272 265956
rect 404372 265946 404400 266319
rect 404360 265940 404412 265946
rect 404360 265882 404412 265888
rect 398840 265804 398892 265810
rect 398840 265746 398892 265752
rect 405752 265674 405780 266319
rect 407132 266082 407160 266319
rect 407120 266076 407172 266082
rect 407120 266018 407172 266024
rect 408512 265742 408540 266319
rect 409892 266218 409920 266319
rect 411272 266286 411300 266319
rect 411260 266280 411312 266286
rect 411260 266222 411312 266228
rect 409880 266212 409932 266218
rect 409880 266154 409932 266160
rect 408500 265736 408552 265742
rect 408500 265678 408552 265684
rect 405740 265668 405792 265674
rect 405740 265610 405792 265616
rect 411364 265538 411392 266455
rect 412914 266384 412970 266393
rect 412914 266319 412970 266328
rect 416778 266384 416834 266393
rect 416778 266319 416834 266328
rect 418158 266384 418214 266393
rect 418158 266319 418214 266328
rect 411352 265532 411404 265538
rect 411352 265474 411404 265480
rect 412928 264858 412956 266319
rect 416792 264926 416820 266319
rect 416780 264920 416832 264926
rect 416780 264862 416832 264868
rect 412916 264852 412968 264858
rect 412916 264794 412968 264800
rect 418172 264586 418200 266319
rect 418264 264654 418292 266455
rect 419538 266384 419594 266393
rect 419538 266319 419594 266328
rect 420918 266384 420974 266393
rect 420918 266319 420974 266328
rect 419552 264722 419580 266319
rect 420932 264790 420960 266319
rect 420920 264784 420972 264790
rect 420920 264726 420972 264732
rect 419540 264716 419592 264722
rect 419540 264658 419592 264664
rect 418252 264648 418304 264654
rect 418252 264590 418304 264596
rect 418160 264580 418212 264586
rect 418160 264522 418212 264528
rect 421576 251122 421604 267854
rect 432144 267844 432196 267850
rect 432144 267786 432196 267792
rect 432156 267753 432184 267786
rect 432142 267744 432198 267753
rect 432142 267679 432198 267688
rect 422574 267064 422630 267073
rect 422574 266999 422630 267008
rect 422588 266966 422616 266999
rect 422576 266960 422628 266966
rect 422576 266902 422628 266908
rect 434272 266422 434300 268087
rect 435732 267912 435784 267918
rect 435732 267854 435784 267860
rect 435744 267753 435772 267854
rect 435730 267744 435786 267753
rect 435730 267679 435786 267688
rect 435914 267744 435970 267753
rect 435914 267679 435970 267688
rect 445758 267744 445814 267753
rect 445758 267679 445814 267688
rect 447138 267744 447194 267753
rect 447138 267679 447194 267688
rect 449898 267744 449954 267753
rect 449898 267679 449954 267688
rect 435928 267374 435956 267679
rect 445772 267578 445800 267679
rect 445760 267572 445812 267578
rect 445760 267514 445812 267520
rect 447152 267442 447180 267679
rect 449912 267510 449940 267679
rect 455800 267646 455828 268087
rect 473372 267753 473400 268466
rect 480916 268462 480944 269583
rect 483386 268968 483442 268977
rect 483386 268903 483442 268912
rect 480904 268456 480956 268462
rect 480904 268398 480956 268404
rect 483400 268394 483428 268903
rect 483388 268388 483440 268394
rect 483388 268330 483440 268336
rect 458178 267744 458234 267753
rect 458178 267679 458180 267688
rect 458232 267679 458234 267688
rect 473358 267744 473414 267753
rect 473358 267679 473414 267688
rect 458180 267650 458232 267656
rect 455788 267640 455840 267646
rect 455788 267582 455840 267588
rect 449900 267504 449952 267510
rect 449900 267446 449952 267452
rect 503534 267472 503590 267481
rect 447140 267436 447192 267442
rect 503534 267407 503590 267416
rect 447140 267378 447192 267384
rect 435916 267368 435968 267374
rect 435916 267310 435968 267316
rect 437478 267336 437534 267345
rect 437478 267271 437480 267280
rect 437532 267271 437534 267280
rect 442998 267336 443054 267345
rect 442998 267271 443054 267280
rect 503442 267336 503498 267345
rect 503442 267271 503498 267280
rect 437480 267242 437532 267248
rect 443012 267238 443040 267271
rect 443000 267232 443052 267238
rect 440238 267200 440294 267209
rect 443000 267174 443052 267180
rect 440238 267135 440240 267144
rect 440292 267135 440294 267144
rect 440240 267106 440292 267112
rect 503456 267034 503484 267271
rect 503548 267170 503576 267407
rect 503536 267164 503588 267170
rect 503536 267106 503588 267112
rect 503444 267028 503496 267034
rect 503444 266970 503496 266976
rect 425704 266416 425756 266422
rect 434260 266416 434312 266422
rect 425704 266358 425756 266364
rect 429106 266384 429162 266393
rect 421564 251116 421616 251122
rect 421564 251058 421616 251064
rect 425716 250782 425744 266358
rect 430486 266384 430542 266393
rect 429162 266342 429240 266370
rect 429106 266319 429162 266328
rect 425704 250776 425756 250782
rect 425704 250718 425756 250724
rect 429212 250646 429240 266342
rect 430670 266384 430726 266393
rect 430542 266342 430620 266370
rect 430486 266319 430542 266328
rect 430592 251190 430620 266342
rect 434260 266358 434312 266364
rect 436098 266384 436154 266393
rect 430670 266319 430726 266328
rect 436098 266319 436154 266328
rect 437478 266384 437534 266393
rect 437478 266319 437534 266328
rect 438858 266384 438914 266393
rect 438858 266319 438914 266328
rect 430580 251184 430632 251190
rect 430580 251126 430632 251132
rect 430684 250714 430712 266319
rect 436112 263566 436140 266319
rect 436100 263560 436152 263566
rect 436100 263502 436152 263508
rect 437492 263498 437520 266319
rect 437480 263492 437532 263498
rect 437480 263434 437532 263440
rect 430672 250708 430724 250714
rect 430672 250650 430724 250656
rect 429200 250640 429252 250646
rect 429200 250582 429252 250588
rect 438872 250578 438900 266319
rect 500408 250640 500460 250646
rect 500408 250582 500460 250588
rect 438860 250572 438912 250578
rect 438860 250514 438912 250520
rect 499028 250572 499080 250578
rect 499028 250514 499080 250520
rect 379704 250504 379756 250510
rect 379704 250446 379756 250452
rect 396080 250504 396132 250510
rect 396080 250446 396132 250452
rect 379612 146192 379664 146198
rect 379716 146169 379744 250446
rect 499040 249937 499068 250514
rect 500420 249937 500448 250582
rect 499026 249928 499082 249937
rect 499026 249863 499082 249872
rect 500406 249928 500462 249937
rect 500406 249863 500462 249872
rect 510894 249928 510950 249937
rect 517532 249898 517560 354690
rect 517624 251122 517652 355438
rect 517716 355434 517744 460906
rect 519556 454714 519584 516122
rect 580264 515432 580316 515438
rect 580264 515374 580316 515380
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 520924 487212 520976 487218
rect 520924 487154 520976 487160
rect 519544 454708 519596 454714
rect 519544 454650 519596 454656
rect 518898 454200 518954 454209
rect 518898 454135 518954 454144
rect 518440 371884 518492 371890
rect 518440 371826 518492 371832
rect 518452 371346 518480 371826
rect 517888 371340 517940 371346
rect 517888 371282 517940 371288
rect 518440 371340 518492 371346
rect 518440 371282 518492 371288
rect 517704 355428 517756 355434
rect 517704 355370 517756 355376
rect 517716 354674 517744 355370
rect 517716 354646 517836 354674
rect 517704 266416 517756 266422
rect 517704 266358 517756 266364
rect 517612 251116 517664 251122
rect 517612 251058 517664 251064
rect 510894 249863 510896 249872
rect 510948 249863 510950 249872
rect 517520 249892 517572 249898
rect 510896 249834 510948 249840
rect 517520 249834 517572 249840
rect 425978 164792 426034 164801
rect 425978 164727 426034 164736
rect 434350 164792 434406 164801
rect 434350 164727 434406 164736
rect 451002 164792 451058 164801
rect 451002 164727 451058 164736
rect 423494 164656 423550 164665
rect 423494 164591 423550 164600
rect 416042 164248 416098 164257
rect 416042 164183 416098 164192
rect 421010 164248 421066 164257
rect 421010 164183 421066 164192
rect 393320 164144 393372 164150
rect 393320 164086 393372 164092
rect 394516 164144 394568 164150
rect 394516 164086 394568 164092
rect 379888 160132 379940 160138
rect 379888 160074 379940 160080
rect 379796 146192 379848 146198
rect 379612 146134 379664 146140
rect 379702 146160 379758 146169
rect 379796 146134 379848 146140
rect 379702 146095 379758 146104
rect 379716 57254 379744 146095
rect 379704 57248 379756 57254
rect 379704 57190 379756 57196
rect 379428 56296 379480 56302
rect 379428 56238 379480 56244
rect 379808 56166 379836 146134
rect 379900 56234 379928 160074
rect 379980 148368 380032 148374
rect 379980 148310 380032 148316
rect 379888 56228 379940 56234
rect 379888 56170 379940 56176
rect 379796 56160 379848 56166
rect 379796 56102 379848 56108
rect 379152 56024 379204 56030
rect 379152 55966 379204 55972
rect 378968 55956 379020 55962
rect 378968 55898 379020 55904
rect 379992 54874 380020 148310
rect 393332 145382 393360 164086
rect 394528 163130 394556 164086
rect 416056 163946 416084 164183
rect 421024 164014 421052 164183
rect 423508 164082 423536 164591
rect 425992 164422 426020 164727
rect 434364 164490 434392 164727
rect 436926 164656 436982 164665
rect 436926 164591 436982 164600
rect 438030 164656 438086 164665
rect 438030 164591 438086 164600
rect 434352 164484 434404 164490
rect 434352 164426 434404 164432
rect 425980 164416 426032 164422
rect 425980 164358 426032 164364
rect 428186 164248 428242 164257
rect 428186 164183 428242 164192
rect 430946 164248 431002 164257
rect 430946 164183 431002 164192
rect 423496 164076 423548 164082
rect 423496 164018 423548 164024
rect 421012 164008 421064 164014
rect 421012 163950 421064 163956
rect 416044 163940 416096 163946
rect 416044 163882 416096 163888
rect 428200 163878 428228 164183
rect 428188 163872 428240 163878
rect 428188 163814 428240 163820
rect 430960 163810 430988 164183
rect 430948 163804 431000 163810
rect 430948 163746 431000 163752
rect 396724 163192 396776 163198
rect 396724 163134 396776 163140
rect 401598 163160 401654 163169
rect 394516 163124 394568 163130
rect 394516 163066 394568 163072
rect 396078 162752 396134 162761
rect 396078 162687 396134 162696
rect 396092 145518 396120 162687
rect 396170 162208 396226 162217
rect 396170 162143 396226 162152
rect 396080 145512 396132 145518
rect 396080 145454 396132 145460
rect 396184 145450 396212 162143
rect 396736 146130 396764 163134
rect 401598 163095 401654 163104
rect 415308 163124 415360 163130
rect 397458 162752 397514 162761
rect 397458 162687 397514 162696
rect 398838 162752 398894 162761
rect 398838 162687 398894 162696
rect 400218 162752 400274 162761
rect 400218 162687 400274 162696
rect 397472 148510 397500 162687
rect 397460 148504 397512 148510
rect 397460 148446 397512 148452
rect 398852 148442 398880 162687
rect 400232 148918 400260 162687
rect 401612 148986 401640 163095
rect 415308 163066 415360 163072
rect 415320 162858 415348 163066
rect 431960 163056 432012 163062
rect 431960 162998 432012 163004
rect 418158 162888 418214 162897
rect 415308 162852 415360 162858
rect 418158 162823 418160 162832
rect 415308 162794 415360 162800
rect 418212 162823 418214 162832
rect 418160 162794 418212 162800
rect 431972 162761 432000 162998
rect 436940 162926 436968 164591
rect 438044 162994 438072 164591
rect 451016 164354 451044 164727
rect 480902 164656 480958 164665
rect 480902 164591 480958 164600
rect 451004 164348 451056 164354
rect 451004 164290 451056 164296
rect 480916 164286 480944 164591
rect 480904 164280 480956 164286
rect 473450 164248 473506 164257
rect 473450 164183 473506 164192
rect 475842 164248 475898 164257
rect 475842 164183 475898 164192
rect 478418 164248 478474 164257
rect 480904 164222 480956 164228
rect 478418 164183 478474 164192
rect 470598 163840 470654 163849
rect 470598 163775 470654 163784
rect 470612 163742 470640 163775
rect 470600 163736 470652 163742
rect 470600 163678 470652 163684
rect 473464 163674 473492 164183
rect 473452 163668 473504 163674
rect 473452 163610 473504 163616
rect 475856 163606 475884 164183
rect 475844 163600 475896 163606
rect 475844 163542 475896 163548
rect 478432 163538 478460 164183
rect 517532 163674 517560 249834
rect 517716 171134 517744 266358
rect 517808 250578 517836 354646
rect 517900 267170 517928 371282
rect 517980 371272 518032 371278
rect 517980 371214 518032 371220
rect 517888 267164 517940 267170
rect 517888 267106 517940 267112
rect 517900 266422 517928 267106
rect 517992 267034 518020 371214
rect 518912 349217 518940 454135
rect 518990 393816 519046 393825
rect 518990 393751 519046 393760
rect 519004 362234 519032 393751
rect 519358 392184 519414 392193
rect 519358 392119 519414 392128
rect 519174 390824 519230 390833
rect 519174 390759 519230 390768
rect 519082 389328 519138 389337
rect 519082 389263 519138 389272
rect 518992 362228 519044 362234
rect 518992 362170 519044 362176
rect 519096 359582 519124 389263
rect 519188 365022 519216 390759
rect 519266 388104 519322 388113
rect 519266 388039 519322 388048
rect 519176 365016 519228 365022
rect 519176 364958 519228 364964
rect 519280 364334 519308 388039
rect 519188 364306 519308 364334
rect 519188 363662 519216 364306
rect 519176 363656 519228 363662
rect 519176 363598 519228 363604
rect 519084 359576 519136 359582
rect 519084 359518 519136 359524
rect 518898 349208 518954 349217
rect 518898 349143 518954 349152
rect 517980 267028 518032 267034
rect 517980 266970 518032 266976
rect 517888 266416 517940 266422
rect 517888 266358 517940 266364
rect 517888 251116 517940 251122
rect 517888 251058 517940 251064
rect 517900 250646 517928 251058
rect 517888 250640 517940 250646
rect 517888 250582 517940 250588
rect 517796 250572 517848 250578
rect 517796 250514 517848 250520
rect 517624 171106 517744 171134
rect 510528 163668 510580 163674
rect 510528 163610 510580 163616
rect 517520 163668 517572 163674
rect 517520 163610 517572 163616
rect 478420 163532 478472 163538
rect 478420 163474 478472 163480
rect 455786 163160 455842 163169
rect 455786 163095 455842 163104
rect 438032 162988 438084 162994
rect 438032 162930 438084 162936
rect 436928 162920 436980 162926
rect 436928 162862 436980 162868
rect 455800 162790 455828 163095
rect 455788 162784 455840 162790
rect 403070 162752 403126 162761
rect 403070 162687 403126 162696
rect 404358 162752 404414 162761
rect 404358 162687 404414 162696
rect 405738 162752 405794 162761
rect 405738 162687 405794 162696
rect 407210 162752 407266 162761
rect 407210 162687 407266 162696
rect 408314 162752 408370 162761
rect 408314 162687 408370 162696
rect 408498 162752 408554 162761
rect 408498 162687 408554 162696
rect 409970 162752 410026 162761
rect 409970 162687 410026 162696
rect 410614 162752 410670 162761
rect 410614 162687 410670 162696
rect 411350 162752 411406 162761
rect 411350 162687 411406 162696
rect 412638 162752 412694 162761
rect 412638 162687 412694 162696
rect 413650 162752 413706 162761
rect 413650 162687 413706 162696
rect 414018 162752 414074 162761
rect 414018 162687 414074 162696
rect 415398 162752 415454 162761
rect 415398 162687 415454 162696
rect 416778 162752 416834 162761
rect 416778 162687 416834 162696
rect 418158 162752 418214 162761
rect 418158 162687 418214 162696
rect 419538 162752 419594 162761
rect 419538 162687 419594 162696
rect 420918 162752 420974 162761
rect 420918 162687 420974 162696
rect 422298 162752 422354 162761
rect 422298 162687 422354 162696
rect 423678 162752 423734 162761
rect 423678 162687 423734 162696
rect 425058 162752 425114 162761
rect 425058 162687 425114 162696
rect 426438 162752 426494 162761
rect 426438 162687 426494 162696
rect 429106 162752 429162 162761
rect 429106 162687 429162 162696
rect 429290 162752 429346 162761
rect 429290 162687 429346 162696
rect 430578 162752 430634 162761
rect 430578 162687 430634 162696
rect 431958 162752 432014 162761
rect 431958 162687 432014 162696
rect 434626 162752 434682 162761
rect 434626 162687 434682 162696
rect 435362 162752 435418 162761
rect 435362 162687 435418 162696
rect 435914 162752 435970 162761
rect 435914 162687 435970 162696
rect 438490 162752 438546 162761
rect 438490 162687 438546 162696
rect 439042 162752 439098 162761
rect 439042 162687 439098 162696
rect 440882 162752 440938 162761
rect 440882 162687 440938 162696
rect 443458 162752 443514 162761
rect 443458 162687 443514 162696
rect 445850 162752 445906 162761
rect 445850 162687 445906 162696
rect 448242 162752 448298 162761
rect 448242 162687 448298 162696
rect 453210 162752 453266 162761
rect 455788 162726 455840 162732
rect 458362 162752 458418 162761
rect 453210 162687 453266 162696
rect 458362 162687 458364 162696
rect 402978 162208 403034 162217
rect 402978 162143 403034 162152
rect 401600 148980 401652 148986
rect 401600 148922 401652 148928
rect 400220 148912 400272 148918
rect 400220 148854 400272 148860
rect 398840 148436 398892 148442
rect 398840 148378 398892 148384
rect 396724 146124 396776 146130
rect 396724 146066 396776 146072
rect 402992 145790 403020 162143
rect 402980 145784 403032 145790
rect 402980 145726 403032 145732
rect 403084 145722 403112 162687
rect 403072 145716 403124 145722
rect 403072 145658 403124 145664
rect 404372 145654 404400 162687
rect 404360 145648 404412 145654
rect 404360 145590 404412 145596
rect 405752 145586 405780 162687
rect 407224 145926 407252 162687
rect 408328 162110 408356 162687
rect 408316 162104 408368 162110
rect 408316 162046 408368 162052
rect 407212 145920 407264 145926
rect 407212 145862 407264 145868
rect 408512 145858 408540 162687
rect 409984 146062 410012 162687
rect 410628 161974 410656 162687
rect 411258 162208 411314 162217
rect 411258 162143 411314 162152
rect 410616 161968 410668 161974
rect 410616 161910 410668 161916
rect 409972 146056 410024 146062
rect 409972 145998 410024 146004
rect 408500 145852 408552 145858
rect 408500 145794 408552 145800
rect 405740 145580 405792 145586
rect 405740 145522 405792 145528
rect 396172 145444 396224 145450
rect 396172 145386 396224 145392
rect 393320 145376 393372 145382
rect 393320 145318 393372 145324
rect 411272 145314 411300 162143
rect 411364 145994 411392 162687
rect 412652 146033 412680 162687
rect 413664 162178 413692 162687
rect 413652 162172 413704 162178
rect 413652 162114 413704 162120
rect 414032 146198 414060 162687
rect 414020 146192 414072 146198
rect 415412 146169 415440 162687
rect 414020 146134 414072 146140
rect 415398 146160 415454 146169
rect 416792 146130 416820 162687
rect 418172 159934 418200 162687
rect 418434 162208 418490 162217
rect 418434 162143 418490 162152
rect 418448 162042 418476 162143
rect 418436 162036 418488 162042
rect 418436 161978 418488 161984
rect 419552 160002 419580 162687
rect 420932 160070 420960 162687
rect 421564 161628 421616 161634
rect 421564 161570 421616 161576
rect 420920 160064 420972 160070
rect 420920 160006 420972 160012
rect 419540 159996 419592 160002
rect 419540 159938 419592 159944
rect 418160 159928 418212 159934
rect 418160 159870 418212 159876
rect 415398 146095 415454 146104
rect 416780 146124 416832 146130
rect 416780 146066 416832 146072
rect 412638 146024 412694 146033
rect 411352 145988 411404 145994
rect 412638 145959 412694 145968
rect 411352 145930 411404 145936
rect 411260 145308 411312 145314
rect 411260 145250 411312 145256
rect 421576 144906 421604 161570
rect 422312 161294 422340 162687
rect 422300 161288 422352 161294
rect 422300 161230 422352 161236
rect 423692 145625 423720 162687
rect 425072 146305 425100 162687
rect 426452 161362 426480 162687
rect 426530 162208 426586 162217
rect 426530 162143 426586 162152
rect 426440 161356 426492 161362
rect 426440 161298 426492 161304
rect 426544 147626 426572 162143
rect 429120 161474 429148 162687
rect 429120 161446 429240 161474
rect 429212 148374 429240 161446
rect 429304 160818 429332 162687
rect 429292 160812 429344 160818
rect 429292 160754 429344 160760
rect 430592 160750 430620 162687
rect 433524 162308 433576 162314
rect 433524 162250 433576 162256
rect 433536 162217 433564 162250
rect 433522 162208 433578 162217
rect 433522 162143 433578 162152
rect 434640 161430 434668 162687
rect 435376 161566 435404 162687
rect 435928 162246 435956 162687
rect 438504 162450 438532 162687
rect 438492 162444 438544 162450
rect 438492 162386 438544 162392
rect 435916 162240 435968 162246
rect 435916 162182 435968 162188
rect 439056 161634 439084 162687
rect 440896 162518 440924 162687
rect 440884 162512 440936 162518
rect 440884 162454 440936 162460
rect 443472 162382 443500 162687
rect 445864 162586 445892 162687
rect 448256 162654 448284 162687
rect 448244 162648 448296 162654
rect 448244 162590 448296 162596
rect 445852 162580 445904 162586
rect 445852 162522 445904 162528
rect 443460 162376 443512 162382
rect 443460 162318 443512 162324
rect 453224 161906 453252 162687
rect 458416 162687 458418 162696
rect 503258 162752 503314 162761
rect 503258 162687 503314 162696
rect 458364 162658 458416 162664
rect 503272 162314 503300 162687
rect 503626 162616 503682 162625
rect 503626 162551 503682 162560
rect 503260 162308 503312 162314
rect 503260 162250 503312 162256
rect 503640 162178 503668 162551
rect 503628 162172 503680 162178
rect 503628 162114 503680 162120
rect 453212 161900 453264 161906
rect 453212 161842 453264 161848
rect 439044 161628 439096 161634
rect 439044 161570 439096 161576
rect 435364 161560 435416 161566
rect 435364 161502 435416 161508
rect 434720 161492 434772 161498
rect 434720 161434 434772 161440
rect 434628 161424 434680 161430
rect 434628 161366 434680 161372
rect 430580 160744 430632 160750
rect 430580 160686 430632 160692
rect 434732 149054 434760 161434
rect 434720 149048 434772 149054
rect 434720 148990 434772 148996
rect 429200 148368 429252 148374
rect 429200 148310 429252 148316
rect 426532 147620 426584 147626
rect 426532 147562 426584 147568
rect 425058 146296 425114 146305
rect 510540 146282 510568 163610
rect 517624 163554 517652 171106
rect 517532 163526 517652 163554
rect 517532 162178 517560 163526
rect 517612 162852 517664 162858
rect 517612 162794 517664 162800
rect 517624 162314 517652 162794
rect 517612 162308 517664 162314
rect 517612 162250 517664 162256
rect 517520 162172 517572 162178
rect 517520 162114 517572 162120
rect 510540 146266 510660 146282
rect 510540 146260 510672 146266
rect 510540 146254 510620 146260
rect 425058 146231 425114 146240
rect 510620 146202 510672 146208
rect 498660 146192 498712 146198
rect 510632 146169 510660 146202
rect 498660 146134 498712 146140
rect 510618 146160 510674 146169
rect 423678 145616 423734 145625
rect 423678 145551 423734 145560
rect 498672 144945 498700 146134
rect 499856 146124 499908 146130
rect 510618 146095 510674 146104
rect 499856 146066 499908 146072
rect 499868 144945 499896 146066
rect 498658 144936 498714 144945
rect 421564 144900 421616 144906
rect 498658 144871 498714 144880
rect 499854 144936 499910 144945
rect 499854 144871 499910 144880
rect 421564 144842 421616 144848
rect 397092 59832 397144 59838
rect 396078 59800 396134 59809
rect 396078 59735 396080 59744
rect 396132 59735 396134 59744
rect 397090 59800 397092 59809
rect 397144 59800 397146 59809
rect 397090 59735 397146 59744
rect 416962 59800 417018 59809
rect 416962 59735 417018 59744
rect 418434 59800 418490 59809
rect 418434 59735 418490 59744
rect 422850 59800 422906 59809
rect 422850 59735 422906 59744
rect 423954 59800 424010 59809
rect 423954 59735 424010 59744
rect 396080 59706 396132 59712
rect 416976 59702 417004 59735
rect 416964 59696 417016 59702
rect 403070 59664 403126 59673
rect 403070 59599 403126 59608
rect 404174 59664 404230 59673
rect 404174 59599 404230 59608
rect 412546 59664 412602 59673
rect 416964 59638 417016 59644
rect 412546 59599 412602 59608
rect 418160 59628 418212 59634
rect 403084 59294 403112 59599
rect 403072 59288 403124 59294
rect 403072 59230 403124 59236
rect 404188 58614 404216 59599
rect 404176 58608 404228 58614
rect 404176 58550 404228 58556
rect 397458 57896 397514 57905
rect 397458 57831 397514 57840
rect 399482 57896 399538 57905
rect 399482 57831 399538 57840
rect 400218 57896 400274 57905
rect 400218 57831 400274 57840
rect 401690 57896 401746 57905
rect 401690 57831 401746 57840
rect 404358 57896 404414 57905
rect 404358 57831 404414 57840
rect 405830 57896 405886 57905
rect 405830 57831 405886 57840
rect 407210 57896 407266 57905
rect 407210 57831 407266 57840
rect 408314 57896 408370 57905
rect 408314 57831 408370 57840
rect 408682 57896 408738 57905
rect 408682 57831 408738 57840
rect 409878 57896 409934 57905
rect 409878 57831 409934 57840
rect 411350 57896 411406 57905
rect 411350 57831 411406 57840
rect 379980 54868 380032 54874
rect 379980 54810 380032 54816
rect 377220 54732 377272 54738
rect 377220 54674 377272 54680
rect 376576 54596 376628 54602
rect 376576 54538 376628 54544
rect 376208 54528 376260 54534
rect 376208 54470 376260 54476
rect 397472 54398 397500 57831
rect 399496 56574 399524 57831
rect 399484 56568 399536 56574
rect 399484 56510 399536 56516
rect 400232 54466 400260 57831
rect 401704 55894 401732 57831
rect 401692 55888 401744 55894
rect 401692 55830 401744 55836
rect 404372 54534 404400 57831
rect 405844 54670 405872 57831
rect 405832 54664 405884 54670
rect 405832 54606 405884 54612
rect 407224 54602 407252 57831
rect 408328 55826 408356 57831
rect 408696 55962 408724 57831
rect 408684 55956 408736 55962
rect 408684 55898 408736 55904
rect 408316 55820 408368 55826
rect 408316 55762 408368 55768
rect 409892 54738 409920 57831
rect 411258 56944 411314 56953
rect 411258 56879 411314 56888
rect 411272 56030 411300 56879
rect 411260 56024 411312 56030
rect 411260 55966 411312 55972
rect 411364 54806 411392 57831
rect 412560 56953 412588 59599
rect 418160 59570 418212 59576
rect 418172 59537 418200 59570
rect 418158 59528 418214 59537
rect 418158 59463 418214 59472
rect 418448 59430 418476 59735
rect 422864 59566 422892 59735
rect 423494 59664 423550 59673
rect 423494 59599 423550 59608
rect 422852 59560 422904 59566
rect 422852 59502 422904 59508
rect 418436 59424 418488 59430
rect 418436 59366 418488 59372
rect 420642 59392 420698 59401
rect 420642 59327 420698 59336
rect 421746 59392 421802 59401
rect 421746 59327 421802 59336
rect 420656 59158 420684 59327
rect 421760 59226 421788 59327
rect 421748 59220 421800 59226
rect 421748 59162 421800 59168
rect 420644 59152 420696 59158
rect 420644 59094 420696 59100
rect 423508 59022 423536 59599
rect 423968 59498 423996 59735
rect 480902 59664 480958 59673
rect 480902 59599 480958 59608
rect 423956 59492 424008 59498
rect 423956 59434 424008 59440
rect 425978 59392 426034 59401
rect 425978 59327 426034 59336
rect 428186 59392 428242 59401
rect 428186 59327 428242 59336
rect 453394 59392 453450 59401
rect 453394 59327 453450 59336
rect 463514 59392 463570 59401
rect 463514 59327 463570 59336
rect 425992 59090 426020 59327
rect 425980 59084 426032 59090
rect 425980 59026 426032 59032
rect 423496 59016 423548 59022
rect 423496 58958 423548 58964
rect 428200 58682 428228 59327
rect 453408 58954 453436 59327
rect 453396 58948 453448 58954
rect 453396 58890 453448 58896
rect 463528 58886 463556 59327
rect 463516 58880 463568 58886
rect 463516 58822 463568 58828
rect 480916 58818 480944 59599
rect 485962 59256 486018 59265
rect 485962 59191 486018 59200
rect 480904 58812 480956 58818
rect 480904 58754 480956 58760
rect 485976 58750 486004 59191
rect 485964 58744 486016 58750
rect 485964 58686 486016 58692
rect 428188 58676 428240 58682
rect 428188 58618 428240 58624
rect 478420 57928 478472 57934
rect 414570 57896 414626 57905
rect 414570 57831 414626 57840
rect 415490 57896 415546 57905
rect 415490 57831 415546 57840
rect 416042 57896 416098 57905
rect 416042 57831 416098 57840
rect 426438 57896 426494 57905
rect 426438 57831 426494 57840
rect 427634 57896 427690 57905
rect 427634 57831 427690 57840
rect 427818 57896 427874 57905
rect 427818 57831 427874 57840
rect 429198 57896 429254 57905
rect 429198 57831 429254 57840
rect 430578 57896 430634 57905
rect 430578 57831 430634 57840
rect 432234 57896 432290 57905
rect 432234 57831 432290 57840
rect 433338 57896 433394 57905
rect 433338 57831 433394 57840
rect 433614 57896 433670 57905
rect 433614 57831 433670 57840
rect 435914 57896 435970 57905
rect 435914 57831 435970 57840
rect 436098 57896 436154 57905
rect 436098 57831 436154 57840
rect 438214 57896 438270 57905
rect 438214 57831 438270 57840
rect 438490 57896 438546 57905
rect 438490 57831 438546 57840
rect 438858 57896 438914 57905
rect 438858 57831 438914 57840
rect 440882 57896 440938 57905
rect 440882 57831 440938 57840
rect 443458 57896 443514 57905
rect 443458 57831 443514 57840
rect 448242 57896 448298 57905
rect 448242 57831 448298 57840
rect 470874 57896 470930 57905
rect 470874 57831 470876 57840
rect 412546 56944 412602 56953
rect 412546 56879 412602 56888
rect 412638 56808 412694 56817
rect 412638 56743 412694 56752
rect 412652 56098 412680 56743
rect 414584 56166 414612 57831
rect 415504 57254 415532 57831
rect 416056 57322 416084 57831
rect 416044 57316 416096 57322
rect 416044 57258 416096 57264
rect 415492 57248 415544 57254
rect 415492 57190 415544 57196
rect 426452 56234 426480 57831
rect 427648 56302 427676 57831
rect 427636 56296 427688 56302
rect 427636 56238 427688 56244
rect 426440 56228 426492 56234
rect 426440 56170 426492 56176
rect 414572 56160 414624 56166
rect 414572 56102 414624 56108
rect 412640 56092 412692 56098
rect 412640 56034 412692 56040
rect 427832 54874 427860 57831
rect 429212 54942 429240 57831
rect 430592 55010 430620 57831
rect 430948 57384 431000 57390
rect 430948 57326 431000 57332
rect 430960 57225 430988 57326
rect 430946 57216 431002 57225
rect 430946 57151 431002 57160
rect 432248 56370 432276 57831
rect 432236 56364 432288 56370
rect 432236 56306 432288 56312
rect 433352 55146 433380 57831
rect 433628 57594 433656 57831
rect 433616 57588 433668 57594
rect 433616 57530 433668 57536
rect 435928 57458 435956 57831
rect 435916 57452 435968 57458
rect 435916 57394 435968 57400
rect 433430 57216 433486 57225
rect 433430 57151 433486 57160
rect 435730 57216 435786 57225
rect 435730 57151 435786 57160
rect 433340 55140 433392 55146
rect 433340 55082 433392 55088
rect 433444 55078 433472 57151
rect 435744 56506 435772 57151
rect 435732 56500 435784 56506
rect 435732 56442 435784 56448
rect 436112 55214 436140 57831
rect 438228 56438 438256 57831
rect 438504 57526 438532 57831
rect 438492 57520 438544 57526
rect 438492 57462 438544 57468
rect 438216 56432 438268 56438
rect 438216 56374 438268 56380
rect 436100 55208 436152 55214
rect 438872 55185 438900 57831
rect 440896 57662 440924 57831
rect 443472 57798 443500 57831
rect 443460 57792 443512 57798
rect 443460 57734 443512 57740
rect 448256 57730 448284 57831
rect 470928 57831 470930 57840
rect 478418 57896 478420 57905
rect 503260 57928 503312 57934
rect 478472 57896 478474 57905
rect 478418 57831 478474 57840
rect 503258 57896 503260 57905
rect 503312 57896 503314 57905
rect 503258 57831 503314 57840
rect 503534 57896 503590 57905
rect 517532 57866 517560 162114
rect 517624 57934 517652 162250
rect 517808 146198 517836 250514
rect 517796 146192 517848 146198
rect 517796 146134 517848 146140
rect 517900 146130 517928 250582
rect 517992 162858 518020 266970
rect 518912 244225 518940 349143
rect 518990 288416 519046 288425
rect 518990 288351 519046 288360
rect 519004 287201 519032 288351
rect 518990 287192 519046 287201
rect 518990 287127 519046 287136
rect 518898 244216 518954 244225
rect 518898 244151 518954 244160
rect 518898 184920 518954 184929
rect 518898 184855 518954 184864
rect 517980 162852 518032 162858
rect 517980 162794 518032 162800
rect 518072 146192 518124 146198
rect 518072 146134 518124 146140
rect 517888 146124 517940 146130
rect 517888 146066 517940 146072
rect 518084 145586 518112 146134
rect 518440 146124 518492 146130
rect 518440 146066 518492 146072
rect 518452 145654 518480 146066
rect 518440 145648 518492 145654
rect 518440 145590 518492 145596
rect 518072 145580 518124 145586
rect 518072 145522 518124 145528
rect 518912 79937 518940 184855
rect 519004 182753 519032 287127
rect 519096 285025 519124 359518
rect 519082 285016 519138 285025
rect 519082 284951 519138 284960
rect 518990 182744 519046 182753
rect 518990 182679 519046 182688
rect 518898 79928 518954 79937
rect 518898 79863 518954 79872
rect 519004 78305 519032 182679
rect 519096 179489 519124 284951
rect 519188 284209 519216 363598
rect 519268 362228 519320 362234
rect 519268 362170 519320 362176
rect 519280 289377 519308 362170
rect 519372 358057 519400 392119
rect 520936 388482 520964 487154
rect 580276 458153 580304 515374
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 580264 454708 580316 454714
rect 580264 454650 580316 454656
rect 580276 404977 580304 454650
rect 580262 404968 580318 404977
rect 580262 404903 580318 404912
rect 520924 388476 520976 388482
rect 520924 388418 520976 388424
rect 580356 388476 580408 388482
rect 580356 388418 580408 388424
rect 580264 371272 580316 371278
rect 580264 371214 580316 371220
rect 519452 365016 519504 365022
rect 519452 364958 519504 364964
rect 519358 358048 519414 358057
rect 519358 357983 519414 357992
rect 519266 289368 519322 289377
rect 519266 289303 519322 289312
rect 519174 284200 519230 284209
rect 519174 284135 519230 284144
rect 519188 282946 519216 284135
rect 519176 282940 519228 282946
rect 519176 282882 519228 282888
rect 519082 179480 519138 179489
rect 519082 179415 519138 179424
rect 519082 178800 519138 178809
rect 519188 178786 519216 282882
rect 519280 184929 519308 289303
rect 519372 288425 519400 357983
rect 519358 288416 519414 288425
rect 519358 288351 519414 288360
rect 519464 285841 519492 364958
rect 580276 325281 580304 371214
rect 580368 351937 580396 388418
rect 580446 378448 580502 378457
rect 580446 378383 580502 378392
rect 580460 371890 580488 378383
rect 580448 371884 580500 371890
rect 580448 371826 580500 371832
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 519450 285832 519506 285841
rect 519450 285767 519506 285776
rect 519358 244216 519414 244225
rect 519358 244151 519414 244160
rect 519266 184920 519322 184929
rect 519266 184855 519322 184864
rect 519268 182164 519320 182170
rect 519268 182106 519320 182112
rect 519280 181393 519308 182106
rect 519266 181384 519322 181393
rect 519266 181319 519322 181328
rect 519138 178758 519216 178786
rect 519082 178735 519138 178744
rect 518990 78296 519046 78305
rect 518990 78231 519046 78240
rect 519096 74225 519124 178735
rect 519280 76809 519308 181319
rect 519372 139369 519400 244151
rect 519464 182170 519492 285767
rect 519910 285016 519966 285025
rect 519910 284951 519966 284960
rect 519924 284374 519952 284951
rect 519912 284368 519964 284374
rect 519912 284310 519964 284316
rect 580264 284368 580316 284374
rect 580264 284310 580316 284316
rect 580276 232393 580304 284310
rect 580356 282940 580408 282946
rect 580356 282882 580408 282888
rect 580368 272241 580396 282882
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 520186 182744 520242 182753
rect 520186 182679 520242 182688
rect 520200 182238 520228 182679
rect 520188 182232 520240 182238
rect 520188 182174 520240 182180
rect 580264 182232 580316 182238
rect 580264 182174 580316 182180
rect 519452 182164 519504 182170
rect 519452 182106 519504 182112
rect 519450 179480 519506 179489
rect 519450 179415 519506 179424
rect 519358 139360 519414 139369
rect 519358 139295 519414 139304
rect 519266 76800 519322 76809
rect 519266 76735 519322 76744
rect 519464 75449 519492 179415
rect 580276 152697 580304 182174
rect 580368 182170 580396 192471
rect 580356 182164 580408 182170
rect 580356 182106 580408 182112
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580264 145648 580316 145654
rect 580264 145590 580316 145596
rect 520188 80028 520240 80034
rect 520188 79970 520240 79976
rect 520200 79937 520228 79970
rect 520186 79928 520242 79937
rect 520186 79863 520242 79872
rect 519450 75440 519506 75449
rect 519450 75375 519506 75384
rect 519082 74216 519138 74225
rect 519082 74151 519138 74160
rect 517612 57928 517664 57934
rect 517612 57870 517664 57876
rect 503534 57831 503536 57840
rect 470876 57802 470928 57808
rect 503588 57831 503590 57840
rect 517520 57860 517572 57866
rect 503536 57802 503588 57808
rect 517520 57802 517572 57808
rect 448244 57724 448296 57730
rect 448244 57666 448296 57672
rect 440884 57656 440936 57662
rect 440884 57598 440936 57604
rect 436100 55150 436152 55156
rect 438858 55176 438914 55185
rect 438858 55111 438914 55120
rect 433432 55072 433484 55078
rect 433432 55014 433484 55020
rect 430580 55004 430632 55010
rect 430580 54946 430632 54952
rect 429200 54936 429252 54942
rect 429200 54878 429252 54884
rect 427820 54868 427872 54874
rect 427820 54810 427872 54816
rect 411352 54800 411404 54806
rect 411352 54742 411404 54748
rect 409880 54732 409932 54738
rect 409880 54674 409932 54680
rect 407212 54596 407264 54602
rect 407212 54538 407264 54544
rect 404360 54528 404412 54534
rect 404360 54470 404412 54476
rect 400220 54460 400272 54466
rect 400220 54402 400272 54408
rect 374736 54392 374788 54398
rect 374736 54334 374788 54340
rect 397460 54392 397512 54398
rect 397460 54334 397512 54340
rect 580276 33153 580304 145590
rect 580356 145580 580408 145586
rect 580356 145522 580408 145528
rect 580368 73001 580396 145522
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580460 80034 580488 112775
rect 580448 80028 580500 80034
rect 580448 79970 580500 79976
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 632032 3570 632088
rect 3422 579944 3478 580000
rect 2962 410488 3018 410544
rect 3330 358400 3386 358456
rect 3054 201864 3110 201920
rect 3606 514800 3662 514856
rect 3606 462576 3662 462632
rect 3514 97552 3570 97608
rect 3422 58520 3478 58576
rect 40682 632032 40738 632088
rect 40590 373224 40646 373280
rect 57702 620608 57758 620664
rect 57518 614352 57574 614408
rect 57426 589872 57482 589928
rect 57334 586336 57390 586392
rect 57058 577632 57114 577688
rect 57150 574912 57206 574968
rect 57334 571512 57390 571568
rect 57242 565392 57298 565448
rect 57610 593408 57666 593464
rect 57518 583616 57574 583672
rect 59266 617752 59322 617808
rect 59082 611632 59138 611688
rect 58898 608232 58954 608288
rect 57886 599528 57942 599584
rect 57886 595992 57942 596048
rect 58530 568792 58586 568848
rect 58806 581032 58862 581088
rect 58990 602112 59046 602168
rect 59174 605512 59230 605568
rect 106370 625232 106426 625288
rect 59542 562732 59598 562788
rect 86958 559544 87014 559600
rect 120814 598304 120870 598360
rect 120998 576816 121054 576872
rect 121458 570968 121514 571024
rect 121090 564848 121146 564904
rect 121182 562128 121238 562184
rect 121734 613808 121790 613864
rect 121826 611088 121882 611144
rect 121918 601568 121974 601624
rect 122194 586608 122250 586664
rect 122102 583208 122158 583264
rect 122010 580488 122066 580544
rect 123022 619928 123078 619984
rect 122930 568248 122986 568304
rect 123114 617208 123170 617264
rect 123574 607688 123630 607744
rect 123206 604968 123262 605024
rect 123390 595448 123446 595504
rect 123298 592728 123354 592784
rect 123482 574368 123538 574424
rect 124126 589348 124182 589384
rect 124126 589328 124128 589348
rect 124128 589328 124180 589348
rect 124180 589328 124182 589348
rect 137374 620608 137430 620664
rect 136730 608232 136786 608288
rect 136638 595992 136694 596048
rect 136914 589872 136970 589928
rect 136730 577632 136786 577688
rect 137282 574912 137338 574968
rect 137190 568792 137246 568848
rect 137650 611632 137706 611688
rect 137466 583752 137522 583808
rect 137558 571512 137614 571568
rect 139030 617752 139086 617808
rect 138570 614352 138626 614408
rect 137926 599528 137982 599584
rect 137926 593408 137982 593464
rect 138478 562672 138534 562728
rect 138938 605512 138994 605568
rect 138846 602112 138902 602168
rect 138754 587152 138810 587208
rect 138662 581032 138718 581088
rect 139306 565392 139362 565448
rect 200762 610544 200818 610600
rect 200854 598304 200910 598360
rect 200946 574096 201002 574152
rect 201038 568248 201094 568304
rect 201130 562128 201186 562184
rect 201590 619928 201646 619984
rect 202970 617208 203026 617264
rect 201866 613808 201922 613864
rect 201774 604968 201830 605024
rect 202878 607688 202934 607744
rect 201958 592728 202014 592784
rect 202234 586608 202290 586664
rect 202050 583208 202106 583264
rect 202142 580488 202198 580544
rect 202326 570968 202382 571024
rect 203062 601568 203118 601624
rect 203154 595448 203210 595504
rect 204166 589348 204222 589384
rect 204166 589328 204168 589348
rect 204168 589328 204220 589348
rect 204220 589328 204222 589348
rect 203246 577088 203302 577144
rect 203338 564848 203394 564904
rect 216678 620608 216734 620664
rect 216678 617752 216734 617808
rect 215942 611632 215998 611688
rect 216678 608232 216734 608288
rect 217230 602112 217286 602168
rect 216678 593428 216734 593464
rect 216678 593408 216680 593428
rect 216680 593408 216732 593428
rect 216732 593408 216734 593428
rect 216678 589872 216734 589928
rect 216678 587152 216734 587208
rect 216034 577632 216090 577688
rect 216678 574912 216734 574968
rect 216678 571512 216734 571568
rect 217138 562672 217194 562728
rect 217690 614352 217746 614408
rect 217414 583752 217470 583808
rect 217782 599528 217838 599584
rect 217690 581032 217746 581088
rect 217598 565392 217654 565448
rect 218702 596128 218758 596184
rect 219254 605512 219310 605568
rect 219162 568792 219218 568848
rect 238666 543088 238722 543144
rect 241518 542680 241574 542736
rect 245842 542952 245898 543008
rect 248694 542816 248750 542872
rect 255134 542408 255190 542464
rect 264426 541048 264482 541104
rect 280894 594904 280950 594960
rect 281630 619928 281686 619984
rect 281170 592728 281226 592784
rect 281538 568248 281594 568304
rect 281262 564848 281318 564904
rect 281538 562128 281594 562184
rect 281722 617208 281778 617264
rect 283010 613808 283066 613864
rect 281998 611088 282054 611144
rect 281814 586608 281870 586664
rect 281906 577088 281962 577144
rect 282918 574368 282974 574424
rect 283654 607688 283710 607744
rect 283102 604968 283158 605024
rect 283194 601568 283250 601624
rect 283286 598848 283342 598904
rect 283562 589348 283618 589384
rect 283562 589328 283564 589348
rect 283564 589328 283616 589348
rect 283616 589328 283618 589348
rect 283378 583208 283434 583264
rect 283470 580488 283526 580544
rect 283562 570968 283618 571024
rect 282918 541592 282974 541648
rect 293130 542544 293186 542600
rect 294510 541184 294566 541240
rect 301594 542816 301650 542872
rect 301594 518744 301650 518800
rect 302238 532344 302294 532400
rect 302882 517384 302938 517440
rect 57702 509924 57758 509960
rect 57702 509904 57704 509924
rect 57704 509904 57756 509924
rect 57756 509904 57758 509924
rect 57886 509904 57942 509960
rect 40866 373904 40922 373960
rect 315302 632168 315358 632224
rect 317786 629584 317842 629640
rect 317970 620064 318026 620120
rect 317970 615576 318026 615632
rect 317878 610544 317934 610600
rect 317970 606056 318026 606112
rect 317602 601024 317658 601080
rect 317602 596400 317658 596456
rect 317418 586508 317420 586528
rect 317420 586508 317472 586528
rect 317472 586508 317474 586528
rect 317418 586472 317474 586508
rect 317970 582528 318026 582584
rect 317878 577224 317934 577280
rect 317970 571784 318026 571840
rect 317050 568248 317106 568304
rect 317418 557640 317474 557696
rect 317970 553444 318026 553480
rect 317970 553424 317972 553444
rect 317972 553424 318024 553444
rect 318024 553424 318026 553444
rect 317510 549072 317566 549128
rect 317970 543804 317972 543824
rect 317972 543804 318024 543824
rect 318024 543804 318026 543824
rect 317970 543768 318026 543804
rect 316866 541592 316922 541648
rect 318154 625232 318210 625288
rect 318798 592728 318854 592784
rect 318338 562264 318394 562320
rect 318062 542952 318118 543008
rect 318246 542544 318302 542600
rect 317234 541184 317290 541240
rect 318062 539280 318118 539336
rect 317602 534928 317658 534984
rect 317602 529760 317658 529816
rect 317602 525408 317658 525464
rect 319626 632304 319682 632360
rect 346398 632032 346454 632088
rect 392122 632304 392178 632360
rect 419170 632168 419226 632224
rect 328090 630808 328146 630864
rect 405370 630672 405426 630728
rect 428370 558184 428426 558240
rect 319534 542408 319590 542464
rect 319350 518472 319406 518528
rect 319902 518336 319958 518392
rect 337658 518336 337714 518392
rect 427818 520240 427874 520296
rect 356242 518472 356298 518528
rect 374458 518608 374514 518664
rect 302974 502424 303030 502480
rect 302882 487464 302938 487520
rect 43902 472640 43958 472696
rect 42614 472504 42670 472560
rect 43442 469784 43498 469840
rect 43534 267008 43590 267064
rect 45282 469920 45338 469976
rect 50066 478352 50122 478408
rect 46018 374992 46074 375048
rect 46478 267552 46534 267608
rect 46754 475496 46810 475552
rect 47398 268540 47400 268560
rect 47400 268540 47452 268560
rect 47452 268540 47454 268560
rect 47398 268504 47454 268540
rect 47306 268404 47308 268424
rect 47308 268404 47360 268424
rect 47360 268404 47362 268424
rect 47306 268368 47362 268404
rect 49514 478080 49570 478136
rect 47858 267144 47914 267200
rect 47858 144744 47914 144800
rect 48686 459584 48742 459640
rect 49054 267416 49110 267472
rect 49514 162560 49570 162616
rect 50710 477672 50766 477728
rect 50434 475632 50490 475688
rect 50710 465840 50766 465896
rect 50618 462848 50674 462904
rect 50894 477536 50950 477592
rect 50894 463256 50950 463312
rect 50618 161880 50674 161936
rect 51446 383560 51502 383616
rect 51354 267316 51356 267336
rect 51356 267316 51408 267336
rect 51408 267316 51410 267336
rect 51354 267280 51410 267316
rect 51630 459584 51686 459640
rect 53562 466112 53618 466168
rect 52366 459584 52422 459640
rect 52826 375264 52882 375320
rect 52366 374856 52422 374912
rect 52366 267280 52422 267336
rect 52734 264832 52790 264888
rect 53378 459584 53434 459640
rect 53194 264832 53250 264888
rect 53470 162424 53526 162480
rect 54298 145696 54354 145752
rect 55954 459584 56010 459640
rect 55678 371320 55734 371376
rect 55126 162696 55182 162752
rect 56322 162288 56378 162344
rect 56966 412256 57022 412312
rect 57058 410352 57114 410408
rect 57058 408584 57114 408640
rect 56966 407360 57022 407416
rect 57058 405748 57114 405784
rect 57058 405728 57060 405748
rect 57060 405728 57112 405748
rect 57112 405728 57114 405748
rect 57058 404388 57114 404424
rect 57058 404368 57060 404388
rect 57060 404368 57112 404388
rect 57112 404368 57114 404388
rect 57058 403028 57114 403064
rect 57058 403008 57060 403028
rect 57060 403008 57112 403028
rect 57112 403008 57114 403028
rect 56598 384956 56600 384976
rect 56600 384956 56652 384976
rect 56652 384956 56654 384976
rect 56598 384920 56654 384956
rect 56598 383016 56654 383072
rect 57242 383288 57298 383344
rect 56874 304952 56930 305008
rect 56874 201320 56930 201376
rect 56874 198736 56930 198792
rect 55954 160112 56010 160168
rect 56414 145560 56470 145616
rect 57150 307672 57206 307728
rect 57150 306856 57206 306912
rect 57518 307672 57574 307728
rect 57334 303592 57390 303648
rect 57242 278704 57298 278760
rect 57058 201864 57114 201920
rect 56966 195200 57022 195256
rect 56874 93744 56930 93800
rect 57150 201320 57206 201376
rect 57058 97416 57114 97472
rect 57518 302232 57574 302288
rect 57426 299512 57482 299568
rect 57426 298152 57482 298208
rect 57334 198736 57390 198792
rect 57334 197376 57390 197432
rect 57150 96464 57206 96520
rect 57702 303592 57758 303648
rect 57610 301280 57666 301336
rect 58990 475904 59046 475960
rect 58438 383560 58494 383616
rect 58530 372816 58586 372872
rect 58622 372680 58678 372736
rect 57886 305904 57942 305960
rect 57886 304952 57942 305008
rect 57886 278704 57942 278760
rect 57518 197376 57574 197432
rect 57702 196016 57758 196072
rect 57518 195200 57574 195256
rect 57426 193160 57482 193216
rect 57334 93336 57390 93392
rect 58530 275984 58586 276040
rect 58714 279928 58770 279984
rect 58806 278024 58862 278080
rect 58622 267008 58678 267064
rect 58346 175208 58402 175264
rect 57886 173304 57942 173360
rect 57702 91024 57758 91080
rect 57518 90480 57574 90536
rect 57426 88168 57482 88224
rect 2778 19352 2834 19408
rect 57886 68856 57942 68912
rect 59082 466384 59138 466440
rect 58990 175208 59046 175264
rect 59174 466248 59230 466304
rect 58622 145832 58678 145888
rect 58530 145696 58586 145752
rect 59910 465976 59966 466032
rect 59818 276120 59874 276176
rect 59818 268776 59874 268832
rect 59818 267144 59874 267200
rect 59818 266328 59874 266384
rect 61474 471144 61530 471200
rect 66350 478624 66406 478680
rect 68650 478760 68706 478816
rect 68926 478760 68982 478816
rect 67822 460128 67878 460184
rect 67730 459992 67786 460048
rect 67638 459040 67694 459096
rect 69202 463120 69258 463176
rect 69110 460400 69166 460456
rect 70490 463392 70546 463448
rect 71778 460808 71834 460864
rect 71962 463256 72018 463312
rect 73802 477944 73858 478000
rect 73342 461488 73398 461544
rect 75826 478624 75882 478680
rect 75918 460672 75974 460728
rect 77758 478488 77814 478544
rect 77298 478352 77354 478408
rect 78678 478624 78734 478680
rect 79506 478760 79562 478816
rect 80150 462984 80206 463040
rect 74722 460536 74778 460592
rect 74630 460264 74686 460320
rect 69018 458904 69074 458960
rect 84290 465840 84346 465896
rect 85762 466112 85818 466168
rect 91374 478216 91430 478272
rect 89810 466384 89866 466440
rect 91282 466248 91338 466304
rect 89902 465704 89958 465760
rect 94042 478080 94098 478136
rect 92662 465976 92718 466032
rect 95790 475904 95846 475960
rect 93858 462848 93914 462904
rect 107750 462848 107806 462904
rect 120078 475496 120134 475552
rect 119158 472640 119214 472696
rect 121366 475768 121422 475824
rect 120906 475632 120962 475688
rect 123574 472504 123630 472560
rect 126610 475360 126666 475416
rect 125874 469920 125930 469976
rect 125782 469784 125838 469840
rect 127070 468424 127126 468480
rect 145102 475360 145158 475416
rect 144734 474136 144790 474192
rect 146022 478080 146078 478136
rect 146482 475496 146538 475552
rect 147310 478352 147366 478408
rect 146942 474272 146998 474328
rect 145562 471280 145618 471336
rect 148230 478216 148286 478272
rect 148690 475632 148746 475688
rect 149978 471552 150034 471608
rect 147678 462984 147734 463040
rect 143538 460264 143594 460320
rect 152646 474000 152702 474056
rect 154854 476856 154910 476912
rect 153934 472504 153990 472560
rect 150530 469784 150586 469840
rect 156050 469920 156106 469976
rect 155958 468560 156014 468616
rect 154670 463120 154726 463176
rect 158810 472776 158866 472832
rect 157430 467064 157486 467120
rect 160282 471416 160338 471472
rect 160190 467200 160246 467256
rect 154578 460400 154634 460456
rect 150438 460128 150494 460184
rect 80242 458768 80298 458824
rect 161662 465976 161718 466032
rect 163594 478488 163650 478544
rect 164514 472640 164570 472696
rect 162858 465840 162914 465896
rect 167182 478624 167238 478680
rect 167090 465704 167146 465760
rect 166998 460672 167054 460728
rect 165618 460536 165674 460592
rect 169850 466112 169906 466168
rect 169942 463392 169998 463448
rect 169758 463256 169814 463312
rect 171230 460808 171286 460864
rect 172886 478760 172942 478816
rect 171322 459312 171378 459368
rect 172610 461488 172666 461544
rect 172518 459176 172574 459232
rect 178314 461352 178370 461408
rect 179970 477944 180026 478000
rect 179602 461624 179658 461680
rect 183558 466248 183614 466304
rect 182822 459992 182878 460048
rect 190918 460964 190974 461000
rect 190918 460944 190920 460964
rect 190920 460944 190972 460964
rect 190972 460944 190974 460964
rect 171138 459040 171194 459096
rect 164238 458904 164294 458960
rect 161478 458768 161534 458824
rect 163410 374584 163466 374640
rect 165986 374604 166042 374640
rect 165986 374584 165988 374604
rect 165988 374584 166040 374604
rect 166040 374584 166042 374604
rect 93582 374448 93638 374504
rect 103518 374448 103574 374504
rect 116030 374448 116086 374504
rect 143538 374448 143594 374504
rect 146206 374448 146262 374504
rect 153474 374448 153530 374504
rect 156510 374448 156566 374504
rect 158534 374468 158590 374504
rect 158534 374448 158536 374468
rect 158536 374448 158588 374468
rect 158588 374448 158590 374468
rect 160926 374448 160982 374504
rect 148966 374196 149022 374232
rect 148966 374176 148968 374196
rect 148968 374176 149020 374196
rect 149020 374176 149022 374196
rect 100850 373668 100852 373688
rect 100852 373668 100904 373688
rect 100904 373668 100906 373688
rect 100850 373632 100906 373668
rect 107842 373632 107898 373688
rect 113546 373632 113602 373688
rect 118330 373652 118386 373688
rect 118330 373632 118332 373652
rect 118332 373632 118384 373652
rect 118384 373632 118386 373652
rect 121366 373632 121422 373688
rect 125782 373632 125838 373688
rect 128910 373652 128966 373688
rect 128910 373632 128912 373652
rect 128912 373632 128964 373652
rect 128964 373632 128966 373652
rect 105450 373496 105506 373552
rect 110418 373516 110474 373552
rect 110418 373496 110420 373516
rect 110420 373496 110472 373516
rect 110472 373496 110474 373516
rect 131026 373668 131028 373688
rect 131028 373668 131080 373688
rect 131080 373668 131082 373688
rect 131026 373632 131082 373668
rect 133694 373632 133750 373688
rect 136454 373632 136510 373688
rect 139214 373632 139270 373688
rect 141606 373632 141662 373688
rect 151726 373632 151782 373688
rect 88338 373360 88394 373416
rect 96066 373360 96122 373416
rect 98274 373380 98330 373416
rect 98274 373360 98276 373380
rect 98276 373360 98328 373380
rect 98328 373360 98330 373380
rect 122930 373360 122986 373416
rect 90178 373108 90234 373144
rect 90178 373088 90180 373108
rect 90180 373088 90232 373108
rect 90232 373088 90234 373108
rect 92386 373088 92442 373144
rect 60738 372816 60794 372872
rect 77206 372544 77262 372600
rect 81990 372544 82046 372600
rect 84750 372564 84806 372600
rect 84750 372544 84752 372564
rect 84752 372544 84804 372564
rect 84804 372544 84806 372564
rect 78494 372408 78550 372464
rect 79966 372408 80022 372464
rect 80150 372408 80206 372464
rect 77022 371864 77078 371920
rect 86774 372544 86830 372600
rect 88062 372544 88118 372600
rect 89350 372544 89406 372600
rect 90730 372544 90786 372600
rect 92202 372544 92258 372600
rect 85486 372408 85542 372464
rect 93582 372544 93638 372600
rect 102046 372544 102102 372600
rect 112902 372544 112958 372600
rect 114466 372544 114522 372600
rect 95238 371592 95294 371648
rect 99286 371592 99342 371648
rect 100482 371592 100538 371648
rect 97722 371456 97778 371512
rect 95238 369688 95294 369744
rect 101126 371456 101182 371512
rect 104622 372136 104678 372192
rect 104622 369552 104678 369608
rect 106094 371592 106150 371648
rect 182822 371592 182878 371648
rect 183466 371592 183522 371648
rect 107566 371320 107622 371376
rect 197358 477980 197360 478000
rect 197360 477980 197412 478000
rect 197412 477980 197414 478000
rect 197358 477944 197414 477980
rect 197450 477808 197506 477864
rect 197266 373360 197322 373416
rect 179142 355272 179198 355328
rect 191470 355308 191472 355328
rect 191472 355308 191524 355328
rect 191524 355308 191526 355328
rect 191470 355272 191526 355308
rect 179694 354748 179750 354784
rect 179694 354728 179696 354748
rect 179696 354728 179748 354748
rect 179748 354728 179750 354748
rect 107566 269864 107622 269920
rect 110970 269864 111026 269920
rect 108302 269728 108358 269784
rect 83094 269592 83150 269648
rect 93582 269592 93638 269648
rect 94502 269592 94558 269648
rect 60922 269048 60978 269104
rect 76010 269048 76066 269104
rect 77114 269048 77170 269104
rect 60738 268912 60794 268968
rect 61014 268776 61070 268832
rect 60922 268640 60978 268696
rect 90730 269048 90786 269104
rect 108670 269592 108726 269648
rect 133418 269728 133474 269784
rect 135902 269728 135958 269784
rect 138478 269728 138534 269784
rect 95882 269048 95938 269104
rect 96066 269048 96122 269104
rect 98458 269048 98514 269104
rect 99378 269048 99434 269104
rect 85394 268096 85450 268152
rect 64878 267280 64934 267336
rect 77298 266872 77354 266928
rect 80058 266892 80114 266928
rect 80058 266872 80060 266892
rect 80060 266872 80112 266892
rect 80112 266872 80114 266892
rect 62118 266328 62174 266384
rect 84198 267688 84254 267744
rect 92386 268096 92442 268152
rect 86958 267688 87014 267744
rect 88338 267144 88394 267200
rect 91098 266600 91154 266656
rect 85578 266328 85634 266384
rect 88338 266328 88394 266384
rect 89718 266328 89774 266384
rect 103518 268096 103574 268152
rect 102690 267724 102692 267744
rect 102692 267724 102744 267744
rect 102744 267724 102746 267744
rect 102690 267688 102746 267724
rect 100758 267144 100814 267200
rect 140870 269592 140926 269648
rect 143538 269592 143594 269648
rect 145930 269592 145986 269648
rect 128358 268096 128414 268152
rect 153566 268096 153622 268152
rect 113270 267960 113326 268016
rect 105266 267688 105322 267744
rect 106370 267688 106426 267744
rect 113178 267688 113234 267744
rect 104898 267164 104954 267200
rect 104898 267144 104900 267164
rect 104900 267144 104952 267164
rect 104952 267144 104954 267164
rect 100758 266464 100814 266520
rect 92478 266328 92534 266384
rect 96618 266328 96674 266384
rect 97998 266328 98054 266384
rect 100850 266328 100906 266384
rect 111798 266328 111854 266384
rect 117134 267724 117136 267744
rect 117136 267724 117188 267744
rect 117188 267724 117190 267744
rect 117134 267688 117190 267724
rect 122838 267708 122894 267744
rect 122838 267688 122840 267708
rect 122840 267688 122892 267708
rect 122892 267688 122894 267708
rect 125598 267552 125654 267608
rect 129738 267688 129794 267744
rect 155958 267688 156014 267744
rect 158534 267708 158590 267744
rect 158534 267688 158536 267708
rect 158536 267688 158588 267708
rect 158588 267688 158590 267708
rect 163502 267688 163558 267744
rect 117318 267416 117374 267472
rect 120078 267436 120134 267472
rect 120078 267416 120080 267436
rect 120080 267416 120132 267436
rect 120132 267416 120134 267436
rect 160926 267416 160982 267472
rect 166170 267436 166226 267472
rect 166170 267416 166172 267436
rect 166172 267416 166224 267436
rect 166224 267416 166226 267436
rect 183466 267416 183522 267472
rect 115938 267300 115994 267336
rect 115938 267280 115940 267300
rect 115940 267280 115992 267300
rect 115992 267280 115994 267300
rect 183282 267280 183338 267336
rect 147678 266328 147734 266384
rect 179326 249872 179382 249928
rect 180246 249872 180302 249928
rect 190918 249872 190974 249928
rect 96066 164736 96122 164792
rect 140870 164736 140926 164792
rect 103518 164600 103574 164656
rect 105910 164600 105966 164656
rect 117042 164600 117098 164656
rect 98458 164192 98514 164248
rect 101034 164192 101090 164248
rect 108210 164192 108266 164248
rect 153382 164600 153438 164656
rect 163318 164600 163374 164656
rect 145930 164192 145986 164248
rect 148506 164192 148562 164248
rect 150898 164192 150954 164248
rect 99378 163104 99434 163160
rect 113546 163104 113602 163160
rect 59358 140800 59414 140856
rect 75918 162696 75974 162752
rect 77298 162696 77354 162752
rect 78678 162696 78734 162752
rect 80058 162696 80114 162752
rect 81438 162696 81494 162752
rect 82818 162696 82874 162752
rect 84198 162696 84254 162752
rect 85578 162696 85634 162752
rect 86958 162696 87014 162752
rect 88430 162696 88486 162752
rect 89810 162696 89866 162752
rect 90730 162696 90786 162752
rect 91190 162696 91246 162752
rect 92478 162696 92534 162752
rect 93674 162696 93730 162752
rect 93858 162696 93914 162752
rect 95238 162696 95294 162752
rect 96894 162696 96950 162752
rect 97998 162696 98054 162752
rect 73802 146240 73858 146296
rect 76010 162152 76066 162208
rect 84290 161472 84346 161528
rect 88338 162152 88394 162208
rect 87602 145968 87658 146024
rect 91098 162152 91154 162208
rect 100758 162696 100814 162752
rect 102138 162696 102194 162752
rect 103518 162696 103574 162752
rect 104898 162696 104954 162752
rect 106278 162696 106334 162752
rect 107658 162696 107714 162752
rect 109038 162696 109094 162752
rect 110418 162696 110474 162752
rect 111798 162696 111854 162752
rect 92478 145832 92534 145888
rect 100850 162152 100906 162208
rect 100850 146240 100906 146296
rect 106370 162152 106426 162208
rect 110970 162188 110972 162208
rect 110972 162188 111024 162208
rect 111024 162188 111026 162208
rect 110970 162152 111026 162188
rect 114466 162696 114522 162752
rect 114742 162696 114798 162752
rect 115938 162696 115994 162752
rect 114650 162016 114706 162072
rect 128358 163104 128414 163160
rect 117318 162696 117374 162752
rect 118330 162696 118386 162752
rect 118698 162696 118754 162752
rect 120722 162696 120778 162752
rect 122838 162696 122894 162752
rect 125874 162696 125930 162752
rect 130842 162732 130844 162752
rect 130844 162732 130896 162752
rect 130896 162732 130898 162752
rect 130842 162696 130898 162732
rect 133418 162696 133474 162752
rect 183466 162696 183522 162752
rect 183190 162424 183246 162480
rect 102138 145696 102194 145752
rect 100758 145560 100814 145616
rect 191746 145424 191802 145480
rect 179050 144880 179106 144936
rect 179694 144880 179750 144936
rect 77114 59744 77170 59800
rect 83094 59744 83150 59800
rect 99470 59744 99526 59800
rect 113546 59744 113602 59800
rect 120906 59744 120962 59800
rect 94502 59608 94558 59664
rect 102782 59608 102838 59664
rect 113270 59608 113326 59664
rect 95882 59336 95938 59392
rect 98090 59336 98146 59392
rect 100758 59336 100814 59392
rect 101770 59336 101826 59392
rect 116950 59608 117006 59664
rect 148506 59200 148562 59256
rect 150898 59200 150954 59256
rect 84198 57976 84254 58032
rect 76010 57840 76066 57896
rect 78218 57840 78274 57896
rect 79506 57840 79562 57896
rect 80058 57840 80114 57896
rect 81806 57840 81862 57896
rect 85394 57840 85450 57896
rect 86498 57840 86554 57896
rect 86958 57840 87014 57896
rect 88338 57840 88394 57896
rect 88706 57840 88762 57896
rect 89718 57840 89774 57896
rect 90730 57840 90786 57896
rect 91190 57840 91246 57896
rect 92110 57840 92166 57896
rect 92478 57840 92534 57896
rect 103794 57840 103850 57896
rect 104990 57840 105046 57896
rect 106370 57840 106426 57896
rect 106738 57840 106794 57896
rect 108026 57840 108082 57896
rect 109222 57840 109278 57896
rect 111154 57840 111210 57896
rect 115754 57840 115810 57896
rect 123482 57840 123538 57896
rect 125874 57840 125930 57896
rect 128358 57840 128414 57896
rect 130842 57840 130898 57896
rect 133418 57840 133474 57896
rect 145562 57860 145618 57896
rect 145562 57840 145564 57860
rect 145564 57840 145616 57860
rect 145616 57840 145618 57860
rect 111798 57568 111854 57624
rect 113178 57568 113234 57624
rect 115938 57568 115994 57624
rect 118698 57568 118754 57624
rect 153290 57840 153346 57896
rect 183282 57860 183338 57896
rect 183282 57840 183284 57860
rect 183284 57840 183336 57860
rect 183336 57840 183338 57860
rect 198646 375264 198702 375320
rect 199014 454688 199070 454744
rect 200762 478524 200764 478544
rect 200764 478524 200816 478544
rect 200816 478524 200818 478544
rect 200762 478488 200818 478524
rect 200486 477536 200542 477592
rect 199198 390768 199254 390824
rect 199474 389000 199530 389056
rect 199658 393760 199714 393816
rect 199842 388456 199898 388512
rect 199474 373904 199530 373960
rect 198738 349560 198794 349616
rect 199014 349560 199070 349616
rect 198830 289720 198886 289776
rect 198738 244160 198794 244216
rect 199474 286320 199530 286376
rect 199014 284824 199070 284880
rect 198922 283056 198978 283112
rect 198830 184320 198886 184376
rect 198738 179424 198794 179480
rect 199750 357992 199806 358048
rect 199658 289720 199714 289776
rect 200026 373224 200082 373280
rect 199750 287680 199806 287736
rect 199566 283056 199622 283112
rect 199198 244160 199254 244216
rect 199106 181328 199162 181384
rect 199014 179424 199070 179480
rect 198830 178608 198886 178664
rect 198738 74840 198794 74896
rect 201406 375264 201462 375320
rect 200762 266736 200818 266792
rect 199382 184320 199438 184376
rect 199290 182688 199346 182744
rect 199198 139168 199254 139224
rect 199382 79328 199438 79384
rect 199290 77696 199346 77752
rect 199106 76336 199162 76392
rect 198830 73616 198886 73672
rect 201590 478352 201646 478408
rect 202234 459312 202290 459368
rect 203246 373224 203302 373280
rect 205638 478488 205694 478544
rect 205638 477672 205694 477728
rect 204902 466112 204958 466168
rect 205086 465976 205142 466032
rect 205546 375264 205602 375320
rect 206466 465840 206522 465896
rect 206926 408584 206982 408640
rect 206834 374584 206890 374640
rect 208398 477944 208454 478000
rect 207202 373768 207258 373824
rect 207754 459176 207810 459232
rect 208306 382336 208362 382392
rect 208122 372272 208178 372328
rect 208950 265512 209006 265568
rect 209686 374584 209742 374640
rect 209594 373496 209650 373552
rect 209502 372136 209558 372192
rect 209594 371864 209650 371920
rect 209594 371592 209650 371648
rect 209502 371456 209558 371512
rect 209410 267552 209466 267608
rect 209226 267416 209282 267472
rect 183466 57740 183468 57760
rect 183468 57740 183520 57760
rect 183520 57740 183522 57760
rect 183466 57704 183522 57740
rect 155958 57568 156014 57624
rect 160098 57568 160154 57624
rect 165618 57568 165674 57624
rect 210238 478216 210294 478272
rect 210054 373360 210110 373416
rect 210514 458904 210570 458960
rect 211342 478660 211344 478680
rect 211344 478660 211396 478680
rect 211396 478660 211398 478680
rect 211342 478624 211398 478660
rect 211066 374584 211122 374640
rect 210698 265104 210754 265160
rect 210974 264968 211030 265024
rect 211158 373632 211214 373688
rect 211434 373632 211490 373688
rect 211710 371728 211766 371784
rect 211526 270544 211582 270600
rect 211618 270408 211674 270464
rect 211894 463256 211950 463312
rect 212722 373088 212778 373144
rect 212078 267280 212134 267336
rect 212078 265784 212134 265840
rect 212170 265512 212226 265568
rect 212078 264968 212134 265024
rect 212630 369688 212686 369744
rect 212446 265648 212502 265704
rect 212446 264968 212502 265024
rect 153290 56208 153346 56264
rect 165618 55120 165674 55176
rect 160098 54984 160154 55040
rect 155958 54848 156014 54904
rect 118698 54712 118754 54768
rect 213090 264968 213146 265024
rect 213366 458768 213422 458824
rect 213826 369144 213882 369200
rect 213734 269048 213790 269104
rect 214930 372000 214986 372056
rect 214838 368328 214894 368384
rect 215850 374312 215906 374368
rect 215206 372408 215262 372464
rect 215390 371184 215446 371240
rect 215114 267008 215170 267064
rect 214562 145832 214618 145888
rect 214654 145696 214710 145752
rect 214930 146240 214986 146296
rect 215850 369552 215906 369608
rect 215574 266328 215630 266384
rect 216402 267144 216458 267200
rect 215850 145560 215906 145616
rect 216954 477536 217010 477592
rect 217414 477536 217470 477592
rect 217782 477536 217838 477592
rect 216770 408720 216826 408776
rect 216678 383288 216734 383344
rect 216862 404948 216864 404968
rect 216864 404948 216916 404968
rect 216916 404948 216918 404968
rect 216862 404912 216918 404948
rect 217322 403144 217378 403200
rect 216954 384956 216956 384976
rect 216956 384956 217008 384976
rect 217008 384956 217010 384976
rect 216954 384920 217010 384956
rect 216862 375264 216918 375320
rect 216770 374992 216826 375048
rect 216586 371320 216642 371376
rect 216586 369144 216642 369200
rect 216494 266872 216550 266928
rect 216494 266328 216550 266384
rect 216402 265104 216458 265160
rect 216494 251096 216550 251152
rect 216678 307672 216734 307728
rect 217046 383016 217102 383072
rect 217138 375264 217194 375320
rect 216862 374856 216918 374912
rect 216770 303728 216826 303784
rect 217046 305904 217102 305960
rect 216954 299920 217010 299976
rect 216862 299376 216918 299432
rect 216678 279928 216734 279984
rect 216678 278316 216734 278352
rect 216678 278296 216680 278316
rect 216680 278296 216732 278316
rect 216732 278296 216734 278316
rect 216862 278024 216918 278080
rect 216678 202816 216734 202872
rect 216678 174936 216734 174992
rect 216678 173304 216734 173360
rect 216862 202816 216918 202872
rect 216862 201864 216918 201920
rect 217782 411848 217838 411904
rect 217690 410896 217746 410952
rect 217598 406000 217654 406056
rect 217230 302776 217286 302832
rect 217046 200912 217102 200968
rect 216862 96872 216918 96928
rect 217046 173032 217102 173088
rect 217874 407768 217930 407824
rect 217782 307672 217838 307728
rect 217782 306856 217838 306912
rect 217690 303728 217746 303784
rect 217506 301008 217562 301064
rect 217414 299920 217470 299976
rect 217230 197784 217286 197840
rect 216954 95920 217010 95976
rect 216678 68312 216734 68368
rect 217598 299376 217654 299432
rect 217598 298152 217654 298208
rect 217506 196016 217562 196072
rect 217414 194928 217470 194984
rect 217230 92792 217286 92848
rect 217690 198736 217746 198792
rect 217690 196016 217746 196072
rect 217598 193160 217654 193216
rect 217414 89936 217470 89992
rect 218702 462984 218758 463040
rect 218334 459720 218390 459776
rect 218242 374176 218298 374232
rect 218150 372272 218206 372328
rect 218334 270408 218390 270464
rect 217966 198736 218022 198792
rect 217690 91024 217746 91080
rect 217506 88168 217562 88224
rect 217874 145968 217930 146024
rect 217966 93744 218022 93800
rect 217966 68312 218022 68368
rect 218886 465704 218942 465760
rect 219254 372680 219310 372736
rect 219622 374040 219678 374096
rect 219898 373088 219954 373144
rect 219530 372000 219586 372056
rect 218978 60560 219034 60616
rect 219622 265920 219678 265976
rect 219254 60560 219310 60616
rect 223118 477536 223174 477592
rect 223578 475496 223634 475552
rect 226154 478216 226210 478272
rect 223670 469784 223726 469840
rect 230110 472776 230166 472832
rect 231490 478352 231546 478408
rect 233238 478488 233294 478544
rect 234066 478216 234122 478272
rect 234526 478080 234582 478136
rect 233698 474000 233754 474056
rect 232778 472640 232834 472696
rect 231858 472504 231914 472560
rect 231030 471144 231086 471200
rect 235906 478760 235962 478816
rect 236274 478624 236330 478680
rect 234618 468424 234674 468480
rect 229098 465704 229154 465760
rect 255686 476720 255742 476776
rect 255318 468560 255374 468616
rect 263690 468696 263746 468752
rect 271142 471280 271198 471336
rect 277490 462984 277546 463040
rect 276110 462848 276166 462904
rect 280250 469920 280306 469976
rect 287242 465840 287298 465896
rect 296718 464344 296774 464400
rect 338302 460964 338358 461000
rect 338302 460944 338304 460964
rect 338304 460944 338356 460964
rect 338356 460944 338358 460964
rect 339774 460980 339776 461000
rect 339776 460980 339828 461000
rect 339828 460980 339830 461000
rect 339774 460944 339830 460980
rect 350998 460964 351054 461000
rect 350998 460944 351000 460964
rect 351000 460944 351052 460964
rect 351052 460944 351054 460964
rect 235998 374448 236054 374504
rect 244278 374448 244334 374504
rect 250074 374448 250130 374504
rect 250718 374448 250774 374504
rect 251270 374448 251326 374504
rect 256054 374448 256110 374504
rect 270498 374448 270554 374504
rect 222014 374176 222070 374232
rect 221922 374040 221978 374096
rect 221830 373632 221886 373688
rect 220818 373224 220874 373280
rect 220726 373108 220782 373144
rect 220726 373088 220728 373108
rect 220728 373088 220780 373108
rect 220780 373088 220782 373108
rect 222014 372136 222070 372192
rect 221922 371864 221978 371920
rect 236458 373360 236514 373416
rect 238114 372544 238170 372600
rect 239310 372544 239366 372600
rect 240414 372544 240470 372600
rect 242898 373360 242954 373416
rect 247130 373088 247186 373144
rect 241702 372544 241758 372600
rect 244278 372544 244334 372600
rect 248418 372544 248474 372600
rect 251178 372544 251234 372600
rect 245658 371728 245714 371784
rect 270222 374040 270278 374096
rect 262770 373768 262826 373824
rect 255410 373496 255466 373552
rect 256698 373496 256754 373552
rect 253938 373108 253994 373144
rect 253938 373088 253940 373108
rect 253940 373088 253992 373108
rect 253992 373088 253994 373108
rect 260010 373380 260066 373416
rect 260010 373360 260012 373380
rect 260012 373360 260064 373380
rect 260064 373360 260066 373380
rect 258078 373088 258134 373144
rect 261298 373088 261354 373144
rect 252558 372680 252614 372736
rect 259458 372544 259514 372600
rect 262218 372544 262274 372600
rect 269210 373360 269266 373416
rect 264978 373088 265034 373144
rect 266358 372580 266360 372600
rect 266360 372580 266412 372600
rect 266412 372580 266414 372600
rect 266358 372544 266414 372580
rect 262862 372272 262918 372328
rect 271878 372564 271934 372600
rect 271878 372544 271880 372564
rect 271880 372544 271932 372564
rect 271932 372544 271934 372564
rect 300858 373088 300914 373144
rect 278686 372408 278742 372464
rect 276938 372272 276994 372328
rect 270498 372136 270554 372192
rect 270222 371864 270278 371920
rect 273442 371728 273498 371784
rect 262770 371592 262826 371648
rect 247038 371320 247094 371376
rect 252558 371320 252614 371376
rect 258170 371320 258226 371376
rect 260838 371320 260894 371376
rect 263598 371320 263654 371376
rect 264978 371320 265034 371376
rect 266358 371320 266414 371376
rect 267738 371320 267794 371376
rect 270498 371320 270554 371376
rect 273258 371320 273314 371376
rect 276018 371456 276074 371512
rect 277674 371456 277730 371512
rect 276018 371320 276074 371376
rect 280158 371320 280214 371376
rect 282918 371320 282974 371376
rect 285678 371320 285734 371376
rect 287334 371320 287390 371376
rect 289818 371320 289874 371376
rect 292578 371320 292634 371376
rect 295338 371320 295394 371376
rect 298098 371320 298154 371376
rect 310518 372544 310574 372600
rect 320914 374468 320970 374504
rect 320914 374448 320916 374468
rect 320916 374448 320968 374468
rect 320968 374448 320970 374468
rect 314658 372564 314714 372600
rect 314658 372544 314660 372564
rect 314660 372544 314712 372564
rect 314712 372544 314714 372564
rect 322938 372544 322994 372600
rect 313278 372428 313334 372464
rect 313278 372408 313280 372428
rect 313280 372408 313332 372428
rect 313332 372408 313334 372428
rect 304998 372272 305054 372328
rect 317418 371728 317474 371784
rect 302238 371320 302294 371376
rect 307758 371320 307814 371376
rect 326158 371320 326214 371376
rect 342902 371320 342958 371376
rect 343362 371340 343418 371376
rect 343362 371320 343364 371340
rect 343364 371320 343416 371340
rect 343416 371320 343418 371340
rect 266358 368328 266414 368384
rect 338486 355000 338542 355056
rect 351734 355000 351790 355056
rect 339774 354748 339830 354784
rect 339774 354728 339776 354748
rect 339776 354728 339828 354748
rect 339828 354728 339830 354748
rect 221002 353368 221058 353424
rect 250718 269864 250774 269920
rect 263506 269864 263562 269920
rect 275742 269728 275798 269784
rect 280894 269728 280950 269784
rect 315854 269728 315910 269784
rect 279146 269592 279202 269648
rect 283470 269592 283526 269648
rect 285954 269592 286010 269648
rect 288254 269592 288310 269648
rect 293406 269592 293462 269648
rect 308494 269592 308550 269648
rect 290922 268912 290978 268968
rect 243082 268776 243138 268832
rect 258078 268776 258134 268832
rect 261666 268776 261722 268832
rect 220726 265956 220728 265976
rect 220728 265956 220780 265976
rect 220780 265956 220782 265976
rect 220726 265920 220782 265956
rect 298466 269048 298522 269104
rect 300858 269048 300914 269104
rect 295890 268912 295946 268968
rect 318430 269592 318486 269648
rect 265162 268096 265218 268152
rect 272154 268096 272210 268152
rect 255778 267688 255834 267744
rect 260838 267688 260894 267744
rect 263598 267688 263654 267744
rect 258262 267144 258318 267200
rect 255318 267008 255374 267064
rect 247038 266872 247094 266928
rect 252558 266892 252614 266928
rect 252558 266872 252560 266892
rect 252560 266872 252612 266892
rect 252612 266872 252614 266892
rect 263598 266872 263654 266928
rect 244370 266464 244426 266520
rect 251270 266464 251326 266520
rect 259550 266464 259606 266520
rect 244278 266328 244334 266384
rect 245658 266328 245714 266384
rect 247038 266328 247094 266384
rect 248510 266328 248566 266384
rect 249798 266328 249854 266384
rect 251178 266328 251234 266384
rect 252558 266328 252614 266384
rect 253938 266328 253994 266384
rect 256698 266328 256754 266384
rect 259458 266328 259514 266384
rect 262218 266348 262274 266384
rect 262218 266328 262220 266348
rect 262220 266328 262272 266348
rect 262272 266328 262274 266348
rect 265806 267688 265862 267744
rect 267094 267688 267150 267744
rect 268198 267688 268254 267744
rect 270866 267688 270922 267744
rect 269762 267144 269818 267200
rect 271234 267144 271290 267200
rect 267738 266872 267794 266928
rect 273258 267688 273314 267744
rect 276018 267688 276074 267744
rect 302238 267688 302294 267744
rect 343454 267416 343510 267472
rect 343546 267280 343602 267336
rect 277122 267144 277178 267200
rect 278134 267164 278190 267200
rect 278134 267144 278136 267164
rect 278136 267144 278188 267164
rect 278188 267144 278190 267164
rect 273258 267028 273314 267064
rect 273258 267008 273260 267028
rect 273260 267008 273312 267028
rect 273312 267008 273314 267028
rect 310518 266872 310574 266928
rect 279974 266328 280030 266384
rect 338486 249872 338542 249928
rect 340234 249872 340290 249928
rect 350998 249872 351054 249928
rect 258446 164736 258502 164792
rect 282182 164736 282238 164792
rect 249154 164464 249210 164520
rect 261022 164600 261078 164656
rect 276110 164600 276166 164656
rect 249154 164192 249210 164248
rect 262862 164464 262918 164520
rect 262862 164192 262918 164248
rect 235998 163104 236054 163160
rect 264978 163104 265034 163160
rect 236090 162696 236146 162752
rect 237378 162696 237434 162752
rect 240138 162696 240194 162752
rect 241518 162696 241574 162752
rect 242898 162696 242954 162752
rect 244278 162696 244334 162752
rect 245658 162696 245714 162752
rect 247130 162696 247186 162752
rect 247866 162696 247922 162752
rect 248418 162696 248474 162752
rect 249798 162696 249854 162752
rect 251270 162696 251326 162752
rect 252558 162696 252614 162752
rect 253938 162696 253994 162752
rect 255410 162696 255466 162752
rect 255962 162696 256018 162752
rect 256698 162696 256754 162752
rect 259550 162696 259606 162752
rect 260838 162696 260894 162752
rect 262218 162696 262274 162752
rect 263598 162696 263654 162752
rect 238758 161472 238814 161528
rect 237378 145832 237434 145888
rect 244370 162152 244426 162208
rect 251178 162424 251234 162480
rect 259458 162560 259514 162616
rect 258078 162152 258134 162208
rect 263690 162560 263746 162616
rect 265438 162696 265494 162752
rect 266358 162696 266414 162752
rect 267554 162696 267610 162752
rect 267738 162696 267794 162752
rect 269118 162696 269174 162752
rect 270498 162696 270554 162752
rect 271878 162696 271934 162752
rect 273258 162696 273314 162752
rect 276018 162696 276074 162752
rect 268290 162560 268346 162616
rect 269118 146240 269174 146296
rect 270498 145696 270554 145752
rect 274546 162560 274602 162616
rect 273442 162288 273498 162344
rect 305918 164600 305974 164656
rect 318430 164600 318486 164656
rect 282182 164192 282238 164248
rect 298466 164192 298522 164248
rect 300858 164192 300914 164248
rect 278410 162696 278466 162752
rect 280066 162696 280122 162752
rect 280802 162696 280858 162752
rect 283746 162696 283802 162752
rect 285954 162696 286010 162752
rect 293314 162696 293370 162752
rect 303434 162716 303490 162752
rect 303434 162696 303436 162716
rect 303436 162696 303488 162716
rect 303488 162696 303490 162716
rect 278042 161472 278098 161528
rect 278226 148960 278282 149016
rect 278226 148280 278282 148336
rect 276018 146376 276074 146432
rect 308586 162732 308588 162752
rect 308588 162732 308640 162752
rect 308640 162732 308642 162752
rect 308586 162696 308642 162732
rect 343454 162696 343510 162752
rect 320914 162560 320970 162616
rect 343362 162560 343418 162616
rect 356794 269048 356850 269104
rect 271878 145560 271934 145616
rect 338486 144880 338542 144936
rect 340234 144880 340290 144936
rect 351642 144880 351698 144936
rect 237102 59764 237158 59800
rect 237102 59744 237104 59764
rect 237104 59744 237156 59764
rect 237156 59744 237158 59764
rect 255870 59744 255926 59800
rect 259458 59744 259514 59800
rect 260654 59744 260710 59800
rect 261758 59744 261814 59800
rect 263874 59744 263930 59800
rect 256974 59608 257030 59664
rect 258078 59608 258134 59664
rect 262770 59472 262826 59528
rect 265254 59608 265310 59664
rect 315854 59608 315910 59664
rect 295890 59200 295946 59256
rect 298466 59200 298522 59256
rect 303434 59200 303490 59256
rect 323306 59200 323362 59256
rect 325882 58112 325938 58168
rect 235998 57840 236054 57896
rect 237378 57840 237434 57896
rect 239218 57840 239274 57896
rect 242898 57840 242954 57896
rect 244370 57840 244426 57896
rect 246394 57840 246450 57896
rect 248602 57840 248658 57896
rect 251178 57840 251234 57896
rect 253386 57840 253442 57896
rect 265346 57840 265402 57896
rect 266358 57840 266414 57896
rect 267002 57840 267058 57896
rect 269762 57840 269818 57896
rect 272154 57840 272210 57896
rect 273626 57840 273682 57896
rect 274638 57840 274694 57896
rect 279054 57840 279110 57896
rect 283654 57840 283710 57896
rect 287610 57840 287666 57896
rect 293314 57840 293370 57896
rect 300858 57840 300914 57896
rect 305826 57840 305882 57896
rect 310978 57840 311034 57896
rect 313370 57840 313426 57896
rect 318338 57860 318394 57896
rect 318338 57840 318340 57860
rect 318340 57840 318392 57860
rect 318392 57840 318394 57860
rect 240138 57432 240194 57488
rect 241518 57432 241574 57488
rect 239862 57296 239918 57352
rect 239862 56888 239918 56944
rect 244278 57432 244334 57488
rect 247038 57432 247094 57488
rect 249798 57432 249854 57488
rect 251362 57432 251418 57488
rect 249798 54848 249854 54904
rect 253938 57432 253994 57488
rect 267738 57568 267794 57624
rect 270498 57568 270554 57624
rect 273350 57568 273406 57624
rect 277398 57568 277454 57624
rect 320914 57840 320970 57896
rect 343178 57876 343180 57896
rect 343180 57876 343232 57896
rect 343232 57876 343234 57896
rect 343178 57840 343234 57876
rect 343454 57860 343510 57896
rect 343454 57840 343456 57860
rect 343456 57840 343508 57860
rect 343508 57840 343510 57860
rect 307758 57568 307814 57624
rect 356794 148960 356850 149016
rect 358910 454688 358966 454744
rect 359002 393760 359058 393816
rect 359094 392128 359150 392184
rect 359186 389272 359242 389328
rect 359738 390768 359794 390824
rect 359830 388048 359886 388104
rect 358910 349560 358966 349616
rect 358910 288360 358966 288416
rect 358910 287680 358966 287736
rect 358818 243752 358874 243808
rect 359002 286320 359058 286376
rect 359278 357992 359334 358048
rect 359186 289720 359242 289776
rect 359278 288360 359334 288416
rect 359554 289720 359610 289776
rect 359462 284824 359518 284880
rect 359094 283056 359150 283112
rect 359370 283056 359426 283112
rect 359002 184864 359058 184920
rect 358910 182688 358966 182744
rect 358910 179424 358966 179480
rect 358818 78240 358874 78296
rect 359278 243752 359334 243808
rect 359186 181328 359242 181384
rect 359094 178064 359150 178120
rect 359002 79872 359058 79928
rect 358910 75384 358966 75440
rect 359554 184864 359610 184920
rect 359462 179424 359518 179480
rect 359370 178064 359426 178120
rect 359278 139304 359334 139360
rect 359186 76880 359242 76936
rect 359094 74024 359150 74080
rect 361486 408584 361542 408640
rect 364246 372680 364302 372736
rect 365350 164056 365406 164112
rect 371146 372680 371202 372736
rect 370778 163920 370834 163976
rect 371238 372272 371294 372328
rect 371790 265240 371846 265296
rect 307758 55120 307814 55176
rect 277398 54984 277454 55040
rect 372434 144064 372490 144120
rect 373538 266872 373594 266928
rect 373906 269320 373962 269376
rect 374182 267416 374238 267472
rect 374366 266328 374422 266384
rect 373906 146240 373962 146296
rect 374734 162424 374790 162480
rect 375194 267144 375250 267200
rect 375194 266328 375250 266384
rect 375378 265104 375434 265160
rect 375470 264968 375526 265024
rect 375470 158752 375526 158808
rect 375838 265104 375894 265160
rect 375930 264968 375986 265024
rect 375930 145560 375986 145616
rect 376206 162560 376262 162616
rect 377034 408720 377090 408776
rect 376942 407788 376998 407824
rect 376942 407768 376944 407788
rect 376944 407768 376996 407788
rect 376996 407768 376998 407788
rect 376666 383288 376722 383344
rect 376666 373224 376722 373280
rect 376942 384956 376944 384976
rect 376944 384956 376996 384976
rect 376996 384956 376998 384976
rect 376942 384920 376998 384956
rect 376942 383016 376998 383072
rect 377586 411848 377642 411904
rect 377494 410896 377550 410952
rect 377310 408720 377366 408776
rect 377218 406000 377274 406056
rect 376942 368464 376998 368520
rect 376850 307672 376906 307728
rect 376850 306856 376906 306912
rect 376758 302776 376814 302832
rect 376758 301008 376814 301064
rect 376482 265240 376538 265296
rect 376942 304952 376998 305008
rect 376850 202816 376906 202872
rect 377310 404948 377312 404968
rect 377312 404948 377364 404968
rect 377364 404948 377366 404968
rect 377310 404912 377366 404948
rect 377218 303728 377274 303784
rect 377034 279928 377090 279984
rect 377034 278024 377090 278080
rect 376942 200912 376998 200968
rect 376758 196016 376814 196072
rect 376850 174936 376906 174992
rect 376850 173304 376906 173360
rect 376758 173032 376814 173088
rect 376482 146240 376538 146296
rect 376482 145560 376538 145616
rect 377402 371864 377458 371920
rect 377678 406000 377734 406056
rect 377586 307672 377642 307728
rect 377494 305904 377550 305960
rect 377494 304952 377550 305008
rect 377586 302776 377642 302832
rect 377310 299920 377366 299976
rect 377218 198736 377274 198792
rect 377402 278316 377458 278352
rect 377402 278296 377404 278316
rect 377404 278296 377456 278316
rect 377456 278296 377458 278316
rect 377494 202816 377550 202872
rect 377494 201864 377550 201920
rect 377310 194928 377366 194984
rect 376942 95920 376998 95976
rect 376942 69944 376998 70000
rect 376942 68332 376998 68368
rect 376942 68312 376944 68332
rect 376944 68312 376996 68332
rect 376996 68312 376998 68332
rect 430946 626456 431002 626512
rect 430854 621968 430910 622024
rect 456798 618976 456854 619032
rect 430762 616800 430818 616856
rect 430670 612448 430726 612504
rect 456798 610816 456854 610872
rect 430578 607144 430634 607200
rect 580170 683848 580226 683904
rect 457442 602656 457498 602712
rect 431222 601704 431278 601760
rect 429474 587968 429530 588024
rect 429382 582664 429438 582720
rect 429290 530236 429346 530292
rect 391938 485016 391994 485072
rect 430670 578312 430726 578368
rect 429566 549344 429622 549400
rect 430578 539552 430634 539608
rect 430578 524864 430634 524920
rect 430762 572736 430818 572792
rect 430670 520104 430726 520160
rect 430854 567704 430910 567760
rect 430946 563080 431002 563136
rect 431038 553424 431094 553480
rect 431130 543904 431186 543960
rect 457442 594496 457498 594552
rect 431314 534384 431370 534440
rect 457534 586336 457590 586392
rect 457626 578176 457682 578232
rect 510618 615576 510674 615632
rect 580170 630828 580226 630864
rect 580170 630808 580172 630828
rect 580172 630808 580224 630828
rect 580224 630808 580226 630828
rect 511998 607416 512054 607472
rect 511998 599256 512054 599312
rect 511262 582936 511318 582992
rect 377770 403144 377826 403200
rect 377678 301008 377734 301064
rect 377770 298152 377826 298208
rect 377586 197784 377642 197840
rect 377494 96872 377550 96928
rect 377862 198736 377918 198792
rect 377770 196016 377826 196072
rect 377678 193160 377734 193216
rect 377586 92792 377642 92848
rect 377310 89936 377366 89992
rect 378506 270408 378562 270464
rect 378046 263492 378102 263528
rect 378046 263472 378048 263492
rect 378048 263472 378100 263492
rect 378100 263472 378102 263492
rect 378414 164192 378470 164248
rect 378046 158752 378102 158808
rect 377954 144064 378010 144120
rect 377954 143656 378010 143712
rect 377862 93744 377918 93800
rect 377770 91024 377826 91080
rect 377678 88168 377734 88224
rect 377310 68040 377366 68096
rect 378966 267552 379022 267608
rect 378966 265512 379022 265568
rect 378874 161880 378930 161936
rect 379242 270272 379298 270328
rect 379058 162288 379114 162344
rect 378874 145968 378930 146024
rect 512090 591096 512146 591152
rect 580170 577632 580226 577688
rect 512182 574776 512238 574832
rect 511262 462168 511318 462224
rect 498382 460964 498438 461000
rect 498382 460944 498384 460964
rect 498384 460944 498436 460964
rect 498436 460944 498438 460964
rect 499854 460980 499856 461000
rect 499856 460980 499908 461000
rect 499908 460980 499910 461000
rect 499854 460944 499910 460980
rect 516598 454688 516654 454744
rect 405922 374992 405978 375048
rect 407762 374992 407818 375048
rect 425058 374992 425114 375048
rect 440330 374992 440386 375048
rect 443090 374992 443146 375048
rect 452842 374992 452898 375048
rect 410706 374584 410762 374640
rect 433614 374448 433670 374504
rect 436006 374448 436062 374504
rect 438490 374448 438546 374504
rect 416042 374040 416098 374096
rect 418250 373632 418306 373688
rect 423034 373668 423036 373688
rect 423036 373668 423088 373688
rect 423088 373668 423090 373688
rect 423034 373632 423090 373668
rect 426898 373652 426954 373688
rect 426898 373632 426900 373652
rect 426900 373632 426952 373652
rect 426952 373632 426954 373652
rect 445850 373632 445906 373688
rect 450266 373516 450322 373552
rect 450266 373496 450268 373516
rect 450268 373496 450320 373516
rect 450320 373496 450322 373516
rect 455418 373496 455474 373552
rect 447690 373380 447746 373416
rect 447690 373360 447692 373380
rect 447692 373360 447744 373380
rect 447744 373360 447746 373380
rect 462778 373360 462834 373416
rect 400218 372544 400274 372600
rect 402886 372580 402888 372600
rect 402888 372580 402940 372600
rect 402940 372580 402942 372600
rect 402886 372544 402942 372580
rect 470598 372272 470654 372328
rect 396078 372156 396134 372192
rect 396078 372136 396080 372156
rect 396080 372136 396132 372156
rect 396132 372136 396134 372156
rect 397458 372020 397514 372056
rect 397458 372000 397460 372020
rect 397460 372000 397512 372020
rect 397512 372000 397514 372020
rect 404358 372000 404414 372056
rect 407118 372000 407174 372056
rect 422298 372000 422354 372056
rect 401598 371748 401654 371784
rect 401598 371728 401600 371748
rect 401600 371728 401652 371748
rect 401652 371728 401654 371748
rect 409878 371728 409934 371784
rect 398838 371612 398894 371648
rect 398838 371592 398840 371612
rect 398840 371592 398892 371612
rect 398892 371592 398894 371612
rect 411258 371592 411314 371648
rect 465078 371592 465134 371648
rect 411350 371476 411406 371512
rect 411350 371456 411352 371476
rect 411352 371456 411404 371476
rect 411404 371456 411406 371476
rect 418250 371456 418306 371512
rect 421010 371456 421066 371512
rect 423678 371456 423734 371512
rect 426438 371456 426494 371512
rect 430670 371456 430726 371512
rect 396078 371320 396134 371376
rect 402978 371320 403034 371376
rect 412638 371320 412694 371376
rect 413190 371320 413246 371376
rect 414018 371320 414074 371376
rect 415398 371320 415454 371376
rect 416778 371320 416834 371376
rect 418158 371320 418214 371376
rect 419538 371320 419594 371376
rect 420918 371320 420974 371376
rect 425058 371320 425114 371376
rect 427818 371320 427874 371376
rect 429198 371320 429254 371376
rect 430578 371320 430634 371376
rect 431958 371320 432014 371376
rect 433338 371320 433394 371376
rect 434718 371320 434774 371376
rect 436098 371320 436154 371376
rect 458178 371320 458234 371376
rect 503166 372136 503222 372192
rect 503534 372136 503590 372192
rect 483018 371864 483074 371920
rect 473358 371320 473414 371376
rect 474738 371320 474794 371376
rect 477498 371320 477554 371376
rect 480258 371320 480314 371376
rect 498842 355000 498898 355056
rect 500866 354864 500922 354920
rect 510894 354748 510950 354784
rect 510894 354728 510896 354748
rect 510896 354728 510948 354748
rect 510948 354728 510950 354748
rect 418434 269728 418490 269784
rect 425242 269728 425298 269784
rect 423494 269592 423550 269648
rect 426438 269592 426494 269648
rect 433614 269592 433670 269648
rect 453394 269592 453450 269648
rect 468482 269592 468538 269648
rect 480902 269592 480958 269648
rect 430946 268912 431002 268968
rect 433338 268912 433394 268968
rect 475842 268912 475898 268968
rect 478418 268912 478474 268968
rect 415858 268776 415914 268832
rect 421010 268796 421066 268832
rect 421010 268776 421012 268796
rect 421012 268776 421064 268796
rect 421064 268776 421066 268796
rect 398194 268096 398250 268152
rect 401690 268096 401746 268152
rect 379978 267008 380034 267064
rect 388166 265240 388222 265296
rect 389178 265104 389234 265160
rect 390558 264968 390614 265024
rect 398838 266328 398894 266384
rect 400218 266328 400274 266384
rect 416042 268096 416098 268152
rect 402978 267688 403034 267744
rect 414386 267688 414442 267744
rect 434258 268096 434314 268152
rect 455786 268096 455842 268152
rect 407118 267008 407174 267064
rect 409878 267028 409934 267064
rect 409878 267008 409880 267028
rect 409880 267008 409932 267028
rect 409932 267008 409934 267028
rect 412914 267008 412970 267064
rect 411350 266464 411406 266520
rect 418250 266464 418306 266520
rect 403162 266348 403218 266384
rect 403162 266328 403164 266348
rect 403164 266328 403216 266348
rect 403216 266328 403218 266348
rect 404358 266328 404414 266384
rect 405738 266328 405794 266384
rect 407118 266328 407174 266384
rect 408498 266328 408554 266384
rect 409878 266328 409934 266384
rect 411258 266328 411314 266384
rect 412914 266328 412970 266384
rect 416778 266328 416834 266384
rect 418158 266328 418214 266384
rect 419538 266328 419594 266384
rect 420918 266328 420974 266384
rect 432142 267688 432198 267744
rect 422574 267008 422630 267064
rect 435730 267688 435786 267744
rect 435914 267688 435970 267744
rect 445758 267688 445814 267744
rect 447138 267688 447194 267744
rect 449898 267688 449954 267744
rect 483386 268912 483442 268968
rect 458178 267708 458234 267744
rect 458178 267688 458180 267708
rect 458180 267688 458232 267708
rect 458232 267688 458234 267708
rect 473358 267688 473414 267744
rect 503534 267416 503590 267472
rect 437478 267300 437534 267336
rect 437478 267280 437480 267300
rect 437480 267280 437532 267300
rect 437532 267280 437534 267300
rect 442998 267280 443054 267336
rect 503442 267280 503498 267336
rect 440238 267164 440294 267200
rect 440238 267144 440240 267164
rect 440240 267144 440292 267164
rect 440292 267144 440294 267164
rect 429106 266328 429162 266384
rect 430486 266328 430542 266384
rect 430670 266328 430726 266384
rect 436098 266328 436154 266384
rect 437478 266328 437534 266384
rect 438858 266328 438914 266384
rect 499026 249872 499082 249928
rect 500406 249872 500462 249928
rect 510894 249892 510950 249928
rect 580170 511264 580226 511320
rect 518898 454144 518954 454200
rect 510894 249872 510896 249892
rect 510896 249872 510948 249892
rect 510948 249872 510950 249892
rect 425978 164736 426034 164792
rect 434350 164736 434406 164792
rect 451002 164736 451058 164792
rect 423494 164600 423550 164656
rect 416042 164192 416098 164248
rect 421010 164192 421066 164248
rect 379702 146104 379758 146160
rect 436926 164600 436982 164656
rect 438030 164600 438086 164656
rect 428186 164192 428242 164248
rect 430946 164192 431002 164248
rect 396078 162696 396134 162752
rect 396170 162152 396226 162208
rect 401598 163104 401654 163160
rect 397458 162696 397514 162752
rect 398838 162696 398894 162752
rect 400218 162696 400274 162752
rect 418158 162852 418214 162888
rect 418158 162832 418160 162852
rect 418160 162832 418212 162852
rect 418212 162832 418214 162852
rect 480902 164600 480958 164656
rect 473450 164192 473506 164248
rect 475842 164192 475898 164248
rect 478418 164192 478474 164248
rect 470598 163784 470654 163840
rect 518990 393760 519046 393816
rect 519358 392128 519414 392184
rect 519174 390768 519230 390824
rect 519082 389272 519138 389328
rect 519266 388048 519322 388104
rect 518898 349152 518954 349208
rect 455786 163104 455842 163160
rect 403070 162696 403126 162752
rect 404358 162696 404414 162752
rect 405738 162696 405794 162752
rect 407210 162696 407266 162752
rect 408314 162696 408370 162752
rect 408498 162696 408554 162752
rect 409970 162696 410026 162752
rect 410614 162696 410670 162752
rect 411350 162696 411406 162752
rect 412638 162696 412694 162752
rect 413650 162696 413706 162752
rect 414018 162696 414074 162752
rect 415398 162696 415454 162752
rect 416778 162696 416834 162752
rect 418158 162696 418214 162752
rect 419538 162696 419594 162752
rect 420918 162696 420974 162752
rect 422298 162696 422354 162752
rect 423678 162696 423734 162752
rect 425058 162696 425114 162752
rect 426438 162696 426494 162752
rect 429106 162696 429162 162752
rect 429290 162696 429346 162752
rect 430578 162696 430634 162752
rect 431958 162696 432014 162752
rect 434626 162696 434682 162752
rect 435362 162696 435418 162752
rect 435914 162696 435970 162752
rect 438490 162696 438546 162752
rect 439042 162696 439098 162752
rect 440882 162696 440938 162752
rect 443458 162696 443514 162752
rect 445850 162696 445906 162752
rect 448242 162696 448298 162752
rect 453210 162696 453266 162752
rect 458362 162716 458418 162752
rect 458362 162696 458364 162716
rect 458364 162696 458416 162716
rect 458416 162696 458418 162716
rect 402978 162152 403034 162208
rect 411258 162152 411314 162208
rect 415398 146104 415454 146160
rect 418434 162152 418490 162208
rect 412638 145968 412694 146024
rect 426530 162152 426586 162208
rect 433522 162152 433578 162208
rect 503258 162696 503314 162752
rect 503626 162560 503682 162616
rect 425058 146240 425114 146296
rect 423678 145560 423734 145616
rect 510618 146104 510674 146160
rect 498658 144880 498714 144936
rect 499854 144880 499910 144936
rect 396078 59764 396134 59800
rect 396078 59744 396080 59764
rect 396080 59744 396132 59764
rect 396132 59744 396134 59764
rect 397090 59780 397092 59800
rect 397092 59780 397144 59800
rect 397144 59780 397146 59800
rect 397090 59744 397146 59780
rect 416962 59744 417018 59800
rect 418434 59744 418490 59800
rect 422850 59744 422906 59800
rect 423954 59744 424010 59800
rect 403070 59608 403126 59664
rect 404174 59608 404230 59664
rect 412546 59608 412602 59664
rect 397458 57840 397514 57896
rect 399482 57840 399538 57896
rect 400218 57840 400274 57896
rect 401690 57840 401746 57896
rect 404358 57840 404414 57896
rect 405830 57840 405886 57896
rect 407210 57840 407266 57896
rect 408314 57840 408370 57896
rect 408682 57840 408738 57896
rect 409878 57840 409934 57896
rect 411350 57840 411406 57896
rect 411258 56888 411314 56944
rect 418158 59472 418214 59528
rect 423494 59608 423550 59664
rect 420642 59336 420698 59392
rect 421746 59336 421802 59392
rect 480902 59608 480958 59664
rect 425978 59336 426034 59392
rect 428186 59336 428242 59392
rect 453394 59336 453450 59392
rect 463514 59336 463570 59392
rect 485962 59200 486018 59256
rect 414570 57840 414626 57896
rect 415490 57840 415546 57896
rect 416042 57840 416098 57896
rect 426438 57840 426494 57896
rect 427634 57840 427690 57896
rect 427818 57840 427874 57896
rect 429198 57840 429254 57896
rect 430578 57840 430634 57896
rect 432234 57840 432290 57896
rect 433338 57840 433394 57896
rect 433614 57840 433670 57896
rect 435914 57840 435970 57896
rect 436098 57840 436154 57896
rect 438214 57840 438270 57896
rect 438490 57840 438546 57896
rect 438858 57840 438914 57896
rect 440882 57840 440938 57896
rect 443458 57840 443514 57896
rect 448242 57840 448298 57896
rect 470874 57860 470930 57896
rect 470874 57840 470876 57860
rect 470876 57840 470928 57860
rect 470928 57840 470930 57860
rect 412546 56888 412602 56944
rect 412638 56752 412694 56808
rect 430946 57160 431002 57216
rect 433430 57160 433486 57216
rect 435730 57160 435786 57216
rect 478418 57876 478420 57896
rect 478420 57876 478472 57896
rect 478472 57876 478474 57896
rect 478418 57840 478474 57876
rect 503258 57876 503260 57896
rect 503260 57876 503312 57896
rect 503312 57876 503314 57896
rect 503258 57840 503314 57876
rect 503534 57860 503590 57896
rect 518990 288360 519046 288416
rect 518990 287136 519046 287192
rect 518898 244160 518954 244216
rect 518898 184864 518954 184920
rect 519082 284960 519138 285016
rect 518990 182688 519046 182744
rect 518898 79872 518954 79928
rect 580262 458088 580318 458144
rect 580262 404912 580318 404968
rect 519358 357992 519414 358048
rect 519266 289312 519322 289368
rect 519174 284144 519230 284200
rect 519082 179424 519138 179480
rect 519082 178744 519138 178800
rect 519358 288360 519414 288416
rect 580446 378392 580502 378448
rect 580354 351872 580410 351928
rect 580262 325216 580318 325272
rect 519450 285776 519506 285832
rect 519358 244160 519414 244216
rect 519266 184864 519322 184920
rect 519266 181328 519322 181384
rect 518990 78240 519046 78296
rect 519910 284960 519966 285016
rect 580354 272176 580410 272232
rect 580262 232328 580318 232384
rect 580354 192480 580410 192536
rect 520186 182688 520242 182744
rect 519450 179424 519506 179480
rect 519358 139304 519414 139360
rect 519266 76744 519322 76800
rect 580262 152632 580318 152688
rect 520186 79872 520242 79928
rect 519450 75384 519506 75440
rect 519082 74160 519138 74216
rect 503534 57840 503536 57860
rect 503536 57840 503588 57860
rect 503588 57840 503590 57860
rect 438858 55120 438914 55176
rect 580446 112784 580502 112840
rect 580354 72936 580410 72992
rect 580262 33088 580318 33144
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect 319621 632362 319687 632365
rect 392117 632362 392183 632365
rect 319621 632360 392183 632362
rect 319621 632304 319626 632360
rect 319682 632304 392122 632360
rect 392178 632304 392183 632360
rect 319621 632302 392183 632304
rect 319621 632299 319687 632302
rect 392117 632299 392183 632302
rect 315297 632226 315363 632229
rect 419165 632226 419231 632229
rect 315297 632224 419231 632226
rect -960 632090 480 632180
rect 315297 632168 315302 632224
rect 315358 632168 419170 632224
rect 419226 632168 419231 632224
rect 315297 632166 419231 632168
rect 315297 632163 315363 632166
rect 419165 632163 419231 632166
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 40677 632090 40743 632093
rect 346393 632090 346459 632093
rect 40677 632088 346459 632090
rect 40677 632032 40682 632088
rect 40738 632032 346398 632088
rect 346454 632032 346459 632088
rect 40677 632030 346459 632032
rect 40677 632027 40743 632030
rect 346393 632027 346459 632030
rect 53046 630804 53052 630868
rect 53116 630866 53122 630868
rect 328085 630866 328151 630869
rect 53116 630864 328151 630866
rect 53116 630808 328090 630864
rect 328146 630808 328151 630864
rect 53116 630806 328151 630808
rect 53116 630804 53122 630806
rect 328085 630803 328151 630806
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 54334 630668 54340 630732
rect 54404 630730 54410 630732
rect 405365 630730 405431 630733
rect 54404 630728 405431 630730
rect 54404 630672 405370 630728
rect 405426 630672 405431 630728
rect 583520 630716 584960 630806
rect 54404 630670 405431 630672
rect 54404 630668 54410 630670
rect 405365 630667 405431 630670
rect 317781 629642 317847 629645
rect 320038 629642 320098 630224
rect 317781 629640 320098 629642
rect 317781 629584 317786 629640
rect 317842 629584 320098 629640
rect 317781 629582 320098 629584
rect 317781 629579 317847 629582
rect 430941 626514 431007 626517
rect 428782 626512 431007 626514
rect 428782 626456 430946 626512
rect 431002 626456 431007 626512
rect 428782 626454 431007 626456
rect 428782 626144 428842 626454
rect 430941 626451 431007 626454
rect 106365 625290 106431 625293
rect 120022 625290 120028 625292
rect 106365 625288 120028 625290
rect 106365 625232 106370 625288
rect 106426 625232 120028 625288
rect 106365 625230 120028 625232
rect 106365 625227 106431 625230
rect 120022 625228 120028 625230
rect 120092 625228 120098 625292
rect 318149 625290 318215 625293
rect 320038 625290 320098 625464
rect 318149 625288 320098 625290
rect 318149 625232 318154 625288
rect 318210 625232 320098 625288
rect 318149 625230 320098 625232
rect 318149 625227 318215 625230
rect 430849 622026 430915 622029
rect 428782 622024 430915 622026
rect 428782 621968 430854 622024
rect 430910 621968 430915 622024
rect 428782 621966 430915 621968
rect 428782 621384 428842 621966
rect 430849 621963 430915 621966
rect 57697 620666 57763 620669
rect 137369 620666 137435 620669
rect 216673 620666 216739 620669
rect 57697 620664 60076 620666
rect 57697 620608 57702 620664
rect 57758 620608 60076 620664
rect 57697 620606 60076 620608
rect 137369 620664 140116 620666
rect 137369 620608 137374 620664
rect 137430 620608 140116 620664
rect 137369 620606 140116 620608
rect 216673 620664 220156 620666
rect 216673 620608 216678 620664
rect 216734 620608 220156 620664
rect 216673 620606 220156 620608
rect 57697 620603 57763 620606
rect 137369 620603 137435 620606
rect 216673 620603 216739 620606
rect 317965 620122 318031 620125
rect 320038 620122 320098 620704
rect 317965 620120 320098 620122
rect 317965 620064 317970 620120
rect 318026 620064 320098 620120
rect 317965 620062 320098 620064
rect 317965 620059 318031 620062
rect 123017 619986 123083 619989
rect 201585 619986 201651 619989
rect 281625 619986 281691 619989
rect 120796 619984 123083 619986
rect 120796 619928 123022 619984
rect 123078 619928 123083 619984
rect 120796 619926 123083 619928
rect 200836 619984 201651 619986
rect 200836 619928 201590 619984
rect 201646 619928 201651 619984
rect 200836 619926 201651 619928
rect 280876 619984 281691 619986
rect 280876 619928 281630 619984
rect 281686 619928 281691 619984
rect 280876 619926 281691 619928
rect 123017 619923 123083 619926
rect 201585 619923 201651 619926
rect 281625 619923 281691 619926
rect -960 619020 480 619260
rect 456793 619034 456859 619037
rect 456793 619032 460092 619034
rect 456793 618976 456798 619032
rect 456854 618976 460092 619032
rect 456793 618974 460092 618976
rect 456793 618971 456859 618974
rect 59261 617810 59327 617813
rect 59494 617810 60076 617870
rect 139350 617818 140032 617878
rect 219390 617818 220064 617878
rect 139025 617810 139091 617813
rect 139350 617810 139410 617818
rect 59261 617808 59554 617810
rect 59261 617752 59266 617808
rect 59322 617752 59554 617808
rect 59261 617750 59554 617752
rect 139025 617808 139410 617810
rect 139025 617752 139030 617808
rect 139086 617752 139410 617808
rect 139025 617750 139410 617752
rect 216673 617810 216739 617813
rect 219390 617810 219450 617818
rect 216673 617808 219450 617810
rect 216673 617752 216678 617808
rect 216734 617752 219450 617808
rect 216673 617750 219450 617752
rect 59261 617747 59327 617750
rect 139025 617747 139091 617750
rect 216673 617747 216739 617750
rect 583520 617388 584960 617628
rect 123109 617266 123175 617269
rect 202965 617266 203031 617269
rect 281717 617266 281783 617269
rect 120796 617264 123175 617266
rect 120796 617208 123114 617264
rect 123170 617208 123175 617264
rect 120796 617206 123175 617208
rect 200836 617264 203031 617266
rect 200836 617208 202970 617264
rect 203026 617208 203031 617264
rect 200836 617206 203031 617208
rect 280876 617264 281783 617266
rect 280876 617208 281722 617264
rect 281778 617208 281783 617264
rect 280876 617206 281783 617208
rect 123109 617203 123175 617206
rect 202965 617203 203031 617206
rect 281717 617203 281783 617206
rect 430757 616858 430823 616861
rect 428782 616856 430823 616858
rect 428782 616800 430762 616856
rect 430818 616800 430823 616856
rect 428782 616798 430823 616800
rect 428782 616624 428842 616798
rect 430757 616795 430823 616798
rect 317965 615634 318031 615637
rect 320038 615634 320098 615944
rect 510613 615634 510679 615637
rect 317965 615632 320098 615634
rect 317965 615576 317970 615632
rect 318026 615576 320098 615632
rect 317965 615574 320098 615576
rect 509956 615632 510679 615634
rect 509956 615576 510618 615632
rect 510674 615576 510679 615632
rect 509956 615574 510679 615576
rect 317965 615571 318031 615574
rect 510613 615571 510679 615574
rect 57513 614410 57579 614413
rect 59494 614410 60076 614470
rect 139350 614418 140032 614478
rect 219390 614418 220064 614478
rect 138565 614410 138631 614413
rect 139350 614410 139410 614418
rect 57513 614408 59554 614410
rect 57513 614352 57518 614408
rect 57574 614352 59554 614408
rect 57513 614350 59554 614352
rect 138565 614408 139410 614410
rect 138565 614352 138570 614408
rect 138626 614352 139410 614408
rect 138565 614350 139410 614352
rect 217685 614410 217751 614413
rect 219390 614410 219450 614418
rect 217685 614408 219450 614410
rect 217685 614352 217690 614408
rect 217746 614352 219450 614408
rect 217685 614350 219450 614352
rect 57513 614347 57579 614350
rect 138565 614347 138631 614350
rect 217685 614347 217751 614350
rect 121729 613866 121795 613869
rect 201861 613866 201927 613869
rect 283005 613866 283071 613869
rect 120796 613864 121795 613866
rect 120796 613808 121734 613864
rect 121790 613808 121795 613864
rect 120796 613806 121795 613808
rect 200836 613864 201927 613866
rect 200836 613808 201866 613864
rect 201922 613808 201927 613864
rect 200836 613806 201927 613808
rect 280876 613864 283071 613866
rect 280876 613808 283010 613864
rect 283066 613808 283071 613864
rect 280876 613806 283071 613808
rect 121729 613803 121795 613806
rect 201861 613803 201927 613806
rect 283005 613803 283071 613806
rect 430665 612506 430731 612509
rect 428782 612504 430731 612506
rect 428782 612448 430670 612504
rect 430726 612448 430731 612504
rect 428782 612446 430731 612448
rect 428782 611864 428842 612446
rect 430665 612443 430731 612446
rect 59077 611690 59143 611693
rect 59494 611690 60076 611750
rect 139350 611698 140032 611758
rect 219390 611698 220064 611758
rect 137645 611690 137711 611693
rect 139350 611690 139410 611698
rect 59077 611688 59554 611690
rect 59077 611632 59082 611688
rect 59138 611632 59554 611688
rect 59077 611630 59554 611632
rect 137645 611688 139410 611690
rect 137645 611632 137650 611688
rect 137706 611632 139410 611688
rect 137645 611630 139410 611632
rect 215937 611690 216003 611693
rect 219390 611690 219450 611698
rect 215937 611688 219450 611690
rect 215937 611632 215942 611688
rect 215998 611632 219450 611688
rect 215937 611630 219450 611632
rect 59077 611627 59143 611630
rect 137645 611627 137711 611630
rect 215937 611627 216003 611630
rect 121821 611146 121887 611149
rect 281993 611146 282059 611149
rect 120796 611144 121887 611146
rect 120796 611088 121826 611144
rect 121882 611088 121887 611144
rect 280876 611144 282059 611146
rect 120796 611086 121887 611088
rect 121821 611083 121887 611086
rect 200806 610605 200866 611116
rect 280876 611088 281998 611144
rect 282054 611088 282059 611144
rect 280876 611086 282059 611088
rect 281993 611083 282059 611086
rect 200757 610600 200866 610605
rect 200757 610544 200762 610600
rect 200818 610544 200866 610600
rect 200757 610542 200866 610544
rect 317873 610602 317939 610605
rect 320038 610602 320098 611184
rect 456793 610874 456859 610877
rect 456793 610872 460092 610874
rect 456793 610816 456798 610872
rect 456854 610816 460092 610872
rect 456793 610814 460092 610816
rect 456793 610811 456859 610814
rect 317873 610600 320098 610602
rect 317873 610544 317878 610600
rect 317934 610544 320098 610600
rect 317873 610542 320098 610544
rect 200757 610539 200823 610542
rect 317873 610539 317939 610542
rect 58893 608290 58959 608293
rect 59494 608290 60076 608350
rect 139350 608298 140032 608358
rect 219390 608298 220064 608358
rect 136725 608290 136791 608293
rect 139350 608290 139410 608298
rect 58893 608288 59554 608290
rect 58893 608232 58898 608288
rect 58954 608232 59554 608288
rect 58893 608230 59554 608232
rect 136725 608288 139410 608290
rect 136725 608232 136730 608288
rect 136786 608232 139410 608288
rect 136725 608230 139410 608232
rect 216673 608290 216739 608293
rect 219390 608290 219450 608298
rect 216673 608288 219450 608290
rect 216673 608232 216678 608288
rect 216734 608232 219450 608288
rect 216673 608230 219450 608232
rect 58893 608227 58959 608230
rect 136725 608227 136791 608230
rect 216673 608227 216739 608230
rect 123569 607746 123635 607749
rect 202873 607746 202939 607749
rect 283649 607746 283715 607749
rect 120796 607744 123635 607746
rect 120796 607688 123574 607744
rect 123630 607688 123635 607744
rect 120796 607686 123635 607688
rect 200836 607744 202939 607746
rect 200836 607688 202878 607744
rect 202934 607688 202939 607744
rect 200836 607686 202939 607688
rect 280876 607744 283715 607746
rect 280876 607688 283654 607744
rect 283710 607688 283715 607744
rect 280876 607686 283715 607688
rect 123569 607683 123635 607686
rect 202873 607683 202939 607686
rect 283649 607683 283715 607686
rect 511993 607474 512059 607477
rect 509956 607472 512059 607474
rect 509956 607416 511998 607472
rect 512054 607416 512059 607472
rect 509956 607414 512059 607416
rect 511993 607411 512059 607414
rect 430573 607202 430639 607205
rect 428782 607200 430639 607202
rect 428782 607144 430578 607200
rect 430634 607144 430639 607200
rect 428782 607142 430639 607144
rect 428782 607104 428842 607142
rect 430573 607139 430639 607142
rect -960 605964 480 606204
rect 317965 606114 318031 606117
rect 320038 606114 320098 606424
rect 317965 606112 320098 606114
rect 317965 606056 317970 606112
rect 318026 606056 320098 606112
rect 317965 606054 320098 606056
rect 317965 606051 318031 606054
rect 59169 605570 59235 605573
rect 59494 605570 60076 605630
rect 139350 605578 140032 605638
rect 219390 605578 220064 605638
rect 138933 605570 138999 605573
rect 139350 605570 139410 605578
rect 59169 605568 59554 605570
rect 59169 605512 59174 605568
rect 59230 605512 59554 605568
rect 59169 605510 59554 605512
rect 138933 605568 139410 605570
rect 138933 605512 138938 605568
rect 138994 605512 139410 605568
rect 138933 605510 139410 605512
rect 219249 605570 219315 605573
rect 219390 605570 219450 605578
rect 219249 605568 219450 605570
rect 219249 605512 219254 605568
rect 219310 605512 219450 605568
rect 219249 605510 219450 605512
rect 59169 605507 59235 605510
rect 138933 605507 138999 605510
rect 219249 605507 219315 605510
rect 123201 605026 123267 605029
rect 201769 605026 201835 605029
rect 283097 605026 283163 605029
rect 120796 605024 123267 605026
rect 120796 604968 123206 605024
rect 123262 604968 123267 605024
rect 120796 604966 123267 604968
rect 200836 605024 201835 605026
rect 200836 604968 201774 605024
rect 201830 604968 201835 605024
rect 200836 604966 201835 604968
rect 280876 605024 283163 605026
rect 280876 604968 283102 605024
rect 283158 604968 283163 605024
rect 280876 604966 283163 604968
rect 123201 604963 123267 604966
rect 201769 604963 201835 604966
rect 283097 604963 283163 604966
rect 583520 604060 584960 604300
rect 457437 602714 457503 602717
rect 457437 602712 460092 602714
rect 457437 602656 457442 602712
rect 457498 602656 460092 602712
rect 457437 602654 460092 602656
rect 457437 602651 457503 602654
rect 58985 602170 59051 602173
rect 59494 602170 60076 602230
rect 139350 602178 140032 602238
rect 219390 602178 220064 602238
rect 138841 602170 138907 602173
rect 139350 602170 139410 602178
rect 58985 602168 59554 602170
rect 58985 602112 58990 602168
rect 59046 602112 59554 602168
rect 58985 602110 59554 602112
rect 138841 602168 139410 602170
rect 138841 602112 138846 602168
rect 138902 602112 139410 602168
rect 138841 602110 139410 602112
rect 217225 602170 217291 602173
rect 219390 602170 219450 602178
rect 217225 602168 219450 602170
rect 217225 602112 217230 602168
rect 217286 602112 219450 602168
rect 217225 602110 219450 602112
rect 58985 602107 59051 602110
rect 138841 602107 138907 602110
rect 217225 602107 217291 602110
rect 428782 601762 428842 602344
rect 431217 601762 431283 601765
rect 428782 601760 431283 601762
rect 428782 601704 431222 601760
rect 431278 601704 431283 601760
rect 428782 601702 431283 601704
rect 431217 601699 431283 601702
rect 121913 601626 121979 601629
rect 203057 601626 203123 601629
rect 283189 601626 283255 601629
rect 120796 601624 121979 601626
rect 120796 601568 121918 601624
rect 121974 601568 121979 601624
rect 120796 601566 121979 601568
rect 200836 601624 203123 601626
rect 200836 601568 203062 601624
rect 203118 601568 203123 601624
rect 200836 601566 203123 601568
rect 280876 601624 283255 601626
rect 280876 601568 283194 601624
rect 283250 601568 283255 601624
rect 280876 601566 283255 601568
rect 121913 601563 121979 601566
rect 203057 601563 203123 601566
rect 283189 601563 283255 601566
rect 317597 601082 317663 601085
rect 320038 601082 320098 601664
rect 317597 601080 320098 601082
rect 317597 601024 317602 601080
rect 317658 601024 320098 601080
rect 317597 601022 320098 601024
rect 317597 601019 317663 601022
rect 57881 599586 57947 599589
rect 137921 599586 137987 599589
rect 217777 599586 217843 599589
rect 57881 599584 59554 599586
rect 57881 599528 57886 599584
rect 57942 599566 59554 599584
rect 137921 599584 139594 599586
rect 57942 599528 60076 599566
rect 57881 599526 60076 599528
rect 57881 599523 57947 599526
rect 59494 599506 60076 599526
rect 137921 599528 137926 599584
rect 137982 599566 139594 599584
rect 217777 599584 219818 599586
rect 137982 599528 140116 599566
rect 137921 599526 140116 599528
rect 137921 599523 137987 599526
rect 139534 599506 140116 599526
rect 217777 599528 217782 599584
rect 217838 599566 219818 599584
rect 217838 599528 220156 599566
rect 217777 599526 220156 599528
rect 217777 599523 217843 599526
rect 219758 599506 220156 599526
rect 511993 599314 512059 599317
rect 509956 599312 512059 599314
rect 509956 599256 511998 599312
rect 512054 599256 512059 599312
rect 509956 599254 512059 599256
rect 511993 599251 512059 599254
rect 283281 598906 283347 598909
rect 280876 598904 283347 598906
rect 120766 598365 120826 598876
rect 200806 598365 200866 598876
rect 280876 598848 283286 598904
rect 283342 598848 283347 598904
rect 280876 598846 283347 598848
rect 283281 598843 283347 598846
rect 120766 598360 120875 598365
rect 120766 598304 120814 598360
rect 120870 598304 120875 598360
rect 120766 598302 120875 598304
rect 200806 598360 200915 598365
rect 200806 598304 200854 598360
rect 200910 598304 200915 598360
rect 200806 598302 200915 598304
rect 120809 598299 120875 598302
rect 200849 598299 200915 598302
rect 430614 597682 430620 597684
rect 428782 597622 430620 597682
rect 428782 597584 428842 597622
rect 430614 597620 430620 597622
rect 430684 597620 430690 597684
rect 317597 596458 317663 596461
rect 320038 596458 320098 596904
rect 317597 596456 320098 596458
rect 317597 596400 317602 596456
rect 317658 596400 320098 596456
rect 317597 596398 320098 596400
rect 317597 596395 317663 596398
rect 218697 596186 218763 596189
rect 218697 596184 219818 596186
rect 218697 596128 218702 596184
rect 218758 596166 219818 596184
rect 218758 596128 220156 596166
rect 218697 596126 220156 596128
rect 218697 596123 218763 596126
rect 57881 596050 57947 596053
rect 59494 596050 60076 596110
rect 136633 596050 136699 596053
rect 139534 596050 140116 596110
rect 219758 596106 220156 596126
rect 57881 596048 59554 596050
rect 57881 595992 57886 596048
rect 57942 595992 59554 596048
rect 57881 595990 59554 595992
rect 136633 596048 139594 596050
rect 136633 595992 136638 596048
rect 136694 595992 139594 596048
rect 136633 595990 139594 595992
rect 57881 595987 57947 595990
rect 136633 595987 136699 595990
rect 123385 595506 123451 595509
rect 203149 595506 203215 595509
rect 120796 595504 123451 595506
rect 120796 595448 123390 595504
rect 123446 595448 123451 595504
rect 120796 595446 123451 595448
rect 200836 595504 203215 595506
rect 200836 595448 203154 595504
rect 203210 595448 203215 595504
rect 200836 595446 203215 595448
rect 123385 595443 123451 595446
rect 203149 595443 203215 595446
rect 280846 594965 280906 595476
rect 280846 594960 280955 594965
rect 280846 594904 280894 594960
rect 280950 594904 280955 594960
rect 280846 594902 280955 594904
rect 280889 594899 280955 594902
rect 457437 594554 457503 594557
rect 457437 594552 460092 594554
rect 457437 594496 457442 594552
rect 457498 594496 460092 594552
rect 457437 594494 460092 594496
rect 457437 594491 457503 594494
rect 57605 593466 57671 593469
rect 137921 593466 137987 593469
rect 216673 593466 216739 593469
rect 57605 593464 59554 593466
rect 57605 593408 57610 593464
rect 57666 593446 59554 593464
rect 137921 593464 139594 593466
rect 57666 593408 60076 593446
rect 57605 593406 60076 593408
rect 57605 593403 57671 593406
rect 59494 593386 60076 593406
rect 137921 593408 137926 593464
rect 137982 593446 139594 593464
rect 216673 593464 219818 593466
rect 137982 593408 140116 593446
rect 137921 593406 140116 593408
rect 137921 593403 137987 593406
rect 139534 593386 140116 593406
rect 216673 593408 216678 593464
rect 216734 593446 219818 593464
rect 216734 593408 220156 593446
rect 216673 593406 220156 593408
rect 216673 593403 216739 593406
rect 219758 593386 220156 593406
rect -960 592908 480 593148
rect 123293 592786 123359 592789
rect 201953 592786 202019 592789
rect 281165 592786 281231 592789
rect 120796 592784 123359 592786
rect 120796 592728 123298 592784
rect 123354 592728 123359 592784
rect 120796 592726 123359 592728
rect 200836 592784 202019 592786
rect 200836 592728 201958 592784
rect 202014 592728 202019 592784
rect 200836 592726 202019 592728
rect 280876 592784 281231 592786
rect 280876 592728 281170 592784
rect 281226 592728 281231 592784
rect 280876 592726 281231 592728
rect 123293 592723 123359 592726
rect 201953 592723 202019 592726
rect 281165 592723 281231 592726
rect 318793 592786 318859 592789
rect 318793 592784 320098 592786
rect 318793 592728 318798 592784
rect 318854 592728 320098 592784
rect 318793 592726 320098 592728
rect 318793 592723 318859 592726
rect 320038 592144 320098 592726
rect 428782 592242 428842 592824
rect 430798 592242 430804 592244
rect 428782 592182 430804 592242
rect 430798 592180 430804 592182
rect 430868 592180 430874 592244
rect 512085 591154 512151 591157
rect 509956 591152 512151 591154
rect 509956 591096 512090 591152
rect 512146 591096 512151 591152
rect 509956 591094 512151 591096
rect 512085 591091 512151 591094
rect 583520 590868 584960 591108
rect 57421 589930 57487 589933
rect 59494 589930 60076 589990
rect 139350 589938 140032 589998
rect 219390 589938 220064 589998
rect 136909 589930 136975 589933
rect 139350 589930 139410 589938
rect 57421 589928 59554 589930
rect 57421 589872 57426 589928
rect 57482 589872 59554 589928
rect 57421 589870 59554 589872
rect 136909 589928 139410 589930
rect 136909 589872 136914 589928
rect 136970 589872 139410 589928
rect 136909 589870 139410 589872
rect 216673 589930 216739 589933
rect 219390 589930 219450 589938
rect 216673 589928 219450 589930
rect 216673 589872 216678 589928
rect 216734 589872 219450 589928
rect 216673 589870 219450 589872
rect 57421 589867 57487 589870
rect 136909 589867 136975 589870
rect 216673 589867 216739 589870
rect 124121 589386 124187 589389
rect 204161 589386 204227 589389
rect 283557 589386 283623 589389
rect 120796 589384 124187 589386
rect 120796 589328 124126 589384
rect 124182 589328 124187 589384
rect 120796 589326 124187 589328
rect 200836 589384 204227 589386
rect 200836 589328 204166 589384
rect 204222 589328 204227 589384
rect 200836 589326 204227 589328
rect 280876 589384 283623 589386
rect 280876 589328 283562 589384
rect 283618 589328 283623 589384
rect 280876 589326 283623 589328
rect 124121 589323 124187 589326
rect 204161 589323 204227 589326
rect 283557 589323 283623 589326
rect 428782 588026 428842 588064
rect 429469 588026 429535 588029
rect 428782 588024 429535 588026
rect 428782 587968 429474 588024
rect 429530 587968 429535 588024
rect 428782 587966 429535 587968
rect 429469 587963 429535 587966
rect 59494 587210 60076 587270
rect 139350 587218 140032 587278
rect 219390 587218 220064 587278
rect 138749 587210 138815 587213
rect 139350 587210 139410 587218
rect 57329 586394 57395 586397
rect 59494 586394 59554 587210
rect 138749 587208 139410 587210
rect 138749 587152 138754 587208
rect 138810 587152 139410 587208
rect 138749 587150 139410 587152
rect 216673 587210 216739 587213
rect 219390 587210 219450 587218
rect 216673 587208 219450 587210
rect 216673 587152 216678 587208
rect 216734 587152 219450 587208
rect 216673 587150 219450 587152
rect 138749 587147 138815 587150
rect 216673 587147 216739 587150
rect 122189 586666 122255 586669
rect 202229 586666 202295 586669
rect 281809 586666 281875 586669
rect 120796 586664 122255 586666
rect 120796 586608 122194 586664
rect 122250 586608 122255 586664
rect 120796 586606 122255 586608
rect 200836 586664 202295 586666
rect 200836 586608 202234 586664
rect 202290 586608 202295 586664
rect 200836 586606 202295 586608
rect 280876 586664 281875 586666
rect 280876 586608 281814 586664
rect 281870 586608 281875 586664
rect 280876 586606 281875 586608
rect 122189 586603 122255 586606
rect 202229 586603 202295 586606
rect 281809 586603 281875 586606
rect 317413 586530 317479 586533
rect 317413 586528 317522 586530
rect 317413 586472 317418 586528
rect 317474 586472 317522 586528
rect 317413 586467 317522 586472
rect 57329 586392 59554 586394
rect 57329 586336 57334 586392
rect 57390 586336 59554 586392
rect 57329 586334 59554 586336
rect 317462 586394 317522 586467
rect 320038 586394 320098 587384
rect 317462 586334 320098 586394
rect 457529 586394 457595 586397
rect 457529 586392 460092 586394
rect 457529 586336 457534 586392
rect 457590 586336 460092 586392
rect 457529 586334 460092 586336
rect 57329 586331 57395 586334
rect 457529 586331 457595 586334
rect 59494 583810 60076 583870
rect 139350 583818 140032 583878
rect 219390 583818 220064 583878
rect 137461 583810 137527 583813
rect 139350 583810 139410 583818
rect 57470 583750 59554 583810
rect 137461 583808 139410 583810
rect 137461 583752 137466 583808
rect 137522 583752 139410 583808
rect 137461 583750 139410 583752
rect 217409 583810 217475 583813
rect 219390 583810 219450 583818
rect 217409 583808 219450 583810
rect 217409 583752 217414 583808
rect 217470 583752 219450 583808
rect 217409 583750 219450 583752
rect 57470 583677 57530 583750
rect 137461 583747 137527 583750
rect 217409 583747 217475 583750
rect 57470 583672 57579 583677
rect 57470 583616 57518 583672
rect 57574 583616 57579 583672
rect 57470 583614 57579 583616
rect 57513 583611 57579 583614
rect 122097 583266 122163 583269
rect 202045 583266 202111 583269
rect 283373 583266 283439 583269
rect 120796 583264 122163 583266
rect 120796 583208 122102 583264
rect 122158 583208 122163 583264
rect 120796 583206 122163 583208
rect 200836 583264 202111 583266
rect 200836 583208 202050 583264
rect 202106 583208 202111 583264
rect 200836 583206 202111 583208
rect 280876 583264 283439 583266
rect 280876 583208 283378 583264
rect 283434 583208 283439 583264
rect 280876 583206 283439 583208
rect 122097 583203 122163 583206
rect 202045 583203 202111 583206
rect 283373 583203 283439 583206
rect 428782 582722 428842 583304
rect 511257 582994 511323 582997
rect 509956 582992 511323 582994
rect 509956 582936 511262 582992
rect 511318 582936 511323 582992
rect 509956 582934 511323 582936
rect 511257 582931 511323 582934
rect 429377 582722 429443 582725
rect 428782 582720 429443 582722
rect 428782 582664 429382 582720
rect 429438 582664 429443 582720
rect 428782 582662 429443 582664
rect 429377 582659 429443 582662
rect 317965 582586 318031 582589
rect 320038 582586 320098 582624
rect 317965 582584 320098 582586
rect 317965 582528 317970 582584
rect 318026 582528 320098 582584
rect 317965 582526 320098 582528
rect 317965 582523 318031 582526
rect 58801 581090 58867 581093
rect 59494 581090 60076 581150
rect 139350 581098 140032 581158
rect 219390 581098 220064 581158
rect 138657 581090 138723 581093
rect 139350 581090 139410 581098
rect 58801 581088 59554 581090
rect 58801 581032 58806 581088
rect 58862 581032 59554 581088
rect 58801 581030 59554 581032
rect 138657 581088 139410 581090
rect 138657 581032 138662 581088
rect 138718 581032 139410 581088
rect 138657 581030 139410 581032
rect 217685 581090 217751 581093
rect 219390 581090 219450 581098
rect 217685 581088 219450 581090
rect 217685 581032 217690 581088
rect 217746 581032 219450 581088
rect 217685 581030 219450 581032
rect 58801 581027 58867 581030
rect 138657 581027 138723 581030
rect 217685 581027 217751 581030
rect 122005 580546 122071 580549
rect 202137 580546 202203 580549
rect 283465 580546 283531 580549
rect 120796 580544 122071 580546
rect 120796 580488 122010 580544
rect 122066 580488 122071 580544
rect 120796 580486 122071 580488
rect 200836 580544 202203 580546
rect 200836 580488 202142 580544
rect 202198 580488 202203 580544
rect 200836 580486 202203 580488
rect 280876 580544 283531 580546
rect 280876 580488 283470 580544
rect 283526 580488 283531 580544
rect 280876 580486 283531 580488
rect 122005 580483 122071 580486
rect 202137 580483 202203 580486
rect 283465 580483 283531 580486
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 428782 578370 428842 578544
rect 430665 578370 430731 578373
rect 428782 578368 430731 578370
rect 428782 578312 430670 578368
rect 430726 578312 430731 578368
rect 428782 578310 430731 578312
rect 430665 578307 430731 578310
rect 457621 578234 457687 578237
rect 457621 578232 460092 578234
rect 457621 578176 457626 578232
rect 457682 578176 460092 578232
rect 457621 578174 460092 578176
rect 457621 578171 457687 578174
rect 57053 577690 57119 577693
rect 59494 577690 60076 577750
rect 139350 577698 140032 577758
rect 219390 577698 220064 577758
rect 136725 577690 136791 577693
rect 139350 577690 139410 577698
rect 57053 577688 59554 577690
rect 57053 577632 57058 577688
rect 57114 577632 59554 577688
rect 57053 577630 59554 577632
rect 136725 577688 139410 577690
rect 136725 577632 136730 577688
rect 136786 577632 139410 577688
rect 136725 577630 139410 577632
rect 216029 577690 216095 577693
rect 219390 577690 219450 577698
rect 216029 577688 219450 577690
rect 216029 577632 216034 577688
rect 216090 577632 219450 577688
rect 216029 577630 219450 577632
rect 57053 577627 57119 577630
rect 136725 577627 136791 577630
rect 216029 577627 216095 577630
rect 317873 577282 317939 577285
rect 320038 577282 320098 577864
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 317873 577280 320098 577282
rect 317873 577224 317878 577280
rect 317934 577224 320098 577280
rect 317873 577222 320098 577224
rect 317873 577219 317939 577222
rect 203241 577146 203307 577149
rect 281901 577146 281967 577149
rect 200836 577144 203307 577146
rect 120766 576874 120826 577116
rect 200836 577088 203246 577144
rect 203302 577088 203307 577144
rect 200836 577086 203307 577088
rect 280876 577144 281967 577146
rect 280876 577088 281906 577144
rect 281962 577088 281967 577144
rect 280876 577086 281967 577088
rect 203241 577083 203307 577086
rect 281901 577083 281967 577086
rect 120993 576874 121059 576877
rect 120766 576872 121059 576874
rect 120766 576816 120998 576872
rect 121054 576816 121059 576872
rect 120766 576814 121059 576816
rect 120993 576811 121059 576814
rect 57145 574970 57211 574973
rect 59494 574970 60076 575030
rect 139350 574978 140032 575038
rect 219390 574978 220064 575038
rect 137277 574970 137343 574973
rect 139350 574970 139410 574978
rect 57145 574968 59554 574970
rect 57145 574912 57150 574968
rect 57206 574912 59554 574968
rect 57145 574910 59554 574912
rect 137277 574968 139410 574970
rect 137277 574912 137282 574968
rect 137338 574912 139410 574968
rect 137277 574910 139410 574912
rect 216673 574970 216739 574973
rect 219390 574970 219450 574978
rect 216673 574968 219450 574970
rect 216673 574912 216678 574968
rect 216734 574912 219450 574968
rect 216673 574910 219450 574912
rect 57145 574907 57211 574910
rect 137277 574907 137343 574910
rect 216673 574907 216739 574910
rect 512177 574834 512243 574837
rect 509956 574832 512243 574834
rect 509956 574776 512182 574832
rect 512238 574776 512243 574832
rect 509956 574774 512243 574776
rect 512177 574771 512243 574774
rect 123477 574426 123543 574429
rect 282913 574426 282979 574429
rect 120796 574424 123543 574426
rect 120796 574368 123482 574424
rect 123538 574368 123543 574424
rect 280876 574424 282979 574426
rect 120796 574366 123543 574368
rect 123477 574363 123543 574366
rect 200806 574154 200866 574396
rect 280876 574368 282918 574424
rect 282974 574368 282979 574424
rect 280876 574366 282979 574368
rect 282913 574363 282979 574366
rect 200941 574154 201007 574157
rect 200806 574152 201007 574154
rect 200806 574096 200946 574152
rect 201002 574096 201007 574152
rect 200806 574094 201007 574096
rect 200941 574091 201007 574094
rect 428782 572794 428842 573104
rect 430757 572794 430823 572797
rect 428782 572792 430823 572794
rect 428782 572736 430762 572792
rect 430818 572736 430823 572792
rect 428782 572734 430823 572736
rect 430757 572731 430823 572734
rect 317965 571842 318031 571845
rect 320038 571842 320098 572424
rect 317965 571840 320098 571842
rect 317965 571784 317970 571840
rect 318026 571784 320098 571840
rect 317965 571782 320098 571784
rect 317965 571779 318031 571782
rect 57329 571570 57395 571573
rect 59494 571570 60076 571630
rect 139350 571578 140032 571638
rect 219390 571578 220064 571638
rect 137553 571570 137619 571573
rect 139350 571570 139410 571578
rect 57329 571568 59554 571570
rect 57329 571512 57334 571568
rect 57390 571512 59554 571568
rect 57329 571510 59554 571512
rect 137553 571568 139410 571570
rect 137553 571512 137558 571568
rect 137614 571512 139410 571568
rect 137553 571510 139410 571512
rect 216673 571570 216739 571573
rect 219390 571570 219450 571578
rect 216673 571568 219450 571570
rect 216673 571512 216678 571568
rect 216734 571512 219450 571568
rect 216673 571510 219450 571512
rect 57329 571507 57395 571510
rect 137553 571507 137619 571510
rect 216673 571507 216739 571510
rect 121453 571026 121519 571029
rect 202321 571026 202387 571029
rect 283557 571026 283623 571029
rect 120796 571024 121519 571026
rect 120796 570968 121458 571024
rect 121514 570968 121519 571024
rect 120796 570966 121519 570968
rect 200836 571024 202387 571026
rect 200836 570968 202326 571024
rect 202382 570968 202387 571024
rect 200836 570966 202387 570968
rect 280876 571024 283623 571026
rect 280876 570968 283562 571024
rect 283618 570968 283623 571024
rect 280876 570966 283623 570968
rect 121453 570963 121519 570966
rect 202321 570963 202387 570966
rect 283557 570963 283623 570966
rect 58525 568850 58591 568853
rect 59494 568850 60076 568910
rect 139350 568858 140032 568918
rect 219390 568858 220064 568918
rect 137185 568850 137251 568853
rect 139350 568850 139410 568858
rect 58525 568848 59554 568850
rect 58525 568792 58530 568848
rect 58586 568792 59554 568848
rect 58525 568790 59554 568792
rect 137185 568848 139410 568850
rect 137185 568792 137190 568848
rect 137246 568792 139410 568848
rect 137185 568790 139410 568792
rect 219157 568850 219223 568853
rect 219390 568850 219450 568858
rect 219157 568848 219450 568850
rect 219157 568792 219162 568848
rect 219218 568792 219450 568848
rect 219157 568790 219450 568792
rect 58525 568787 58591 568790
rect 137185 568787 137251 568790
rect 219157 568787 219223 568790
rect 122925 568306 122991 568309
rect 201033 568306 201099 568309
rect 281533 568306 281599 568309
rect 120796 568304 122991 568306
rect 120796 568248 122930 568304
rect 122986 568248 122991 568304
rect 120796 568246 122991 568248
rect 200836 568304 201099 568306
rect 200836 568248 201038 568304
rect 201094 568248 201099 568304
rect 200836 568246 201099 568248
rect 280876 568304 281599 568306
rect 280876 568248 281538 568304
rect 281594 568248 281599 568304
rect 280876 568246 281599 568248
rect 122925 568243 122991 568246
rect 201033 568243 201099 568246
rect 281533 568243 281599 568246
rect 317045 568306 317111 568309
rect 317045 568304 320098 568306
rect 317045 568248 317050 568304
rect 317106 568248 320098 568304
rect 317045 568246 320098 568248
rect 317045 568243 317111 568246
rect 320038 567664 320098 568246
rect 428782 567762 428842 568344
rect 430849 567762 430915 567765
rect 428782 567760 430915 567762
rect 428782 567704 430854 567760
rect 430910 567704 430915 567760
rect 428782 567702 430915 567704
rect 430849 567699 430915 567702
rect -960 566796 480 567036
rect 57237 565450 57303 565453
rect 59494 565450 60076 565510
rect 139350 565458 140032 565518
rect 219390 565458 220064 565518
rect 139350 565453 139410 565458
rect 57237 565448 59554 565450
rect 57237 565392 57242 565448
rect 57298 565392 59554 565448
rect 57237 565390 59554 565392
rect 139301 565448 139410 565453
rect 139301 565392 139306 565448
rect 139362 565392 139410 565448
rect 139301 565390 139410 565392
rect 217593 565450 217659 565453
rect 219390 565450 219450 565458
rect 217593 565448 219450 565450
rect 217593 565392 217598 565448
rect 217654 565392 219450 565448
rect 217593 565390 219450 565392
rect 57237 565387 57303 565390
rect 139301 565387 139367 565390
rect 217593 565387 217659 565390
rect 121085 564906 121151 564909
rect 203333 564906 203399 564909
rect 281257 564906 281323 564909
rect 120796 564904 121151 564906
rect 120796 564848 121090 564904
rect 121146 564848 121151 564904
rect 120796 564846 121151 564848
rect 200836 564904 203399 564906
rect 200836 564848 203338 564904
rect 203394 564848 203399 564904
rect 200836 564846 203399 564848
rect 280876 564904 281323 564906
rect 280876 564848 281262 564904
rect 281318 564848 281323 564904
rect 280876 564846 281323 564848
rect 121085 564843 121151 564846
rect 203333 564843 203399 564846
rect 281257 564843 281323 564846
rect 583520 564212 584960 564452
rect 428782 563138 428842 563584
rect 430941 563138 431007 563141
rect 428782 563136 431007 563138
rect 428782 563080 430946 563136
rect 431002 563080 431007 563136
rect 428782 563078 431007 563080
rect 430941 563075 431007 563078
rect 59537 562790 59603 562793
rect 59537 562788 60076 562790
rect 59537 562732 59542 562788
rect 59598 562732 60076 562788
rect 139350 562738 140032 562798
rect 219390 562738 220064 562798
rect 59537 562730 60076 562732
rect 138473 562730 138539 562733
rect 139350 562730 139410 562738
rect 59537 562727 59603 562730
rect 138473 562728 139410 562730
rect 138473 562672 138478 562728
rect 138534 562672 139410 562728
rect 138473 562670 139410 562672
rect 217133 562730 217199 562733
rect 219390 562730 219450 562738
rect 217133 562728 219450 562730
rect 217133 562672 217138 562728
rect 217194 562672 219450 562728
rect 217133 562670 219450 562672
rect 138473 562667 138539 562670
rect 217133 562667 217199 562670
rect 318333 562322 318399 562325
rect 320038 562322 320098 562904
rect 318333 562320 320098 562322
rect 318333 562264 318338 562320
rect 318394 562264 320098 562320
rect 318333 562262 320098 562264
rect 318333 562259 318399 562262
rect 121177 562186 121243 562189
rect 201125 562186 201191 562189
rect 281533 562186 281599 562189
rect 120796 562184 121243 562186
rect 120796 562128 121182 562184
rect 121238 562128 121243 562184
rect 120796 562126 121243 562128
rect 200836 562184 201191 562186
rect 200836 562128 201130 562184
rect 201186 562128 201191 562184
rect 200836 562126 201191 562128
rect 280876 562184 281599 562186
rect 280876 562128 281538 562184
rect 281594 562128 281599 562184
rect 280876 562126 281599 562128
rect 121177 562123 121243 562126
rect 201125 562123 201191 562126
rect 281533 562123 281599 562126
rect 86953 559602 87019 559605
rect 120022 559602 120028 559604
rect 86953 559600 120028 559602
rect 86953 559544 86958 559600
rect 87014 559544 120028 559600
rect 86953 559542 120028 559544
rect 86953 559539 87019 559542
rect 120022 559540 120028 559542
rect 120092 559540 120098 559604
rect 428414 558245 428474 558824
rect 428365 558240 428474 558245
rect 428365 558184 428370 558240
rect 428426 558184 428474 558240
rect 428365 558182 428474 558184
rect 428365 558179 428431 558182
rect 317413 557698 317479 557701
rect 320038 557698 320098 558144
rect 317413 557696 320098 557698
rect 317413 557640 317418 557696
rect 317474 557640 320098 557696
rect 317413 557638 320098 557640
rect 317413 557635 317479 557638
rect -960 553740 480 553980
rect 317965 553482 318031 553485
rect 428782 553482 428842 554064
rect 431033 553482 431099 553485
rect 317965 553480 320098 553482
rect 317965 553424 317970 553480
rect 318026 553424 320098 553480
rect 317965 553422 320098 553424
rect 428782 553480 431099 553482
rect 428782 553424 431038 553480
rect 431094 553424 431099 553480
rect 428782 553422 431099 553424
rect 317965 553419 318031 553422
rect 320038 553384 320098 553422
rect 431033 553419 431099 553422
rect 583520 551020 584960 551260
rect 429561 549402 429627 549405
rect 428782 549400 429627 549402
rect 428782 549344 429566 549400
rect 429622 549344 429627 549400
rect 428782 549342 429627 549344
rect 428782 549304 428842 549342
rect 429561 549339 429627 549342
rect 317505 549130 317571 549133
rect 317505 549128 320098 549130
rect 317505 549072 317510 549128
rect 317566 549072 320098 549128
rect 317505 549070 320098 549072
rect 317505 549067 317571 549070
rect 320038 548624 320098 549070
rect 428782 543962 428842 544544
rect 431125 543962 431191 543965
rect 428782 543960 431191 543962
rect 428782 543904 431130 543960
rect 431186 543904 431191 543960
rect 428782 543902 431191 543904
rect 431125 543899 431191 543902
rect 317965 543826 318031 543829
rect 320038 543826 320098 543864
rect 317965 543824 320098 543826
rect 317965 543768 317970 543824
rect 318026 543768 320098 543824
rect 317965 543766 320098 543768
rect 317965 543763 318031 543766
rect 238661 543146 238727 543149
rect 300158 543146 300164 543148
rect 238661 543144 300164 543146
rect 238661 543088 238666 543144
rect 238722 543088 300164 543144
rect 238661 543086 300164 543088
rect 238661 543083 238727 543086
rect 300158 543084 300164 543086
rect 300228 543084 300234 543148
rect 245837 543010 245903 543013
rect 318057 543010 318123 543013
rect 245837 543008 318123 543010
rect 245837 542952 245842 543008
rect 245898 542952 318062 543008
rect 318118 542952 318123 543008
rect 245837 542950 318123 542952
rect 245837 542947 245903 542950
rect 318057 542947 318123 542950
rect 248689 542874 248755 542877
rect 301589 542874 301655 542877
rect 248689 542872 301655 542874
rect 248689 542816 248694 542872
rect 248750 542816 301594 542872
rect 301650 542816 301655 542872
rect 248689 542814 301655 542816
rect 248689 542811 248755 542814
rect 301589 542811 301655 542814
rect 241513 542738 241579 542741
rect 299974 542738 299980 542740
rect 241513 542736 299980 542738
rect 241513 542680 241518 542736
rect 241574 542680 299980 542736
rect 241513 542678 299980 542680
rect 241513 542675 241579 542678
rect 299974 542676 299980 542678
rect 300044 542676 300050 542740
rect 293125 542602 293191 542605
rect 318241 542602 318307 542605
rect 293125 542600 318307 542602
rect 293125 542544 293130 542600
rect 293186 542544 318246 542600
rect 318302 542544 318307 542600
rect 293125 542542 318307 542544
rect 293125 542539 293191 542542
rect 318241 542539 318307 542542
rect 255129 542466 255195 542469
rect 319529 542466 319595 542469
rect 255129 542464 319595 542466
rect 255129 542408 255134 542464
rect 255190 542408 319534 542464
rect 319590 542408 319595 542464
rect 255129 542406 319595 542408
rect 255129 542403 255195 542406
rect 319529 542403 319595 542406
rect 282913 541650 282979 541653
rect 316861 541650 316927 541653
rect 282913 541648 316927 541650
rect 282913 541592 282918 541648
rect 282974 541592 316866 541648
rect 316922 541592 316927 541648
rect 282913 541590 316927 541592
rect 282913 541587 282979 541590
rect 316861 541587 316927 541590
rect 294505 541242 294571 541245
rect 317229 541242 317295 541245
rect 294505 541240 317295 541242
rect 294505 541184 294510 541240
rect 294566 541184 317234 541240
rect 317290 541184 317295 541240
rect 294505 541182 317295 541184
rect 294505 541179 294571 541182
rect 317229 541179 317295 541182
rect 264421 541106 264487 541109
rect 320582 541106 320588 541108
rect 264421 541104 320588 541106
rect 264421 541048 264426 541104
rect 264482 541048 320588 541104
rect 264421 541046 320588 541048
rect 264421 541043 264487 541046
rect 320582 541044 320588 541046
rect 320652 541044 320658 541108
rect -960 540684 480 540924
rect 428782 539610 428842 539784
rect 430573 539610 430639 539613
rect 428782 539608 430639 539610
rect 428782 539552 430578 539608
rect 430634 539552 430639 539608
rect 428782 539550 430639 539552
rect 430573 539547 430639 539550
rect 318057 539338 318123 539341
rect 318057 539336 320098 539338
rect 318057 539280 318062 539336
rect 318118 539280 320098 539336
rect 318057 539278 320098 539280
rect 318057 539275 318123 539278
rect 320038 539104 320098 539278
rect 583520 537692 584960 537932
rect 317597 534986 317663 534989
rect 317597 534984 320098 534986
rect 317597 534928 317602 534984
rect 317658 534928 320098 534984
rect 317597 534926 320098 534928
rect 317597 534923 317663 534926
rect 320038 534344 320098 534926
rect 428782 534442 428842 535024
rect 431309 534442 431375 534445
rect 428782 534440 431375 534442
rect 428782 534384 431314 534440
rect 431370 534384 431375 534440
rect 428782 534382 431375 534384
rect 431309 534379 431375 534382
rect 302233 532402 302299 532405
rect 299828 532400 302299 532402
rect 299828 532344 302238 532400
rect 302294 532344 302299 532400
rect 299828 532342 302299 532344
rect 302233 532339 302299 532342
rect 429285 530294 429351 530297
rect 428812 530292 429351 530294
rect 428812 530236 429290 530292
rect 429346 530236 429351 530292
rect 428812 530234 429351 530236
rect 429285 530231 429351 530234
rect 317597 529818 317663 529821
rect 317597 529816 320098 529818
rect 317597 529760 317602 529816
rect 317658 529760 320098 529816
rect 317597 529758 320098 529760
rect 317597 529755 317663 529758
rect 320038 529584 320098 529758
rect -960 527764 480 528004
rect 317597 525466 317663 525469
rect 317597 525464 320098 525466
rect 317597 525408 317602 525464
rect 317658 525408 320098 525464
rect 317597 525406 320098 525408
rect 317597 525403 317663 525406
rect 320038 524824 320098 525406
rect 428782 524922 428842 525504
rect 430573 524922 430639 524925
rect 428782 524920 430639 524922
rect 428782 524864 430578 524920
rect 430634 524864 430639 524920
rect 428782 524862 430639 524864
rect 430573 524859 430639 524862
rect 583520 524364 584960 524604
rect 427813 520298 427879 520301
rect 428230 520298 428290 520744
rect 427813 520296 428290 520298
rect 427813 520240 427818 520296
rect 427874 520240 428290 520296
rect 427813 520238 428290 520240
rect 427813 520235 427879 520238
rect 300158 520100 300164 520164
rect 300228 520162 300234 520164
rect 430665 520162 430731 520165
rect 300228 520160 430731 520162
rect 300228 520104 430670 520160
rect 430726 520104 430731 520160
rect 300228 520102 430731 520104
rect 300228 520100 300234 520102
rect 430665 520099 430731 520102
rect 301589 518802 301655 518805
rect 430614 518802 430620 518804
rect 301589 518800 430620 518802
rect 301589 518744 301594 518800
rect 301650 518744 430620 518800
rect 301589 518742 430620 518744
rect 301589 518739 301655 518742
rect 430614 518740 430620 518742
rect 430684 518740 430690 518804
rect 320766 518604 320772 518668
rect 320836 518666 320842 518668
rect 374453 518666 374519 518669
rect 320836 518664 374519 518666
rect 320836 518608 374458 518664
rect 374514 518608 374519 518664
rect 320836 518606 374519 518608
rect 320836 518604 320842 518606
rect 374453 518603 374519 518606
rect 319345 518530 319411 518533
rect 356237 518530 356303 518533
rect 319345 518528 356303 518530
rect 319345 518472 319350 518528
rect 319406 518472 356242 518528
rect 356298 518472 356303 518528
rect 319345 518470 356303 518472
rect 319345 518467 319411 518470
rect 356237 518467 356303 518470
rect 319897 518394 319963 518397
rect 337653 518394 337719 518397
rect 319897 518392 337719 518394
rect 319897 518336 319902 518392
rect 319958 518336 337658 518392
rect 337714 518336 337719 518392
rect 319897 518334 337719 518336
rect 319897 518331 319963 518334
rect 337653 518331 337719 518334
rect 302877 517442 302943 517445
rect 299828 517440 302943 517442
rect 299828 517384 302882 517440
rect 302938 517384 302943 517440
rect 299828 517382 302943 517384
rect 302877 517379 302943 517382
rect 299974 517244 299980 517308
rect 300044 517306 300050 517308
rect 430798 517306 430804 517308
rect 300044 517246 430804 517306
rect 300044 517244 300050 517246
rect 430798 517244 430804 517246
rect 430868 517244 430874 517308
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 57697 509962 57763 509965
rect 57881 509962 57947 509965
rect 57697 509960 60076 509962
rect 57697 509904 57702 509960
rect 57758 509904 57886 509960
rect 57942 509904 60076 509960
rect 57697 509902 60076 509904
rect 57697 509899 57763 509902
rect 57881 509899 57947 509902
rect 302969 502482 303035 502485
rect 299828 502480 303035 502482
rect 299828 502424 302974 502480
rect 303030 502424 303035 502480
rect 299828 502422 303035 502424
rect 302969 502419 303035 502422
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 302877 487522 302943 487525
rect 299828 487520 302943 487522
rect 299828 487464 302882 487520
rect 302938 487464 302943 487520
rect 299828 487462 302943 487464
rect 302877 487459 302943 487462
rect 360694 485012 360700 485076
rect 360764 485074 360770 485076
rect 391933 485074 391999 485077
rect 360764 485072 391999 485074
rect 360764 485016 391938 485072
rect 391994 485016 391999 485072
rect 360764 485014 391999 485016
rect 360764 485012 360770 485014
rect 391933 485011 391999 485014
rect 583520 484516 584960 484756
rect 59302 478756 59308 478820
rect 59372 478818 59378 478820
rect 68645 478818 68711 478821
rect 59372 478816 68711 478818
rect 59372 478760 68650 478816
rect 68706 478760 68711 478816
rect 59372 478758 68711 478760
rect 59372 478756 59378 478758
rect 68645 478755 68711 478758
rect 68921 478818 68987 478821
rect 79501 478818 79567 478821
rect 68921 478816 79567 478818
rect 68921 478760 68926 478816
rect 68982 478760 79506 478816
rect 79562 478760 79567 478816
rect 68921 478758 79567 478760
rect 68921 478755 68987 478758
rect 79501 478755 79567 478758
rect 172881 478818 172947 478821
rect 202454 478818 202460 478820
rect 172881 478816 202460 478818
rect 172881 478760 172886 478816
rect 172942 478760 202460 478816
rect 172881 478758 202460 478760
rect 172881 478755 172947 478758
rect 202454 478756 202460 478758
rect 202524 478756 202530 478820
rect 235901 478818 235967 478821
rect 357934 478818 357940 478820
rect 235901 478816 357940 478818
rect 235901 478760 235906 478816
rect 235962 478760 357940 478816
rect 235901 478758 357940 478760
rect 235901 478755 235967 478758
rect 357934 478756 357940 478758
rect 358004 478756 358010 478820
rect 46790 478620 46796 478684
rect 46860 478682 46866 478684
rect 66345 478682 66411 478685
rect 46860 478680 66411 478682
rect 46860 478624 66350 478680
rect 66406 478624 66411 478680
rect 46860 478622 66411 478624
rect 46860 478620 46866 478622
rect 66345 478619 66411 478622
rect 75821 478682 75887 478685
rect 78673 478682 78739 478685
rect 75821 478680 78739 478682
rect 75821 478624 75826 478680
rect 75882 478624 78678 478680
rect 78734 478624 78739 478680
rect 75821 478622 78739 478624
rect 75821 478619 75887 478622
rect 78673 478619 78739 478622
rect 167177 478682 167243 478685
rect 198038 478682 198044 478684
rect 167177 478680 198044 478682
rect 167177 478624 167182 478680
rect 167238 478624 198044 478680
rect 167177 478622 198044 478624
rect 167177 478619 167243 478622
rect 198038 478620 198044 478622
rect 198108 478620 198114 478684
rect 211337 478682 211403 478685
rect 211838 478682 211844 478684
rect 211337 478680 211844 478682
rect 211337 478624 211342 478680
rect 211398 478624 211844 478680
rect 211337 478622 211844 478624
rect 211337 478619 211403 478622
rect 211838 478620 211844 478622
rect 211908 478620 211914 478684
rect 236269 478682 236335 478685
rect 360142 478682 360148 478684
rect 236269 478680 360148 478682
rect 236269 478624 236274 478680
rect 236330 478624 360148 478680
rect 236269 478622 360148 478624
rect 236269 478619 236335 478622
rect 360142 478620 360148 478622
rect 360212 478620 360218 478684
rect 53230 478484 53236 478548
rect 53300 478546 53306 478548
rect 77753 478546 77819 478549
rect 53300 478544 77819 478546
rect 53300 478488 77758 478544
rect 77814 478488 77819 478544
rect 53300 478486 77819 478488
rect 53300 478484 53306 478486
rect 77753 478483 77819 478486
rect 163589 478546 163655 478549
rect 196566 478546 196572 478548
rect 163589 478544 196572 478546
rect 163589 478488 163594 478544
rect 163650 478488 196572 478544
rect 163589 478486 196572 478488
rect 163589 478483 163655 478486
rect 196566 478484 196572 478486
rect 196636 478484 196642 478548
rect 200757 478546 200823 478549
rect 201350 478546 201356 478548
rect 200757 478544 201356 478546
rect 200757 478488 200762 478544
rect 200818 478488 201356 478544
rect 200757 478486 201356 478488
rect 200757 478483 200823 478486
rect 201350 478484 201356 478486
rect 201420 478484 201426 478548
rect 205633 478546 205699 478549
rect 206686 478546 206692 478548
rect 205633 478544 206692 478546
rect 205633 478488 205638 478544
rect 205694 478488 206692 478544
rect 205633 478486 206692 478488
rect 205633 478483 205699 478486
rect 206686 478484 206692 478486
rect 206756 478484 206762 478548
rect 233233 478546 233299 478549
rect 367686 478546 367692 478548
rect 233233 478544 367692 478546
rect 233233 478488 233238 478544
rect 233294 478488 367692 478544
rect 233233 478486 367692 478488
rect 233233 478483 233299 478486
rect 367686 478484 367692 478486
rect 367756 478484 367762 478548
rect 50061 478410 50127 478413
rect 77293 478410 77359 478413
rect 50061 478408 77359 478410
rect 50061 478352 50066 478408
rect 50122 478352 77298 478408
rect 77354 478352 77359 478408
rect 50061 478350 77359 478352
rect 50061 478347 50127 478350
rect 77293 478347 77359 478350
rect 147305 478410 147371 478413
rect 197854 478410 197860 478412
rect 147305 478408 197860 478410
rect 147305 478352 147310 478408
rect 147366 478352 197860 478408
rect 147305 478350 197860 478352
rect 147305 478347 147371 478350
rect 197854 478348 197860 478350
rect 197924 478348 197930 478412
rect 201585 478410 201651 478413
rect 202638 478410 202644 478412
rect 201585 478408 202644 478410
rect 201585 478352 201590 478408
rect 201646 478352 202644 478408
rect 201585 478350 202644 478352
rect 201585 478347 201651 478350
rect 202638 478348 202644 478350
rect 202708 478348 202714 478412
rect 231485 478410 231551 478413
rect 371734 478410 371740 478412
rect 231485 478408 371740 478410
rect 231485 478352 231490 478408
rect 231546 478352 371740 478408
rect 231485 478350 371740 478352
rect 231485 478347 231551 478350
rect 371734 478348 371740 478350
rect 371804 478348 371810 478412
rect 57646 478212 57652 478276
rect 57716 478274 57722 478276
rect 91369 478274 91435 478277
rect 57716 478272 91435 478274
rect 57716 478216 91374 478272
rect 91430 478216 91435 478272
rect 57716 478214 91435 478216
rect 57716 478212 57722 478214
rect 91369 478211 91435 478214
rect 148225 478274 148291 478277
rect 202086 478274 202092 478276
rect 148225 478272 202092 478274
rect 148225 478216 148230 478272
rect 148286 478216 202092 478272
rect 148225 478214 202092 478216
rect 148225 478211 148291 478214
rect 202086 478212 202092 478214
rect 202156 478212 202162 478276
rect 210233 478274 210299 478277
rect 210734 478274 210740 478276
rect 210233 478272 210740 478274
rect 210233 478216 210238 478272
rect 210294 478216 210740 478272
rect 210233 478214 210740 478216
rect 210233 478211 210299 478214
rect 210734 478212 210740 478214
rect 210804 478212 210810 478276
rect 219198 478212 219204 478276
rect 219268 478274 219274 478276
rect 226149 478274 226215 478277
rect 219268 478272 226215 478274
rect 219268 478216 226154 478272
rect 226210 478216 226215 478272
rect 219268 478214 226215 478216
rect 219268 478212 219274 478214
rect 226149 478211 226215 478214
rect 234061 478274 234127 478277
rect 374494 478274 374500 478276
rect 234061 478272 374500 478274
rect 234061 478216 234066 478272
rect 234122 478216 374500 478272
rect 234061 478214 374500 478216
rect 234061 478211 234127 478214
rect 374494 478212 374500 478214
rect 374564 478212 374570 478276
rect 49509 478138 49575 478141
rect 94037 478138 94103 478141
rect 49509 478136 94103 478138
rect 49509 478080 49514 478136
rect 49570 478080 94042 478136
rect 94098 478080 94103 478136
rect 49509 478078 94103 478080
rect 49509 478075 49575 478078
rect 94037 478075 94103 478078
rect 146017 478138 146083 478141
rect 200614 478138 200620 478140
rect 146017 478136 200620 478138
rect 146017 478080 146022 478136
rect 146078 478080 200620 478136
rect 146017 478078 200620 478080
rect 146017 478075 146083 478078
rect 200614 478076 200620 478078
rect 200684 478076 200690 478140
rect 234521 478138 234587 478141
rect 375966 478138 375972 478140
rect 234521 478136 375972 478138
rect 234521 478080 234526 478136
rect 234582 478080 375972 478136
rect 234521 478078 375972 478080
rect 234521 478075 234587 478078
rect 375966 478076 375972 478078
rect 376036 478076 376042 478140
rect 54702 477940 54708 478004
rect 54772 478002 54778 478004
rect 73797 478002 73863 478005
rect 54772 478000 73863 478002
rect 54772 477944 73802 478000
rect 73858 477944 73863 478000
rect 54772 477942 73863 477944
rect 54772 477940 54778 477942
rect 73797 477939 73863 477942
rect 179965 478002 180031 478005
rect 197353 478002 197419 478005
rect 198222 478002 198228 478004
rect 179965 478000 180810 478002
rect 179965 477944 179970 478000
rect 180026 477944 180810 478000
rect 179965 477942 180810 477944
rect 179965 477939 180031 477942
rect 50705 477732 50771 477733
rect 50654 477730 50660 477732
rect 50614 477670 50660 477730
rect 50724 477728 50771 477732
rect 50766 477672 50771 477728
rect 50654 477668 50660 477670
rect 50724 477668 50771 477672
rect 180750 477730 180810 477942
rect 197353 478000 198228 478002
rect 197353 477944 197358 478000
rect 197414 477944 198228 478000
rect 197353 477942 198228 477944
rect 197353 477939 197419 477942
rect 198222 477940 198228 477942
rect 198292 477940 198298 478004
rect 208393 478002 208459 478005
rect 209630 478002 209636 478004
rect 208393 478000 209636 478002
rect 208393 477944 208398 478000
rect 208454 477944 209636 478000
rect 208393 477942 209636 477944
rect 208393 477939 208459 477942
rect 209630 477940 209636 477942
rect 209700 477940 209706 478004
rect 197445 477866 197511 477869
rect 198590 477866 198596 477868
rect 197445 477864 198596 477866
rect 197445 477808 197450 477864
rect 197506 477808 198596 477864
rect 197445 477806 198596 477808
rect 197445 477803 197511 477806
rect 198590 477804 198596 477806
rect 198660 477804 198666 477868
rect 199326 477730 199332 477732
rect 180750 477670 199332 477730
rect 199326 477668 199332 477670
rect 199396 477668 199402 477732
rect 205633 477730 205699 477733
rect 206502 477730 206508 477732
rect 205633 477728 206508 477730
rect 205633 477672 205638 477728
rect 205694 477672 206508 477728
rect 205633 477670 206508 477672
rect 50705 477667 50771 477668
rect 205633 477667 205699 477670
rect 206502 477668 206508 477670
rect 206572 477668 206578 477732
rect 50889 477596 50955 477597
rect 50838 477594 50844 477596
rect 50798 477534 50844 477594
rect 50908 477592 50955 477596
rect 50950 477536 50955 477592
rect 50838 477532 50844 477534
rect 50908 477532 50955 477536
rect 50889 477531 50955 477532
rect 200481 477594 200547 477597
rect 216949 477596 217015 477597
rect 217409 477596 217475 477597
rect 200982 477594 200988 477596
rect 200481 477592 200988 477594
rect 200481 477536 200486 477592
rect 200542 477536 200988 477592
rect 200481 477534 200988 477536
rect 200481 477531 200547 477534
rect 200982 477532 200988 477534
rect 201052 477532 201058 477596
rect 216949 477594 216996 477596
rect 216904 477592 216996 477594
rect 216904 477536 216954 477592
rect 216904 477534 216996 477536
rect 216949 477532 216996 477534
rect 217060 477532 217066 477596
rect 217358 477594 217364 477596
rect 217318 477534 217364 477594
rect 217428 477592 217475 477596
rect 217470 477536 217475 477592
rect 217358 477532 217364 477534
rect 217428 477532 217475 477536
rect 217542 477532 217548 477596
rect 217612 477594 217618 477596
rect 217777 477594 217843 477597
rect 217612 477592 217843 477594
rect 217612 477536 217782 477592
rect 217838 477536 217843 477592
rect 217612 477534 217843 477536
rect 217612 477532 217618 477534
rect 216949 477531 217015 477532
rect 217409 477531 217475 477532
rect 217777 477531 217843 477534
rect 219934 477532 219940 477596
rect 220004 477594 220010 477596
rect 223113 477594 223179 477597
rect 220004 477592 223179 477594
rect 220004 477536 223118 477592
rect 223174 477536 223179 477592
rect 220004 477534 223179 477536
rect 220004 477532 220010 477534
rect 223113 477531 223179 477534
rect 154849 476914 154915 476917
rect 154849 476912 161490 476914
rect 154849 476856 154854 476912
rect 154910 476856 161490 476912
rect 154849 476854 161490 476856
rect 154849 476851 154915 476854
rect 161430 476778 161490 476854
rect 208342 476778 208348 476780
rect 161430 476718 208348 476778
rect 208342 476716 208348 476718
rect 208412 476716 208418 476780
rect 255681 476778 255747 476781
rect 377254 476778 377260 476780
rect 255681 476776 377260 476778
rect 255681 476720 255686 476776
rect 255742 476720 377260 476776
rect 255681 476718 377260 476720
rect 255681 476715 255747 476718
rect 377254 476716 377260 476718
rect 377324 476716 377330 476780
rect 58985 475962 59051 475965
rect 95785 475962 95851 475965
rect 58985 475960 95851 475962
rect 58985 475904 58990 475960
rect 59046 475904 95790 475960
rect 95846 475904 95851 475960
rect 58985 475902 95851 475904
rect 58985 475899 59051 475902
rect 95785 475899 95851 475902
rect -960 475540 480 475780
rect 57278 475764 57284 475828
rect 57348 475826 57354 475828
rect 121361 475826 121427 475829
rect 57348 475824 121427 475826
rect 57348 475768 121366 475824
rect 121422 475768 121427 475824
rect 57348 475766 121427 475768
rect 57348 475764 57354 475766
rect 121361 475763 121427 475766
rect 50429 475690 50495 475693
rect 120901 475690 120967 475693
rect 50429 475688 120967 475690
rect 50429 475632 50434 475688
rect 50490 475632 120906 475688
rect 120962 475632 120967 475688
rect 50429 475630 120967 475632
rect 50429 475627 50495 475630
rect 120901 475627 120967 475630
rect 148685 475690 148751 475693
rect 211654 475690 211660 475692
rect 148685 475688 211660 475690
rect 148685 475632 148690 475688
rect 148746 475632 211660 475688
rect 148685 475630 211660 475632
rect 148685 475627 148751 475630
rect 211654 475628 211660 475630
rect 211724 475628 211730 475692
rect 46749 475554 46815 475557
rect 120073 475554 120139 475557
rect 46749 475552 120139 475554
rect 46749 475496 46754 475552
rect 46810 475496 120078 475552
rect 120134 475496 120139 475552
rect 46749 475494 120139 475496
rect 46749 475491 46815 475494
rect 120073 475491 120139 475494
rect 146477 475554 146543 475557
rect 214414 475554 214420 475556
rect 146477 475552 214420 475554
rect 146477 475496 146482 475552
rect 146538 475496 214420 475552
rect 146477 475494 214420 475496
rect 146477 475491 146543 475494
rect 214414 475492 214420 475494
rect 214484 475492 214490 475556
rect 223573 475554 223639 475557
rect 223573 475552 229110 475554
rect 223573 475496 223578 475552
rect 223634 475496 229110 475552
rect 223573 475494 229110 475496
rect 223573 475491 223639 475494
rect 47894 475356 47900 475420
rect 47964 475418 47970 475420
rect 126605 475418 126671 475421
rect 47964 475416 126671 475418
rect 47964 475360 126610 475416
rect 126666 475360 126671 475416
rect 47964 475358 126671 475360
rect 47964 475356 47970 475358
rect 126605 475355 126671 475358
rect 145097 475418 145163 475421
rect 214598 475418 214604 475420
rect 145097 475416 214604 475418
rect 145097 475360 145102 475416
rect 145158 475360 214604 475416
rect 145097 475358 214604 475360
rect 145097 475355 145163 475358
rect 214598 475356 214604 475358
rect 214668 475356 214674 475420
rect 229050 475418 229110 475494
rect 378726 475418 378732 475420
rect 229050 475358 378732 475418
rect 378726 475356 378732 475358
rect 378796 475356 378802 475420
rect 146937 474330 147003 474333
rect 204846 474330 204852 474332
rect 146937 474328 204852 474330
rect 146937 474272 146942 474328
rect 146998 474272 204852 474328
rect 146937 474270 204852 474272
rect 146937 474267 147003 474270
rect 204846 474268 204852 474270
rect 204916 474268 204922 474332
rect 144729 474194 144795 474197
rect 205030 474194 205036 474196
rect 144729 474192 205036 474194
rect 144729 474136 144734 474192
rect 144790 474136 205036 474192
rect 144729 474134 205036 474136
rect 144729 474131 144795 474134
rect 205030 474132 205036 474134
rect 205100 474132 205106 474196
rect 152641 474058 152707 474061
rect 215334 474058 215340 474060
rect 152641 474056 215340 474058
rect 152641 474000 152646 474056
rect 152702 474000 215340 474056
rect 152641 473998 215340 474000
rect 152641 473995 152707 473998
rect 215334 473996 215340 473998
rect 215404 473996 215410 474060
rect 233693 474058 233759 474061
rect 378174 474058 378180 474060
rect 233693 474056 378180 474058
rect 233693 474000 233698 474056
rect 233754 474000 378180 474056
rect 233693 473998 378180 474000
rect 233693 473995 233759 473998
rect 378174 473996 378180 473998
rect 378244 473996 378250 474060
rect 158805 472834 158871 472837
rect 208894 472834 208900 472836
rect 158805 472832 208900 472834
rect 158805 472776 158810 472832
rect 158866 472776 208900 472832
rect 158805 472774 208900 472776
rect 158805 472771 158871 472774
rect 208894 472772 208900 472774
rect 208964 472772 208970 472836
rect 230105 472834 230171 472837
rect 358118 472834 358124 472836
rect 230105 472832 358124 472834
rect 230105 472776 230110 472832
rect 230166 472776 358124 472832
rect 230105 472774 358124 472776
rect 230105 472771 230171 472774
rect 358118 472772 358124 472774
rect 358188 472772 358194 472836
rect 43897 472698 43963 472701
rect 119153 472698 119219 472701
rect 43897 472696 119219 472698
rect 43897 472640 43902 472696
rect 43958 472640 119158 472696
rect 119214 472640 119219 472696
rect 43897 472638 119219 472640
rect 43897 472635 43963 472638
rect 119153 472635 119219 472638
rect 164509 472698 164575 472701
rect 214782 472698 214788 472700
rect 164509 472696 214788 472698
rect 164509 472640 164514 472696
rect 164570 472640 214788 472696
rect 164509 472638 214788 472640
rect 164509 472635 164575 472638
rect 214782 472636 214788 472638
rect 214852 472636 214858 472700
rect 232773 472698 232839 472701
rect 370446 472698 370452 472700
rect 232773 472696 370452 472698
rect 232773 472640 232778 472696
rect 232834 472640 370452 472696
rect 232773 472638 370452 472640
rect 232773 472635 232839 472638
rect 370446 472636 370452 472638
rect 370516 472636 370522 472700
rect 42609 472562 42675 472565
rect 123569 472562 123635 472565
rect 42609 472560 123635 472562
rect 42609 472504 42614 472560
rect 42670 472504 123574 472560
rect 123630 472504 123635 472560
rect 42609 472502 123635 472504
rect 42609 472499 42675 472502
rect 123569 472499 123635 472502
rect 153929 472562 153995 472565
rect 218830 472562 218836 472564
rect 153929 472560 218836 472562
rect 153929 472504 153934 472560
rect 153990 472504 218836 472560
rect 153929 472502 218836 472504
rect 153929 472499 153995 472502
rect 218830 472500 218836 472502
rect 218900 472500 218906 472564
rect 231853 472562 231919 472565
rect 376150 472562 376156 472564
rect 231853 472560 376156 472562
rect 231853 472504 231858 472560
rect 231914 472504 376156 472560
rect 231853 472502 376156 472504
rect 231853 472499 231919 472502
rect 376150 472500 376156 472502
rect 376220 472500 376226 472564
rect 149973 471610 150039 471613
rect 202270 471610 202276 471612
rect 149973 471608 202276 471610
rect 149973 471552 149978 471608
rect 150034 471552 202276 471608
rect 149973 471550 202276 471552
rect 149973 471547 150039 471550
rect 202270 471548 202276 471550
rect 202340 471548 202346 471612
rect 160277 471474 160343 471477
rect 214966 471474 214972 471476
rect 160277 471472 214972 471474
rect 160277 471416 160282 471472
rect 160338 471416 214972 471472
rect 160277 471414 214972 471416
rect 160277 471411 160343 471414
rect 214966 471412 214972 471414
rect 215036 471412 215042 471476
rect 145557 471338 145623 471341
rect 215886 471338 215892 471340
rect 145557 471336 215892 471338
rect 145557 471280 145562 471336
rect 145618 471280 215892 471336
rect 145557 471278 215892 471280
rect 145557 471275 145623 471278
rect 215886 471276 215892 471278
rect 215956 471276 215962 471340
rect 271137 471338 271203 471341
rect 359590 471338 359596 471340
rect 271137 471336 359596 471338
rect 271137 471280 271142 471336
rect 271198 471280 359596 471336
rect 271137 471278 359596 471280
rect 271137 471275 271203 471278
rect 359590 471276 359596 471278
rect 359660 471276 359666 471340
rect 583520 471324 584960 471564
rect 61469 471202 61535 471205
rect 199142 471202 199148 471204
rect 61469 471200 199148 471202
rect 61469 471144 61474 471200
rect 61530 471144 199148 471200
rect 61469 471142 199148 471144
rect 61469 471139 61535 471142
rect 199142 471140 199148 471142
rect 199212 471140 199218 471204
rect 231025 471202 231091 471205
rect 378910 471202 378916 471204
rect 231025 471200 378916 471202
rect 231025 471144 231030 471200
rect 231086 471144 378916 471200
rect 231025 471142 378916 471144
rect 231025 471139 231091 471142
rect 378910 471140 378916 471142
rect 378980 471140 378986 471204
rect 45277 469978 45343 469981
rect 125869 469978 125935 469981
rect 45277 469976 125935 469978
rect 45277 469920 45282 469976
rect 45338 469920 125874 469976
rect 125930 469920 125935 469976
rect 45277 469918 125935 469920
rect 45277 469915 45343 469918
rect 125869 469915 125935 469918
rect 156045 469978 156111 469981
rect 209814 469978 209820 469980
rect 156045 469976 209820 469978
rect 156045 469920 156050 469976
rect 156106 469920 209820 469976
rect 156045 469918 209820 469920
rect 156045 469915 156111 469918
rect 209814 469916 209820 469918
rect 209884 469916 209890 469980
rect 280245 469978 280311 469981
rect 377438 469978 377444 469980
rect 280245 469976 377444 469978
rect 280245 469920 280250 469976
rect 280306 469920 377444 469976
rect 280245 469918 377444 469920
rect 280245 469915 280311 469918
rect 377438 469916 377444 469918
rect 377508 469916 377514 469980
rect 43437 469842 43503 469845
rect 125777 469842 125843 469845
rect 43437 469840 125843 469842
rect 43437 469784 43442 469840
rect 43498 469784 125782 469840
rect 125838 469784 125843 469840
rect 43437 469782 125843 469784
rect 43437 469779 43503 469782
rect 125777 469779 125843 469782
rect 150525 469842 150591 469845
rect 212758 469842 212764 469844
rect 150525 469840 212764 469842
rect 150525 469784 150530 469840
rect 150586 469784 212764 469840
rect 150525 469782 212764 469784
rect 150525 469779 150591 469782
rect 212758 469780 212764 469782
rect 212828 469780 212834 469844
rect 223665 469842 223731 469845
rect 379094 469842 379100 469844
rect 223665 469840 379100 469842
rect 223665 469784 223670 469840
rect 223726 469784 379100 469840
rect 223665 469782 379100 469784
rect 223665 469779 223731 469782
rect 379094 469780 379100 469782
rect 379164 469780 379170 469844
rect 263685 468754 263751 468757
rect 359406 468754 359412 468756
rect 263685 468752 359412 468754
rect 263685 468696 263690 468752
rect 263746 468696 359412 468752
rect 263685 468694 359412 468696
rect 263685 468691 263751 468694
rect 359406 468692 359412 468694
rect 359476 468692 359482 468756
rect 155953 468618 156019 468621
rect 212574 468618 212580 468620
rect 155953 468616 212580 468618
rect 155953 468560 155958 468616
rect 156014 468560 212580 468616
rect 155953 468558 212580 468560
rect 155953 468555 156019 468558
rect 212574 468556 212580 468558
rect 212644 468556 212650 468620
rect 255313 468618 255379 468621
rect 379462 468618 379468 468620
rect 255313 468616 379468 468618
rect 255313 468560 255318 468616
rect 255374 468560 379468 468616
rect 255313 468558 379468 468560
rect 255313 468555 255379 468558
rect 379462 468556 379468 468558
rect 379532 468556 379538 468620
rect 127065 468482 127131 468485
rect 196750 468482 196756 468484
rect 127065 468480 196756 468482
rect 127065 468424 127070 468480
rect 127126 468424 196756 468480
rect 127065 468422 196756 468424
rect 127065 468419 127131 468422
rect 196750 468420 196756 468422
rect 196820 468420 196826 468484
rect 234613 468482 234679 468485
rect 362902 468482 362908 468484
rect 234613 468480 362908 468482
rect 234613 468424 234618 468480
rect 234674 468424 362908 468480
rect 234613 468422 362908 468424
rect 234613 468419 234679 468422
rect 362902 468420 362908 468422
rect 362972 468420 362978 468484
rect 160185 467258 160251 467261
rect 203190 467258 203196 467260
rect 160185 467256 203196 467258
rect 160185 467200 160190 467256
rect 160246 467200 203196 467256
rect 160185 467198 203196 467200
rect 160185 467195 160251 467198
rect 203190 467196 203196 467198
rect 203260 467196 203266 467260
rect 157425 467122 157491 467125
rect 207054 467122 207060 467124
rect 157425 467120 207060 467122
rect 157425 467064 157430 467120
rect 157486 467064 207060 467120
rect 157425 467062 207060 467064
rect 157425 467059 157491 467062
rect 207054 467060 207060 467062
rect 207124 467060 207130 467124
rect 59077 466442 59143 466445
rect 89805 466442 89871 466445
rect 59077 466440 89871 466442
rect 59077 466384 59082 466440
rect 59138 466384 89810 466440
rect 89866 466384 89871 466440
rect 59077 466382 89871 466384
rect 59077 466379 59143 466382
rect 89805 466379 89871 466382
rect 59169 466306 59235 466309
rect 91277 466306 91343 466309
rect 59169 466304 91343 466306
rect 59169 466248 59174 466304
rect 59230 466248 91282 466304
rect 91338 466248 91343 466304
rect 59169 466246 91343 466248
rect 59169 466243 59235 466246
rect 91277 466243 91343 466246
rect 183553 466306 183619 466309
rect 217174 466306 217180 466308
rect 183553 466304 217180 466306
rect 183553 466248 183558 466304
rect 183614 466248 217180 466304
rect 183553 466246 217180 466248
rect 183553 466243 183619 466246
rect 217174 466244 217180 466246
rect 217244 466244 217250 466308
rect 53557 466170 53623 466173
rect 85757 466170 85823 466173
rect 53557 466168 85823 466170
rect 53557 466112 53562 466168
rect 53618 466112 85762 466168
rect 85818 466112 85823 466168
rect 53557 466110 85823 466112
rect 53557 466107 53623 466110
rect 85757 466107 85823 466110
rect 169845 466170 169911 466173
rect 204897 466170 204963 466173
rect 169845 466168 204963 466170
rect 169845 466112 169850 466168
rect 169906 466112 204902 466168
rect 204958 466112 204963 466168
rect 169845 466110 204963 466112
rect 169845 466107 169911 466110
rect 204897 466107 204963 466110
rect 59905 466034 59971 466037
rect 92657 466034 92723 466037
rect 59905 466032 92723 466034
rect 59905 465976 59910 466032
rect 59966 465976 92662 466032
rect 92718 465976 92723 466032
rect 59905 465974 92723 465976
rect 59905 465971 59971 465974
rect 92657 465971 92723 465974
rect 161657 466034 161723 466037
rect 205081 466034 205147 466037
rect 161657 466032 205147 466034
rect 161657 465976 161662 466032
rect 161718 465976 205086 466032
rect 205142 465976 205147 466032
rect 161657 465974 205147 465976
rect 161657 465971 161723 465974
rect 205081 465971 205147 465974
rect 50705 465898 50771 465901
rect 84285 465898 84351 465901
rect 50705 465896 84351 465898
rect 50705 465840 50710 465896
rect 50766 465840 84290 465896
rect 84346 465840 84351 465896
rect 50705 465838 84351 465840
rect 50705 465835 50771 465838
rect 84285 465835 84351 465838
rect 162853 465898 162919 465901
rect 206461 465898 206527 465901
rect 162853 465896 206527 465898
rect 162853 465840 162858 465896
rect 162914 465840 206466 465896
rect 206522 465840 206527 465896
rect 162853 465838 206527 465840
rect 162853 465835 162919 465838
rect 206461 465835 206527 465838
rect 287237 465898 287303 465901
rect 359958 465898 359964 465900
rect 287237 465896 359964 465898
rect 287237 465840 287242 465896
rect 287298 465840 359964 465896
rect 287237 465838 359964 465840
rect 287237 465835 287303 465838
rect 359958 465836 359964 465838
rect 360028 465836 360034 465900
rect 55438 465700 55444 465764
rect 55508 465762 55514 465764
rect 89897 465762 89963 465765
rect 55508 465760 89963 465762
rect 55508 465704 89902 465760
rect 89958 465704 89963 465760
rect 55508 465702 89963 465704
rect 55508 465700 55514 465702
rect 89897 465699 89963 465702
rect 167085 465762 167151 465765
rect 218881 465762 218947 465765
rect 167085 465760 218947 465762
rect 167085 465704 167090 465760
rect 167146 465704 218886 465760
rect 218942 465704 218947 465760
rect 167085 465702 218947 465704
rect 167085 465699 167151 465702
rect 218881 465699 218947 465702
rect 229093 465762 229159 465765
rect 364926 465762 364932 465764
rect 229093 465760 364932 465762
rect 229093 465704 229098 465760
rect 229154 465704 364932 465760
rect 229093 465702 364932 465704
rect 229093 465699 229159 465702
rect 364926 465700 364932 465702
rect 364996 465700 365002 465764
rect 296713 464402 296779 464405
rect 376886 464402 376892 464404
rect 296713 464400 376892 464402
rect 296713 464344 296718 464400
rect 296774 464344 376892 464400
rect 296713 464342 376892 464344
rect 296713 464339 296779 464342
rect 376886 464340 376892 464342
rect 376956 464340 376962 464404
rect 52310 463388 52316 463452
rect 52380 463450 52386 463452
rect 70485 463450 70551 463453
rect 52380 463448 70551 463450
rect 52380 463392 70490 463448
rect 70546 463392 70551 463448
rect 52380 463390 70551 463392
rect 52380 463388 52386 463390
rect 70485 463387 70551 463390
rect 169937 463450 170003 463453
rect 203006 463450 203012 463452
rect 169937 463448 203012 463450
rect 169937 463392 169942 463448
rect 169998 463392 203012 463448
rect 169937 463390 203012 463392
rect 169937 463387 170003 463390
rect 203006 463388 203012 463390
rect 203076 463388 203082 463452
rect 50889 463314 50955 463317
rect 71957 463314 72023 463317
rect 50889 463312 72023 463314
rect 50889 463256 50894 463312
rect 50950 463256 71962 463312
rect 72018 463256 72023 463312
rect 50889 463254 72023 463256
rect 50889 463251 50955 463254
rect 71957 463251 72023 463254
rect 169753 463314 169819 463317
rect 211889 463314 211955 463317
rect 169753 463312 211955 463314
rect 169753 463256 169758 463312
rect 169814 463256 211894 463312
rect 211950 463256 211955 463312
rect 169753 463254 211955 463256
rect 169753 463251 169819 463254
rect 211889 463251 211955 463254
rect 48078 463116 48084 463180
rect 48148 463178 48154 463180
rect 69197 463178 69263 463181
rect 48148 463176 69263 463178
rect 48148 463120 69202 463176
rect 69258 463120 69263 463176
rect 48148 463118 69263 463120
rect 48148 463116 48154 463118
rect 69197 463115 69263 463118
rect 154665 463178 154731 463181
rect 204294 463178 204300 463180
rect 154665 463176 204300 463178
rect 154665 463120 154670 463176
rect 154726 463120 204300 463176
rect 154665 463118 204300 463120
rect 154665 463115 154731 463118
rect 204294 463116 204300 463118
rect 204364 463116 204370 463180
rect 50470 462980 50476 463044
rect 50540 463042 50546 463044
rect 80145 463042 80211 463045
rect 50540 463040 80211 463042
rect 50540 462984 80150 463040
rect 80206 462984 80211 463040
rect 50540 462982 80211 462984
rect 50540 462980 50546 462982
rect 80145 462979 80211 462982
rect 147673 463042 147739 463045
rect 218697 463042 218763 463045
rect 147673 463040 218763 463042
rect 147673 462984 147678 463040
rect 147734 462984 218702 463040
rect 218758 462984 218763 463040
rect 147673 462982 218763 462984
rect 147673 462979 147739 462982
rect 218697 462979 218763 462982
rect 277485 463042 277551 463045
rect 359774 463042 359780 463044
rect 277485 463040 359780 463042
rect 277485 462984 277490 463040
rect 277546 462984 359780 463040
rect 277485 462982 359780 462984
rect 277485 462979 277551 462982
rect 359774 462980 359780 462982
rect 359844 462980 359850 463044
rect 50613 462906 50679 462909
rect 93853 462906 93919 462909
rect 50613 462904 93919 462906
rect 50613 462848 50618 462904
rect 50674 462848 93858 462904
rect 93914 462848 93919 462904
rect 50613 462846 93919 462848
rect 50613 462843 50679 462846
rect 93853 462843 93919 462846
rect 107745 462906 107811 462909
rect 198958 462906 198964 462908
rect 107745 462904 198964 462906
rect 107745 462848 107750 462904
rect 107806 462848 198964 462904
rect 107745 462846 198964 462848
rect 107745 462843 107811 462846
rect 198958 462844 198964 462846
rect 199028 462844 199034 462908
rect 276105 462906 276171 462909
rect 377622 462906 377628 462908
rect 276105 462904 377628 462906
rect 276105 462848 276110 462904
rect 276166 462848 377628 462904
rect 276105 462846 377628 462848
rect 276105 462843 276171 462846
rect 377622 462844 377628 462846
rect 377692 462844 377698 462908
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 510838 462164 510844 462228
rect 510908 462226 510914 462228
rect 511257 462226 511323 462229
rect 510908 462224 511323 462226
rect 510908 462168 511262 462224
rect 511318 462168 511323 462224
rect 510908 462166 511323 462168
rect 510908 462164 510914 462166
rect 511257 462163 511323 462166
rect 179597 461684 179663 461685
rect 179597 461680 179644 461684
rect 179708 461682 179714 461684
rect 179597 461624 179602 461680
rect 179597 461620 179644 461624
rect 179708 461622 179754 461682
rect 179708 461620 179714 461622
rect 179597 461619 179663 461620
rect 58566 461484 58572 461548
rect 58636 461546 58642 461548
rect 73337 461546 73403 461549
rect 58636 461544 73403 461546
rect 58636 461488 73342 461544
rect 73398 461488 73403 461544
rect 58636 461486 73403 461488
rect 58636 461484 58642 461486
rect 73337 461483 73403 461486
rect 172605 461546 172671 461549
rect 200798 461546 200804 461548
rect 172605 461544 200804 461546
rect 172605 461488 172610 461544
rect 172666 461488 200804 461544
rect 172605 461486 200804 461488
rect 172605 461483 172671 461486
rect 200798 461484 200804 461486
rect 200868 461484 200874 461548
rect 178309 461412 178375 461413
rect 178309 461408 178356 461412
rect 178420 461410 178426 461412
rect 178309 461352 178314 461408
rect 178309 461348 178356 461352
rect 178420 461350 178466 461410
rect 178420 461348 178426 461350
rect 178309 461347 178375 461348
rect 190913 461004 190979 461005
rect 338297 461004 338363 461005
rect 339769 461004 339835 461005
rect 350993 461004 351059 461005
rect 190862 461002 190868 461004
rect 190822 460942 190868 461002
rect 190932 461000 190979 461004
rect 338246 461002 338252 461004
rect 190974 460944 190979 461000
rect 190862 460940 190868 460942
rect 190932 460940 190979 460944
rect 338206 460942 338252 461002
rect 338316 461000 338363 461004
rect 339718 461002 339724 461004
rect 338358 460944 338363 461000
rect 338246 460940 338252 460942
rect 338316 460940 338363 460944
rect 339678 460942 339724 461002
rect 339788 461000 339835 461004
rect 350942 461002 350948 461004
rect 339830 460944 339835 461000
rect 339718 460940 339724 460942
rect 339788 460940 339835 460944
rect 350902 460942 350948 461002
rect 351012 461000 351059 461004
rect 351054 460944 351059 461000
rect 350942 460940 350948 460942
rect 351012 460940 351059 460944
rect 190913 460939 190979 460940
rect 338297 460939 338363 460940
rect 339769 460939 339835 460940
rect 350993 460939 351059 460940
rect 498377 461002 498443 461005
rect 499849 461004 499915 461005
rect 498510 461002 498516 461004
rect 498377 461000 498516 461002
rect 498377 460944 498382 461000
rect 498438 460944 498516 461000
rect 498377 460942 498516 460944
rect 498377 460939 498443 460942
rect 498510 460940 498516 460942
rect 498580 460940 498586 461004
rect 499798 461002 499804 461004
rect 499758 460942 499804 461002
rect 499868 461000 499915 461004
rect 499910 460944 499915 461000
rect 499798 460940 499804 460942
rect 499868 460940 499915 460944
rect 499849 460939 499915 460940
rect 55070 460804 55076 460868
rect 55140 460866 55146 460868
rect 71773 460866 71839 460869
rect 55140 460864 71839 460866
rect 55140 460808 71778 460864
rect 71834 460808 71839 460864
rect 55140 460806 71839 460808
rect 55140 460804 55146 460806
rect 71773 460803 71839 460806
rect 171225 460866 171291 460869
rect 206318 460866 206324 460868
rect 171225 460864 206324 460866
rect 171225 460808 171230 460864
rect 171286 460808 206324 460864
rect 171225 460806 206324 460808
rect 171225 460803 171291 460806
rect 206318 460804 206324 460806
rect 206388 460804 206394 460868
rect 54886 460668 54892 460732
rect 54956 460730 54962 460732
rect 75913 460730 75979 460733
rect 54956 460728 75979 460730
rect 54956 460672 75918 460728
rect 75974 460672 75979 460728
rect 54956 460670 75979 460672
rect 54956 460668 54962 460670
rect 75913 460667 75979 460670
rect 166993 460730 167059 460733
rect 210366 460730 210372 460732
rect 166993 460728 210372 460730
rect 166993 460672 166998 460728
rect 167054 460672 210372 460728
rect 166993 460670 210372 460672
rect 166993 460667 167059 460670
rect 210366 460668 210372 460670
rect 210436 460668 210442 460732
rect 53414 460532 53420 460596
rect 53484 460594 53490 460596
rect 74717 460594 74783 460597
rect 53484 460592 74783 460594
rect 53484 460536 74722 460592
rect 74778 460536 74783 460592
rect 53484 460534 74783 460536
rect 53484 460532 53490 460534
rect 74717 460531 74783 460534
rect 165613 460594 165679 460597
rect 213126 460594 213132 460596
rect 165613 460592 213132 460594
rect 165613 460536 165618 460592
rect 165674 460536 213132 460592
rect 165613 460534 213132 460536
rect 165613 460531 165679 460534
rect 213126 460532 213132 460534
rect 213196 460532 213202 460596
rect 46606 460396 46612 460460
rect 46676 460458 46682 460460
rect 69105 460458 69171 460461
rect 46676 460456 69171 460458
rect 46676 460400 69110 460456
rect 69166 460400 69171 460456
rect 46676 460398 69171 460400
rect 46676 460396 46682 460398
rect 69105 460395 69171 460398
rect 154573 460458 154639 460461
rect 205214 460458 205220 460460
rect 154573 460456 205220 460458
rect 154573 460400 154578 460456
rect 154634 460400 205220 460456
rect 154573 460398 205220 460400
rect 154573 460395 154639 460398
rect 205214 460396 205220 460398
rect 205284 460396 205290 460460
rect 51942 460260 51948 460324
rect 52012 460322 52018 460324
rect 74625 460322 74691 460325
rect 52012 460320 74691 460322
rect 52012 460264 74630 460320
rect 74686 460264 74691 460320
rect 52012 460262 74691 460264
rect 52012 460260 52018 460262
rect 74625 460259 74691 460262
rect 143533 460322 143599 460325
rect 206134 460322 206140 460324
rect 143533 460320 206140 460322
rect 143533 460264 143538 460320
rect 143594 460264 206140 460320
rect 143533 460262 206140 460264
rect 143533 460259 143599 460262
rect 206134 460260 206140 460262
rect 206204 460260 206210 460324
rect 44950 460124 44956 460188
rect 45020 460186 45026 460188
rect 67817 460186 67883 460189
rect 45020 460184 67883 460186
rect 45020 460128 67822 460184
rect 67878 460128 67883 460184
rect 45020 460126 67883 460128
rect 45020 460124 45026 460126
rect 67817 460123 67883 460126
rect 150433 460186 150499 460189
rect 215518 460186 215524 460188
rect 150433 460184 215524 460186
rect 150433 460128 150438 460184
rect 150494 460128 215524 460184
rect 150433 460126 215524 460128
rect 150433 460123 150499 460126
rect 215518 460124 215524 460126
rect 215588 460124 215594 460188
rect 59118 459988 59124 460052
rect 59188 460050 59194 460052
rect 67725 460050 67791 460053
rect 59188 460048 67791 460050
rect 59188 459992 67730 460048
rect 67786 459992 67791 460048
rect 59188 459990 67791 459992
rect 59188 459988 59194 459990
rect 67725 459987 67791 459990
rect 182817 460050 182883 460053
rect 198774 460050 198780 460052
rect 182817 460048 198780 460050
rect 182817 459992 182822 460048
rect 182878 459992 198780 460048
rect 182817 459990 198780 459992
rect 182817 459987 182883 459990
rect 198774 459988 198780 459990
rect 198844 459988 198850 460052
rect 218329 459778 218395 459781
rect 218646 459778 218652 459780
rect 218329 459776 218652 459778
rect 218329 459720 218334 459776
rect 218390 459720 218652 459776
rect 218329 459718 218652 459720
rect 218329 459715 218395 459718
rect 218646 459716 218652 459718
rect 218716 459716 218722 459780
rect 48681 459644 48747 459645
rect 51625 459644 51691 459645
rect 48630 459642 48636 459644
rect 48590 459582 48636 459642
rect 48700 459640 48747 459644
rect 51574 459642 51580 459644
rect 48742 459584 48747 459640
rect 48630 459580 48636 459582
rect 48700 459580 48747 459584
rect 51534 459582 51580 459642
rect 51644 459640 51691 459644
rect 51686 459584 51691 459640
rect 51574 459580 51580 459582
rect 51644 459580 51691 459584
rect 52126 459580 52132 459644
rect 52196 459642 52202 459644
rect 52361 459642 52427 459645
rect 52196 459640 52427 459642
rect 52196 459584 52366 459640
rect 52422 459584 52427 459640
rect 52196 459582 52427 459584
rect 52196 459580 52202 459582
rect 48681 459579 48747 459580
rect 51625 459579 51691 459580
rect 52361 459579 52427 459582
rect 53373 459642 53439 459645
rect 53598 459642 53604 459644
rect 53373 459640 53604 459642
rect 53373 459584 53378 459640
rect 53434 459584 53604 459640
rect 53373 459582 53604 459584
rect 53373 459579 53439 459582
rect 53598 459580 53604 459582
rect 53668 459580 53674 459644
rect 55622 459580 55628 459644
rect 55692 459642 55698 459644
rect 55949 459642 56015 459645
rect 55692 459640 56015 459642
rect 55692 459584 55954 459640
rect 56010 459584 56015 459640
rect 55692 459582 56015 459584
rect 55692 459580 55698 459582
rect 55949 459579 56015 459582
rect 171317 459370 171383 459373
rect 202229 459370 202295 459373
rect 171317 459368 202295 459370
rect 171317 459312 171322 459368
rect 171378 459312 202234 459368
rect 202290 459312 202295 459368
rect 171317 459310 202295 459312
rect 171317 459307 171383 459310
rect 202229 459307 202295 459310
rect 172513 459234 172579 459237
rect 207749 459234 207815 459237
rect 172513 459232 207815 459234
rect 172513 459176 172518 459232
rect 172574 459176 207754 459232
rect 207810 459176 207815 459232
rect 172513 459174 207815 459176
rect 172513 459171 172579 459174
rect 207749 459171 207815 459174
rect 58934 459036 58940 459100
rect 59004 459098 59010 459100
rect 67633 459098 67699 459101
rect 59004 459096 67699 459098
rect 59004 459040 67638 459096
rect 67694 459040 67699 459096
rect 59004 459038 67699 459040
rect 59004 459036 59010 459038
rect 67633 459035 67699 459038
rect 171133 459098 171199 459101
rect 207974 459098 207980 459100
rect 171133 459096 207980 459098
rect 171133 459040 171138 459096
rect 171194 459040 207980 459096
rect 171133 459038 207980 459040
rect 171133 459035 171199 459038
rect 207974 459036 207980 459038
rect 208044 459036 208050 459100
rect 58750 458900 58756 458964
rect 58820 458962 58826 458964
rect 69013 458962 69079 458965
rect 58820 458960 69079 458962
rect 58820 458904 69018 458960
rect 69074 458904 69079 458960
rect 58820 458902 69079 458904
rect 58820 458900 58826 458902
rect 69013 458899 69079 458902
rect 164233 458962 164299 458965
rect 210509 458962 210575 458965
rect 164233 458960 210575 458962
rect 164233 458904 164238 458960
rect 164294 458904 210514 458960
rect 210570 458904 210575 458960
rect 164233 458902 210575 458904
rect 164233 458899 164299 458902
rect 210509 458899 210575 458902
rect 57830 458764 57836 458828
rect 57900 458826 57906 458828
rect 80237 458826 80303 458829
rect 57900 458824 80303 458826
rect 57900 458768 80242 458824
rect 80298 458768 80303 458824
rect 57900 458766 80303 458768
rect 57900 458764 57906 458766
rect 80237 458763 80303 458766
rect 161473 458826 161539 458829
rect 213361 458826 213427 458829
rect 161473 458824 213427 458826
rect 161473 458768 161478 458824
rect 161534 458768 213366 458824
rect 213422 458768 213427 458824
rect 161473 458766 213427 458768
rect 161473 458763 161539 458766
rect 213361 458763 213427 458766
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect 199009 454746 199075 454749
rect 358905 454746 358971 454749
rect 516593 454746 516659 454749
rect 196558 454744 199075 454746
rect 196558 454688 199014 454744
rect 199070 454688 199075 454744
rect 196558 454686 199075 454688
rect 196558 454190 196618 454686
rect 199009 454683 199075 454686
rect 356562 454744 358971 454746
rect 356562 454688 358910 454744
rect 358966 454688 358971 454744
rect 356562 454686 358971 454688
rect 356562 454190 356622 454686
rect 358905 454683 358971 454686
rect 516558 454744 516659 454746
rect 516558 454688 516598 454744
rect 516654 454688 516659 454744
rect 516558 454683 516659 454688
rect 516558 454202 516618 454683
rect 518893 454202 518959 454205
rect 516558 454200 518959 454202
rect 516558 454144 518898 454200
rect 518954 454144 518959 454200
rect 516558 454142 518959 454144
rect 518893 454139 518959 454142
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect 56961 412314 57027 412317
rect 56961 412312 60062 412314
rect 56961 412256 56966 412312
rect 57022 412256 60062 412312
rect 56961 412254 60062 412256
rect 56961 412251 57027 412254
rect 60002 411894 60062 412254
rect 217777 411906 217843 411909
rect 219390 411906 220064 411924
rect 217777 411904 220064 411906
rect 217777 411848 217782 411904
rect 217838 411864 220064 411904
rect 377581 411906 377647 411909
rect 379470 411906 380052 411924
rect 377581 411904 380052 411906
rect 217838 411848 219450 411864
rect 217777 411846 219450 411848
rect 377581 411848 377586 411904
rect 377642 411864 380052 411904
rect 377642 411848 379530 411864
rect 377581 411846 379530 411848
rect 217777 411843 217843 411846
rect 377581 411843 377647 411846
rect 217685 410954 217751 410957
rect 219390 410954 220064 410972
rect 217685 410952 220064 410954
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 57053 410410 57119 410413
rect 60002 410410 60062 410942
rect 217685 410896 217690 410952
rect 217746 410912 220064 410952
rect 377489 410954 377555 410957
rect 379470 410954 380052 410972
rect 377489 410952 380052 410954
rect 217746 410896 219450 410912
rect 217685 410894 219450 410896
rect 377489 410896 377494 410952
rect 377550 410912 380052 410952
rect 377550 410896 379530 410912
rect 377489 410894 379530 410896
rect 217685 410891 217751 410894
rect 377489 410891 377555 410894
rect 57053 410408 60062 410410
rect 57053 410352 57058 410408
rect 57114 410352 60062 410408
rect 57053 410350 60062 410352
rect 57053 410347 57119 410350
rect 216765 408778 216831 408781
rect 219390 408778 220064 408796
rect 216765 408776 220064 408778
rect 57053 408642 57119 408645
rect 60002 408642 60062 408766
rect 216765 408720 216770 408776
rect 216826 408736 220064 408776
rect 377029 408778 377095 408781
rect 377305 408778 377371 408781
rect 379470 408778 380052 408796
rect 377029 408776 380052 408778
rect 216826 408720 219450 408736
rect 216765 408718 219450 408720
rect 377029 408720 377034 408776
rect 377090 408720 377310 408776
rect 377366 408736 380052 408776
rect 377366 408720 379530 408736
rect 377029 408718 379530 408720
rect 216765 408715 216831 408718
rect 377029 408715 377095 408718
rect 377305 408715 377371 408718
rect 57053 408640 60062 408642
rect 57053 408584 57058 408640
rect 57114 408584 60062 408640
rect 57053 408582 60062 408584
rect 57053 408579 57119 408582
rect 206686 408580 206692 408644
rect 206756 408642 206762 408644
rect 206921 408642 206987 408645
rect 206756 408640 206987 408642
rect 206756 408584 206926 408640
rect 206982 408584 206987 408640
rect 206756 408582 206987 408584
rect 206756 408580 206762 408582
rect 206921 408579 206987 408582
rect 360142 408580 360148 408644
rect 360212 408642 360218 408644
rect 361481 408642 361547 408645
rect 360212 408640 361547 408642
rect 360212 408584 361486 408640
rect 361542 408584 361547 408640
rect 360212 408582 361547 408584
rect 360212 408580 360218 408582
rect 361481 408579 361547 408582
rect 217869 407826 217935 407829
rect 219390 407826 220064 407844
rect 217869 407824 220064 407826
rect 56961 407418 57027 407421
rect 60002 407418 60062 407814
rect 217869 407768 217874 407824
rect 217930 407784 220064 407824
rect 376937 407826 377003 407829
rect 379470 407826 380052 407844
rect 376937 407824 380052 407826
rect 217930 407768 219450 407784
rect 217869 407766 219450 407768
rect 376937 407768 376942 407824
rect 376998 407784 380052 407824
rect 376998 407768 379530 407784
rect 376937 407766 379530 407768
rect 217869 407763 217935 407766
rect 376937 407763 377003 407766
rect 56961 407416 60062 407418
rect 56961 407360 56966 407416
rect 57022 407360 60062 407416
rect 56961 407358 60062 407360
rect 56961 407355 57027 407358
rect 217593 406058 217659 406061
rect 219390 406058 220064 406076
rect 217593 406056 220064 406058
rect 57053 405786 57119 405789
rect 60002 405786 60062 406046
rect 217593 406000 217598 406056
rect 217654 406016 220064 406056
rect 377213 406058 377279 406061
rect 377673 406058 377739 406061
rect 379470 406058 380052 406076
rect 377213 406056 380052 406058
rect 217654 406000 219450 406016
rect 217593 405998 219450 406000
rect 377213 406000 377218 406056
rect 377274 406000 377678 406056
rect 377734 406016 380052 406056
rect 377734 406000 379530 406016
rect 377213 405998 379530 406000
rect 217593 405995 217659 405998
rect 377213 405995 377279 405998
rect 377673 405995 377739 405998
rect 57053 405784 60062 405786
rect 57053 405728 57058 405784
rect 57114 405728 60062 405784
rect 57053 405726 60062 405728
rect 57053 405723 57119 405726
rect 216857 404970 216923 404973
rect 219390 404970 220064 404988
rect 216857 404968 220064 404970
rect 57053 404426 57119 404429
rect 60002 404426 60062 404958
rect 216857 404912 216862 404968
rect 216918 404928 220064 404968
rect 377305 404970 377371 404973
rect 379470 404970 380052 404988
rect 377305 404968 380052 404970
rect 216918 404912 219450 404928
rect 216857 404910 219450 404912
rect 377305 404912 377310 404968
rect 377366 404928 380052 404968
rect 580257 404970 580323 404973
rect 583520 404970 584960 405060
rect 580257 404968 584960 404970
rect 377366 404912 379530 404928
rect 377305 404910 379530 404912
rect 580257 404912 580262 404968
rect 580318 404912 584960 404968
rect 580257 404910 584960 404912
rect 216857 404907 216923 404910
rect 377305 404907 377371 404910
rect 580257 404907 580323 404910
rect 583520 404820 584960 404910
rect 57053 404424 60062 404426
rect 57053 404368 57058 404424
rect 57114 404368 60062 404424
rect 57053 404366 60062 404368
rect 57053 404363 57119 404366
rect 217317 403202 217383 403205
rect 219390 403202 220064 403220
rect 217317 403200 220064 403202
rect 57053 403066 57119 403069
rect 60002 403066 60062 403190
rect 217317 403144 217322 403200
rect 217378 403160 220064 403200
rect 377765 403202 377831 403205
rect 379470 403202 380052 403220
rect 377765 403200 380052 403202
rect 217378 403144 219450 403160
rect 217317 403142 219450 403144
rect 377765 403144 377770 403200
rect 377826 403160 380052 403200
rect 377826 403144 379530 403160
rect 377765 403142 379530 403144
rect 217317 403139 217383 403142
rect 377765 403139 377831 403142
rect 57053 403064 60062 403066
rect 57053 403008 57058 403064
rect 57114 403008 60062 403064
rect 57053 403006 60062 403008
rect 57053 403003 57119 403006
rect -960 397340 480 397580
rect 196558 393818 196618 394350
rect 199653 393818 199719 393821
rect 196558 393816 199719 393818
rect 196558 393760 199658 393816
rect 199714 393760 199719 393816
rect 196558 393758 199719 393760
rect 356562 393818 356622 394350
rect 358997 393818 359063 393821
rect 356562 393816 359063 393818
rect 356562 393760 359002 393816
rect 359058 393760 359063 393816
rect 356562 393758 359063 393760
rect 516558 393818 516618 394350
rect 518985 393818 519051 393821
rect 516558 393816 519051 393818
rect 516558 393760 518990 393816
rect 519046 393760 519051 393816
rect 516558 393758 519051 393760
rect 199653 393755 199719 393758
rect 358997 393755 359063 393758
rect 518985 393755 519051 393758
rect 199142 392730 199148 392732
rect 196558 392670 199148 392730
rect 199142 392668 199148 392670
rect 199212 392668 199218 392732
rect 356562 392186 356622 392718
rect 359089 392186 359155 392189
rect 356562 392184 359155 392186
rect 356562 392128 359094 392184
rect 359150 392128 359155 392184
rect 356562 392126 359155 392128
rect 516558 392186 516618 392718
rect 519353 392186 519419 392189
rect 516558 392184 519419 392186
rect 516558 392128 519358 392184
rect 519414 392128 519419 392184
rect 516558 392126 519419 392128
rect 359089 392123 359155 392126
rect 519353 392123 519419 392126
rect 199142 391988 199148 392052
rect 199212 392050 199218 392052
rect 199510 392050 199516 392052
rect 199212 391990 199516 392050
rect 199212 391988 199218 391990
rect 199510 391988 199516 391990
rect 199580 391988 199586 392052
rect 583520 391628 584960 391868
rect 196558 390826 196618 391358
rect 199193 390826 199259 390829
rect 196558 390824 199259 390826
rect 196558 390768 199198 390824
rect 199254 390768 199259 390824
rect 196558 390766 199259 390768
rect 356562 390826 356622 391358
rect 359733 390826 359799 390829
rect 356562 390824 359799 390826
rect 356562 390768 359738 390824
rect 359794 390768 359799 390824
rect 356562 390766 359799 390768
rect 516558 390826 516618 391358
rect 519169 390826 519235 390829
rect 516558 390824 519235 390826
rect 516558 390768 519174 390824
rect 519230 390768 519235 390824
rect 516558 390766 519235 390768
rect 199193 390763 199259 390766
rect 359733 390763 359799 390766
rect 519169 390763 519235 390766
rect 196558 389194 196618 389862
rect 356562 389330 356622 389862
rect 359181 389330 359247 389333
rect 356562 389328 359247 389330
rect 356562 389272 359186 389328
rect 359242 389272 359247 389328
rect 356562 389270 359247 389272
rect 516558 389330 516618 389862
rect 519077 389330 519143 389333
rect 516558 389328 519143 389330
rect 516558 389272 519082 389328
rect 519138 389272 519143 389328
rect 516558 389270 519143 389272
rect 359181 389267 359247 389270
rect 519077 389267 519143 389270
rect 196558 389134 199578 389194
rect 199518 389061 199578 389134
rect 199469 389056 199578 389061
rect 199469 389000 199474 389056
rect 199530 389000 199578 389056
rect 199469 388998 199578 389000
rect 199469 388995 199535 388998
rect 196558 388514 196618 388638
rect 199837 388514 199903 388517
rect 196558 388512 199903 388514
rect 196558 388456 199842 388512
rect 199898 388456 199903 388512
rect 196558 388454 199903 388456
rect 199837 388451 199903 388454
rect 356562 388106 356622 388638
rect 359825 388106 359891 388109
rect 356562 388104 359891 388106
rect 356562 388048 359830 388104
rect 359886 388048 359891 388104
rect 356562 388046 359891 388048
rect 516558 388106 516618 388638
rect 519261 388106 519327 388109
rect 516558 388104 519327 388106
rect 516558 388048 519266 388104
rect 519322 388048 519327 388104
rect 516558 388046 519327 388048
rect 359825 388043 359891 388046
rect 519261 388043 519327 388046
rect 56593 384978 56659 384981
rect 216949 384978 217015 384981
rect 219390 384978 220064 384996
rect 56593 384976 60062 384978
rect 56593 384920 56598 384976
rect 56654 384920 60062 384976
rect 56593 384918 60062 384920
rect 216949 384976 220064 384978
rect 216949 384920 216954 384976
rect 217010 384936 220064 384976
rect 376937 384978 377003 384981
rect 379470 384978 380052 384996
rect 376937 384976 380052 384978
rect 217010 384920 219450 384936
rect 216949 384918 219450 384920
rect 376937 384920 376942 384976
rect 376998 384936 380052 384976
rect 376998 384920 379530 384936
rect 376937 384918 379530 384920
rect 56593 384915 56659 384918
rect 216949 384915 217015 384918
rect 376937 384915 377003 384918
rect -960 384284 480 384524
rect 51441 383618 51507 383621
rect 51574 383618 51580 383620
rect 51441 383616 51580 383618
rect 51441 383560 51446 383616
rect 51502 383560 51580 383616
rect 51441 383558 51580 383560
rect 51441 383555 51507 383558
rect 51574 383556 51580 383558
rect 51644 383556 51650 383620
rect 57462 383556 57468 383620
rect 57532 383618 57538 383620
rect 58433 383618 58499 383621
rect 57532 383616 58499 383618
rect 57532 383560 58438 383616
rect 58494 383560 58499 383616
rect 57532 383558 58499 383560
rect 57532 383556 57538 383558
rect 58433 383555 58499 383558
rect 57237 383346 57303 383349
rect 59494 383346 60032 383364
rect 57237 383344 60032 383346
rect 57237 383288 57242 383344
rect 57298 383304 60032 383344
rect 216673 383346 216739 383349
rect 219390 383346 220064 383364
rect 216673 383344 220064 383346
rect 57298 383288 59554 383304
rect 57237 383286 59554 383288
rect 216673 383288 216678 383344
rect 216734 383304 220064 383344
rect 376661 383346 376727 383349
rect 379470 383346 380052 383364
rect 376661 383344 380052 383346
rect 216734 383288 219450 383304
rect 216673 383286 219450 383288
rect 376661 383288 376666 383344
rect 376722 383304 380052 383344
rect 376722 383288 379530 383304
rect 376661 383286 379530 383288
rect 57237 383283 57303 383286
rect 216673 383283 216739 383286
rect 376661 383283 376727 383286
rect 56593 383074 56659 383077
rect 217041 383074 217107 383077
rect 219390 383074 220064 383092
rect 56593 383072 60062 383074
rect 56593 383016 56598 383072
rect 56654 383016 60062 383072
rect 56593 383014 60062 383016
rect 217041 383072 220064 383074
rect 217041 383016 217046 383072
rect 217102 383032 220064 383072
rect 376937 383074 377003 383077
rect 379470 383074 380052 383092
rect 376937 383072 380052 383074
rect 217102 383016 219450 383032
rect 217041 383014 219450 383016
rect 376937 383016 376942 383072
rect 376998 383032 380052 383072
rect 376998 383016 379530 383032
rect 376937 383014 379530 383016
rect 56593 383011 56659 383014
rect 217041 383011 217107 383014
rect 376937 383011 377003 383014
rect 207054 382332 207060 382396
rect 207124 382394 207130 382396
rect 208301 382394 208367 382397
rect 207124 382392 208367 382394
rect 207124 382336 208306 382392
rect 208362 382336 208367 382392
rect 207124 382334 208367 382336
rect 207124 382332 207130 382334
rect 208301 382331 208367 382334
rect 580441 378450 580507 378453
rect 583520 378450 584960 378540
rect 580441 378448 584960 378450
rect 580441 378392 580446 378448
rect 580502 378392 584960 378448
rect 580441 378390 584960 378392
rect 580441 378387 580507 378390
rect 583520 378300 584960 378390
rect 52821 375322 52887 375325
rect 53230 375322 53236 375324
rect 52821 375320 53236 375322
rect 52821 375264 52826 375320
rect 52882 375264 53236 375320
rect 52821 375262 53236 375264
rect 52821 375259 52887 375262
rect 53230 375260 53236 375262
rect 53300 375260 53306 375324
rect 198222 375260 198228 375324
rect 198292 375322 198298 375324
rect 198641 375322 198707 375325
rect 198292 375320 198707 375322
rect 198292 375264 198646 375320
rect 198702 375264 198707 375320
rect 198292 375262 198707 375264
rect 198292 375260 198298 375262
rect 198641 375259 198707 375262
rect 200982 375260 200988 375324
rect 201052 375322 201058 375324
rect 201401 375322 201467 375325
rect 201052 375320 201467 375322
rect 201052 375264 201406 375320
rect 201462 375264 201467 375320
rect 201052 375262 201467 375264
rect 201052 375260 201058 375262
rect 201401 375259 201467 375262
rect 204294 375260 204300 375324
rect 204364 375322 204370 375324
rect 205541 375322 205607 375325
rect 204364 375320 205607 375322
rect 204364 375264 205546 375320
rect 205602 375264 205607 375320
rect 204364 375262 205607 375264
rect 204364 375260 204370 375262
rect 205541 375259 205607 375262
rect 216857 375322 216923 375325
rect 217133 375322 217199 375325
rect 216857 375320 217199 375322
rect 216857 375264 216862 375320
rect 216918 375264 217138 375320
rect 217194 375264 217199 375320
rect 216857 375262 217199 375264
rect 216857 375259 216923 375262
rect 217133 375259 217199 375262
rect 46013 375050 46079 375053
rect 216765 375050 216831 375053
rect 405917 375052 405983 375053
rect 407757 375052 407823 375053
rect 425053 375052 425119 375053
rect 440325 375052 440391 375053
rect 443085 375052 443151 375053
rect 452837 375052 452903 375053
rect 405917 375050 405964 375052
rect 46013 375048 216831 375050
rect 46013 374992 46018 375048
rect 46074 374992 216770 375048
rect 216826 374992 216831 375048
rect 46013 374990 216831 374992
rect 405872 375048 405964 375050
rect 405872 374992 405922 375048
rect 405872 374990 405964 374992
rect 46013 374987 46079 374990
rect 216765 374987 216831 374990
rect 405917 374988 405964 374990
rect 406028 374988 406034 375052
rect 407757 375050 407804 375052
rect 407712 375048 407804 375050
rect 407712 374992 407762 375048
rect 407712 374990 407804 374992
rect 407757 374988 407804 374990
rect 407868 374988 407874 375052
rect 425053 375050 425100 375052
rect 425008 375048 425100 375050
rect 425008 374992 425058 375048
rect 425008 374990 425100 374992
rect 425053 374988 425100 374990
rect 425164 374988 425170 375052
rect 440325 375050 440372 375052
rect 440280 375048 440372 375050
rect 440280 374992 440330 375048
rect 440280 374990 440372 374992
rect 440325 374988 440372 374990
rect 440436 374988 440442 375052
rect 443085 375050 443132 375052
rect 443040 375048 443132 375050
rect 443040 374992 443090 375048
rect 443040 374990 443132 374992
rect 443085 374988 443132 374990
rect 443196 374988 443202 375052
rect 452837 375050 452884 375052
rect 452792 375048 452884 375050
rect 452792 374992 452842 375048
rect 452792 374990 452884 374992
rect 452837 374988 452884 374990
rect 452948 374988 452954 375052
rect 405917 374987 405983 374988
rect 407757 374987 407823 374988
rect 425053 374987 425119 374988
rect 440325 374987 440391 374988
rect 443085 374987 443151 374988
rect 452837 374987 452903 374988
rect 52361 374914 52427 374917
rect 216857 374914 216923 374917
rect 52361 374912 216923 374914
rect 52361 374856 52366 374912
rect 52422 374856 216862 374912
rect 216918 374856 216923 374912
rect 52361 374854 216923 374856
rect 52361 374851 52427 374854
rect 216857 374851 216923 374854
rect 163405 374644 163471 374645
rect 165981 374644 166047 374645
rect 163360 374580 163366 374644
rect 163430 374642 163471 374644
rect 163430 374640 163522 374642
rect 163466 374584 163522 374640
rect 163430 374582 163522 374584
rect 163430 374580 163471 374582
rect 165944 374580 165950 374644
rect 166014 374642 166047 374644
rect 166014 374640 166106 374642
rect 166042 374584 166106 374640
rect 166014 374582 166106 374584
rect 166014 374580 166047 374582
rect 206502 374580 206508 374644
rect 206572 374642 206578 374644
rect 206829 374642 206895 374645
rect 206572 374640 206895 374642
rect 206572 374584 206834 374640
rect 206890 374584 206895 374640
rect 206572 374582 206895 374584
rect 206572 374580 206578 374582
rect 163405 374579 163471 374580
rect 165981 374579 166047 374580
rect 206829 374579 206895 374582
rect 208342 374580 208348 374644
rect 208412 374642 208418 374644
rect 209681 374642 209747 374645
rect 208412 374640 209747 374642
rect 208412 374584 209686 374640
rect 209742 374584 209747 374640
rect 208412 374582 209747 374584
rect 208412 374580 208418 374582
rect 209681 374579 209747 374582
rect 209814 374580 209820 374644
rect 209884 374642 209890 374644
rect 211061 374642 211127 374645
rect 410701 374644 410767 374645
rect 410701 374642 410742 374644
rect 209884 374640 211127 374642
rect 209884 374584 211066 374640
rect 211122 374584 211127 374640
rect 209884 374582 211127 374584
rect 410650 374640 410742 374642
rect 410650 374584 410706 374640
rect 410650 374582 410742 374584
rect 209884 374580 209890 374582
rect 211061 374579 211127 374582
rect 410701 374580 410742 374582
rect 410806 374580 410812 374644
rect 410701 374579 410767 374580
rect 93577 374508 93643 374509
rect 103513 374508 103579 374509
rect 116025 374508 116091 374509
rect 143533 374508 143599 374509
rect 146201 374508 146267 374509
rect 153469 374508 153535 374509
rect 156505 374508 156571 374509
rect 158529 374508 158595 374509
rect 160921 374508 160987 374509
rect 235993 374508 236059 374509
rect 244273 374508 244339 374509
rect 250069 374508 250135 374509
rect 93577 374506 93598 374508
rect 93506 374504 93598 374506
rect 93506 374448 93582 374504
rect 93506 374446 93598 374448
rect 93577 374444 93598 374446
rect 93662 374444 93668 374508
rect 103513 374504 103526 374508
rect 103590 374506 103596 374508
rect 116025 374506 116038 374508
rect 103513 374448 103518 374504
rect 103513 374444 103526 374448
rect 103590 374446 103670 374506
rect 115946 374504 116038 374506
rect 115946 374448 116030 374504
rect 115946 374446 116038 374448
rect 103590 374444 103596 374446
rect 116025 374444 116038 374446
rect 116102 374444 116108 374508
rect 143504 374444 143510 374508
rect 143574 374506 143599 374508
rect 143574 374504 143666 374506
rect 143594 374448 143666 374504
rect 143574 374446 143666 374448
rect 143574 374444 143599 374446
rect 146150 374444 146156 374508
rect 146220 374506 146267 374508
rect 146220 374504 146312 374506
rect 146262 374448 146312 374504
rect 146220 374446 146312 374448
rect 146220 374444 146267 374446
rect 153432 374444 153438 374508
rect 153502 374506 153535 374508
rect 153502 374504 153594 374506
rect 153530 374448 153594 374504
rect 153502 374446 153594 374448
rect 153502 374444 153535 374446
rect 156454 374444 156460 374508
rect 156524 374506 156571 374508
rect 156524 374504 156616 374506
rect 156566 374448 156616 374504
rect 156524 374446 156616 374448
rect 156524 374444 156571 374446
rect 158478 374444 158484 374508
rect 158548 374506 158595 374508
rect 158548 374504 158640 374506
rect 158590 374448 158640 374504
rect 158548 374446 158640 374448
rect 158548 374444 158595 374446
rect 160912 374444 160918 374508
rect 160982 374506 160988 374508
rect 235993 374506 236054 374508
rect 160982 374446 161074 374506
rect 235962 374504 236054 374506
rect 235962 374448 235998 374504
rect 235962 374446 236054 374448
rect 160982 374444 160988 374446
rect 235993 374444 236054 374446
rect 236118 374444 236124 374508
rect 244222 374444 244228 374508
rect 244292 374506 244339 374508
rect 244292 374504 244384 374506
rect 244334 374448 244384 374504
rect 244292 374446 244384 374448
rect 244292 374444 244339 374446
rect 250056 374444 250062 374508
rect 250126 374506 250135 374508
rect 250713 374508 250779 374509
rect 251265 374508 251331 374509
rect 256049 374508 256115 374509
rect 250713 374506 250742 374508
rect 250126 374504 250218 374506
rect 250130 374448 250218 374504
rect 250126 374446 250218 374448
rect 250650 374504 250742 374506
rect 250650 374448 250718 374504
rect 250650 374446 250742 374448
rect 250126 374444 250135 374446
rect 93577 374443 93643 374444
rect 103513 374443 103579 374444
rect 116025 374443 116091 374444
rect 143533 374443 143599 374444
rect 146201 374443 146267 374444
rect 153469 374443 153535 374444
rect 156505 374443 156571 374444
rect 158529 374443 158595 374444
rect 160921 374443 160987 374444
rect 235993 374443 236059 374444
rect 244273 374443 244339 374444
rect 250069 374443 250135 374444
rect 250713 374444 250742 374446
rect 250806 374444 250812 374508
rect 251265 374506 251286 374508
rect 251194 374504 251286 374506
rect 251194 374448 251270 374504
rect 251194 374446 251286 374448
rect 251265 374444 251286 374446
rect 251350 374444 251356 374508
rect 256040 374444 256046 374508
rect 256110 374506 256116 374508
rect 270493 374506 270559 374509
rect 320909 374508 320975 374509
rect 433609 374508 433675 374509
rect 271136 374506 271142 374508
rect 256110 374446 256202 374506
rect 270493 374504 271142 374506
rect 270493 374448 270498 374504
rect 270554 374448 271142 374504
rect 270493 374446 271142 374448
rect 256110 374444 256116 374446
rect 250713 374443 250779 374444
rect 251265 374443 251331 374444
rect 256049 374443 256115 374444
rect 270493 374443 270559 374446
rect 271136 374444 271142 374446
rect 271206 374444 271212 374508
rect 320909 374506 320918 374508
rect 320826 374504 320918 374506
rect 320826 374448 320914 374504
rect 320826 374446 320918 374448
rect 320909 374444 320918 374446
rect 320982 374444 320988 374508
rect 433584 374444 433590 374508
rect 433654 374506 433675 374508
rect 436001 374508 436067 374509
rect 438485 374508 438551 374509
rect 436001 374506 436038 374508
rect 433654 374504 433746 374506
rect 433670 374448 433746 374504
rect 433654 374446 433746 374448
rect 435946 374504 436038 374506
rect 435946 374448 436006 374504
rect 435946 374446 436038 374448
rect 433654 374444 433675 374446
rect 320909 374443 320975 374444
rect 433609 374443 433675 374444
rect 436001 374444 436038 374446
rect 436102 374444 436108 374508
rect 438480 374506 438486 374508
rect 438394 374446 438486 374506
rect 438480 374444 438486 374446
rect 438550 374444 438556 374508
rect 436001 374443 436067 374444
rect 438485 374443 438551 374444
rect 215845 374370 215911 374373
rect 263726 374370 263732 374372
rect 215845 374368 263732 374370
rect 215845 374312 215850 374368
rect 215906 374312 263732 374368
rect 215845 374310 263732 374312
rect 215845 374307 215911 374310
rect 263726 374308 263732 374310
rect 263796 374308 263802 374372
rect 148961 374236 149027 374237
rect 148910 374172 148916 374236
rect 148980 374234 149027 374236
rect 218237 374234 218303 374237
rect 222009 374234 222075 374237
rect 148980 374232 149072 374234
rect 149022 374176 149072 374232
rect 148980 374174 149072 374176
rect 218237 374232 222075 374234
rect 218237 374176 218242 374232
rect 218298 374176 222014 374232
rect 222070 374176 222075 374232
rect 218237 374174 222075 374176
rect 148980 374172 149027 374174
rect 148961 374171 149027 374172
rect 218237 374171 218303 374174
rect 222009 374171 222075 374174
rect 219617 374098 219683 374101
rect 221917 374098 221983 374101
rect 219617 374096 221983 374098
rect 219617 374040 219622 374096
rect 219678 374040 221922 374096
rect 221978 374040 221983 374096
rect 219617 374038 221983 374040
rect 219617 374035 219683 374038
rect 221917 374035 221983 374038
rect 270217 374098 270283 374101
rect 416037 374100 416103 374101
rect 275134 374098 275140 374100
rect 270217 374096 275140 374098
rect 270217 374040 270222 374096
rect 270278 374040 275140 374096
rect 270217 374038 275140 374040
rect 270217 374035 270283 374038
rect 275134 374036 275140 374038
rect 275204 374036 275210 374100
rect 416037 374098 416084 374100
rect 415992 374096 416084 374098
rect 415992 374040 416042 374096
rect 415992 374038 416084 374040
rect 416037 374036 416084 374038
rect 416148 374036 416154 374100
rect 416037 374035 416103 374036
rect 40861 373962 40927 373965
rect 199469 373962 199535 373965
rect 40861 373960 199535 373962
rect 40861 373904 40866 373960
rect 40922 373904 199474 373960
rect 199530 373904 199535 373960
rect 40861 373902 199535 373904
rect 40861 373899 40927 373902
rect 199469 373899 199535 373902
rect 377438 373900 377444 373964
rect 377508 373962 377514 373964
rect 485814 373962 485820 373964
rect 377508 373902 485820 373962
rect 377508 373900 377514 373902
rect 485814 373900 485820 373902
rect 485884 373900 485890 373964
rect 83774 373764 83780 373828
rect 83844 373826 83850 373828
rect 207197 373826 207263 373829
rect 83844 373824 207263 373826
rect 83844 373768 207202 373824
rect 207258 373768 207263 373824
rect 83844 373766 207263 373768
rect 83844 373764 83850 373766
rect 207197 373763 207263 373766
rect 262765 373826 262831 373829
rect 268510 373826 268516 373828
rect 262765 373824 268516 373826
rect 262765 373768 262770 373824
rect 262826 373768 268516 373824
rect 262765 373766 268516 373768
rect 262765 373763 262831 373766
rect 268510 373764 268516 373766
rect 268580 373764 268586 373828
rect 377622 373764 377628 373828
rect 377692 373826 377698 373828
rect 460974 373826 460980 373828
rect 377692 373766 460980 373826
rect 377692 373764 377698 373766
rect 460974 373764 460980 373766
rect 461044 373764 461050 373828
rect 100845 373692 100911 373693
rect 107837 373692 107903 373693
rect 113541 373692 113607 373693
rect 118325 373692 118391 373693
rect 121361 373692 121427 373693
rect 125777 373692 125843 373693
rect 128905 373692 128971 373693
rect 100845 373690 100892 373692
rect 100800 373688 100892 373690
rect 100800 373632 100850 373688
rect 100800 373630 100892 373632
rect 100845 373628 100892 373630
rect 100956 373628 100962 373692
rect 107837 373690 107884 373692
rect 107792 373688 107884 373690
rect 107792 373632 107842 373688
rect 107792 373630 107884 373632
rect 107837 373628 107884 373630
rect 107948 373628 107954 373692
rect 113541 373690 113588 373692
rect 113496 373688 113588 373690
rect 113496 373632 113546 373688
rect 113496 373630 113588 373632
rect 113541 373628 113588 373630
rect 113652 373628 113658 373692
rect 118325 373690 118372 373692
rect 118280 373688 118372 373690
rect 118280 373632 118330 373688
rect 118280 373630 118372 373632
rect 118325 373628 118372 373630
rect 118436 373628 118442 373692
rect 121310 373690 121316 373692
rect 121270 373630 121316 373690
rect 121380 373688 121427 373692
rect 125726 373690 125732 373692
rect 121422 373632 121427 373688
rect 121310 373628 121316 373630
rect 121380 373628 121427 373632
rect 125686 373630 125732 373690
rect 125796 373688 125843 373692
rect 128854 373690 128860 373692
rect 125838 373632 125843 373688
rect 125726 373628 125732 373630
rect 125796 373628 125843 373632
rect 128814 373630 128860 373690
rect 128924 373688 128971 373692
rect 128966 373632 128971 373688
rect 128854 373628 128860 373630
rect 128924 373628 128971 373632
rect 100845 373627 100911 373628
rect 107837 373627 107903 373628
rect 113541 373627 113607 373628
rect 118325 373627 118391 373628
rect 121361 373627 121427 373628
rect 125777 373627 125843 373628
rect 128905 373627 128971 373628
rect 131021 373692 131087 373693
rect 133689 373692 133755 373693
rect 136449 373692 136515 373693
rect 139209 373692 139275 373693
rect 141601 373692 141667 373693
rect 151721 373692 151787 373693
rect 131021 373688 131068 373692
rect 131132 373690 131138 373692
rect 133638 373690 133644 373692
rect 131021 373632 131026 373688
rect 131021 373628 131068 373632
rect 131132 373630 131178 373690
rect 133598 373630 133644 373690
rect 133708 373688 133755 373692
rect 136398 373690 136404 373692
rect 133750 373632 133755 373688
rect 131132 373628 131138 373630
rect 133638 373628 133644 373630
rect 133708 373628 133755 373632
rect 136358 373630 136404 373690
rect 136468 373688 136515 373692
rect 139158 373690 139164 373692
rect 136510 373632 136515 373688
rect 136398 373628 136404 373630
rect 136468 373628 136515 373632
rect 139118 373630 139164 373690
rect 139228 373688 139275 373692
rect 141550 373690 141556 373692
rect 139270 373632 139275 373688
rect 139158 373628 139164 373630
rect 139228 373628 139275 373632
rect 141510 373630 141556 373690
rect 141620 373688 141667 373692
rect 151670 373690 151676 373692
rect 141662 373632 141667 373688
rect 141550 373628 141556 373630
rect 141620 373628 141667 373632
rect 151630 373630 151676 373690
rect 151740 373688 151787 373692
rect 151782 373632 151787 373688
rect 151670 373628 151676 373630
rect 151740 373628 151787 373632
rect 131021 373627 131087 373628
rect 133689 373627 133755 373628
rect 136449 373627 136515 373628
rect 139209 373627 139275 373628
rect 141601 373627 141667 373628
rect 151721 373627 151787 373628
rect 211153 373690 211219 373693
rect 211429 373690 211495 373693
rect 221825 373690 221891 373693
rect 418245 373692 418311 373693
rect 423029 373692 423095 373693
rect 426893 373692 426959 373693
rect 445845 373692 445911 373693
rect 211153 373688 221891 373690
rect 211153 373632 211158 373688
rect 211214 373632 211434 373688
rect 211490 373632 221830 373688
rect 221886 373632 221891 373688
rect 211153 373630 221891 373632
rect 211153 373627 211219 373630
rect 211429 373627 211495 373630
rect 221825 373627 221891 373630
rect 359590 373628 359596 373692
rect 359660 373690 359666 373692
rect 418245 373690 418292 373692
rect 359660 373630 412650 373690
rect 418200 373688 418292 373690
rect 418200 373632 418250 373688
rect 418200 373630 418292 373632
rect 359660 373628 359666 373630
rect 105445 373556 105511 373557
rect 110413 373556 110479 373557
rect 105445 373554 105492 373556
rect 105400 373552 105492 373554
rect 105400 373496 105450 373552
rect 105400 373494 105492 373496
rect 105445 373492 105492 373494
rect 105556 373492 105562 373556
rect 110413 373554 110460 373556
rect 110368 373552 110460 373554
rect 110368 373496 110418 373552
rect 110368 373494 110460 373496
rect 110413 373492 110460 373494
rect 110524 373492 110530 373556
rect 119838 373492 119844 373556
rect 119908 373554 119914 373556
rect 209589 373554 209655 373557
rect 255405 373556 255471 373557
rect 256693 373556 256759 373557
rect 255405 373554 255452 373556
rect 119908 373552 219450 373554
rect 119908 373496 209594 373552
rect 209650 373496 219450 373552
rect 119908 373494 219450 373496
rect 255360 373552 255452 373554
rect 255360 373496 255410 373552
rect 255360 373494 255452 373496
rect 119908 373492 119914 373494
rect 105445 373491 105511 373492
rect 110413 373491 110479 373492
rect 209589 373491 209655 373494
rect 88333 373420 88399 373421
rect 96061 373420 96127 373421
rect 98269 373420 98335 373421
rect 122925 373420 122991 373421
rect 88333 373418 88380 373420
rect 88288 373416 88380 373418
rect 88288 373360 88338 373416
rect 88288 373358 88380 373360
rect 88333 373356 88380 373358
rect 88444 373356 88450 373420
rect 96061 373418 96108 373420
rect 96016 373416 96108 373418
rect 96016 373360 96066 373416
rect 96016 373358 96108 373360
rect 96061 373356 96108 373358
rect 96172 373356 96178 373420
rect 98269 373418 98316 373420
rect 98224 373416 98316 373418
rect 98224 373360 98274 373416
rect 98224 373358 98316 373360
rect 98269 373356 98316 373358
rect 98380 373356 98386 373420
rect 122925 373418 122972 373420
rect 122880 373416 122972 373418
rect 122880 373360 122930 373416
rect 122880 373358 122972 373360
rect 122925 373356 122972 373358
rect 123036 373356 123042 373420
rect 197261 373418 197327 373421
rect 210049 373418 210115 373421
rect 197261 373416 210115 373418
rect 197261 373360 197266 373416
rect 197322 373360 210054 373416
rect 210110 373360 210115 373416
rect 197261 373358 210115 373360
rect 88333 373355 88399 373356
rect 96061 373355 96127 373356
rect 98269 373355 98335 373356
rect 122925 373355 122991 373356
rect 197261 373355 197327 373358
rect 210049 373355 210115 373358
rect 40585 373282 40651 373285
rect 200021 373282 200087 373285
rect 203241 373282 203307 373285
rect 40585 373280 203307 373282
rect 40585 373224 40590 373280
rect 40646 373224 200026 373280
rect 200082 373224 203246 373280
rect 203302 373224 203307 373280
rect 40585 373222 203307 373224
rect 219390 373282 219450 373494
rect 255405 373492 255452 373494
rect 255516 373492 255522 373556
rect 256693 373554 256740 373556
rect 256648 373552 256740 373554
rect 256648 373496 256698 373552
rect 256648 373494 256740 373496
rect 256693 373492 256740 373494
rect 256804 373492 256810 373556
rect 412590 373554 412650 373630
rect 418245 373628 418292 373630
rect 418356 373628 418362 373692
rect 423029 373690 423076 373692
rect 422984 373688 423076 373690
rect 422984 373632 423034 373688
rect 422984 373630 423076 373632
rect 423029 373628 423076 373630
rect 423140 373628 423146 373692
rect 426893 373690 426940 373692
rect 426848 373688 426940 373690
rect 426848 373632 426898 373688
rect 426848 373630 426940 373632
rect 426893 373628 426940 373630
rect 427004 373628 427010 373692
rect 445845 373690 445892 373692
rect 445800 373688 445892 373690
rect 445800 373632 445850 373688
rect 445800 373630 445892 373632
rect 445845 373628 445892 373630
rect 445956 373628 445962 373692
rect 418245 373627 418311 373628
rect 423029 373627 423095 373628
rect 426893 373627 426959 373628
rect 445845 373627 445911 373628
rect 450261 373556 450327 373557
rect 455413 373556 455479 373557
rect 427854 373554 427860 373556
rect 412590 373494 427860 373554
rect 427854 373492 427860 373494
rect 427924 373492 427930 373556
rect 450261 373554 450308 373556
rect 450216 373552 450308 373554
rect 450216 373496 450266 373552
rect 450216 373494 450308 373496
rect 450261 373492 450308 373494
rect 450372 373492 450378 373556
rect 455413 373554 455460 373556
rect 455368 373552 455460 373554
rect 455368 373496 455418 373552
rect 455368 373494 455460 373496
rect 455413 373492 455460 373494
rect 455524 373492 455530 373556
rect 255405 373491 255471 373492
rect 256693 373491 256759 373492
rect 450261 373491 450327 373492
rect 455413 373491 455479 373492
rect 236453 373420 236519 373421
rect 242893 373420 242959 373421
rect 260005 373420 260071 373421
rect 269205 373420 269271 373421
rect 447685 373420 447751 373421
rect 462773 373420 462839 373421
rect 236453 373418 236500 373420
rect 236408 373416 236500 373418
rect 236408 373360 236458 373416
rect 236408 373358 236500 373360
rect 236453 373356 236500 373358
rect 236564 373356 236570 373420
rect 242893 373418 242940 373420
rect 242848 373416 242940 373418
rect 242848 373360 242898 373416
rect 242848 373358 242940 373360
rect 242893 373356 242940 373358
rect 243004 373356 243010 373420
rect 260005 373418 260052 373420
rect 259960 373416 260052 373418
rect 259960 373360 260010 373416
rect 259960 373358 260052 373360
rect 260005 373356 260052 373358
rect 260116 373356 260122 373420
rect 269205 373418 269252 373420
rect 269160 373416 269252 373418
rect 269160 373360 269210 373416
rect 269160 373358 269252 373360
rect 269205 373356 269252 373358
rect 269316 373356 269322 373420
rect 447685 373418 447732 373420
rect 447640 373416 447732 373418
rect 447640 373360 447690 373416
rect 447640 373358 447732 373360
rect 447685 373356 447732 373358
rect 447796 373356 447802 373420
rect 462773 373418 462820 373420
rect 462728 373416 462820 373418
rect 462728 373360 462778 373416
rect 462728 373358 462820 373360
rect 462773 373356 462820 373358
rect 462884 373356 462890 373420
rect 236453 373355 236519 373356
rect 242893 373355 242959 373356
rect 260005 373355 260071 373356
rect 269205 373355 269271 373356
rect 447685 373355 447751 373356
rect 462773 373355 462839 373356
rect 220813 373282 220879 373285
rect 278814 373282 278820 373284
rect 219390 373280 278820 373282
rect 219390 373224 220818 373280
rect 220874 373224 278820 373280
rect 219390 373222 278820 373224
rect 40585 373219 40651 373222
rect 200021 373219 200087 373222
rect 203241 373219 203307 373222
rect 220813 373219 220879 373222
rect 278814 373220 278820 373222
rect 278884 373220 278890 373284
rect 359958 373220 359964 373284
rect 360028 373282 360034 373284
rect 376661 373282 376727 373285
rect 408534 373282 408540 373284
rect 360028 373280 408540 373282
rect 360028 373224 376666 373280
rect 376722 373224 408540 373280
rect 360028 373222 408540 373224
rect 360028 373220 360034 373222
rect 376661 373219 376727 373222
rect 408534 373220 408540 373222
rect 408604 373220 408610 373284
rect 90173 373148 90239 373149
rect 92381 373148 92447 373149
rect 90173 373146 90220 373148
rect 90128 373144 90220 373146
rect 90128 373088 90178 373144
rect 90128 373086 90220 373088
rect 90173 373084 90220 373086
rect 90284 373084 90290 373148
rect 92381 373144 92428 373148
rect 92492 373146 92498 373148
rect 92381 373088 92386 373144
rect 92381 373084 92428 373088
rect 92492 373086 92538 373146
rect 92492 373084 92498 373086
rect 95182 373084 95188 373148
rect 95252 373146 95258 373148
rect 212717 373146 212783 373149
rect 219893 373146 219959 373149
rect 220721 373146 220787 373149
rect 247125 373148 247191 373149
rect 253933 373148 253999 373149
rect 247125 373146 247172 373148
rect 95252 373144 220787 373146
rect 95252 373088 212722 373144
rect 212778 373088 219898 373144
rect 219954 373088 220726 373144
rect 220782 373088 220787 373144
rect 95252 373086 220787 373088
rect 247080 373144 247172 373146
rect 247080 373088 247130 373144
rect 247080 373086 247172 373088
rect 95252 373084 95258 373086
rect 90173 373083 90239 373084
rect 92381 373083 92447 373084
rect 212717 373083 212783 373086
rect 219893 373083 219959 373086
rect 220721 373083 220787 373086
rect 247125 373084 247172 373086
rect 247236 373084 247242 373148
rect 253933 373146 253980 373148
rect 253888 373144 253980 373146
rect 253888 373088 253938 373144
rect 253888 373086 253980 373088
rect 253933 373084 253980 373086
rect 254044 373084 254050 373148
rect 257838 373084 257844 373148
rect 257908 373146 257914 373148
rect 258073 373146 258139 373149
rect 261293 373148 261359 373149
rect 264973 373148 265039 373149
rect 300853 373148 300919 373149
rect 261293 373146 261340 373148
rect 257908 373144 258139 373146
rect 257908 373088 258078 373144
rect 258134 373088 258139 373144
rect 257908 373086 258139 373088
rect 261248 373144 261340 373146
rect 261248 373088 261298 373144
rect 261248 373086 261340 373088
rect 257908 373084 257914 373086
rect 247125 373083 247191 373084
rect 253933 373083 253999 373084
rect 258073 373083 258139 373086
rect 261293 373084 261340 373086
rect 261404 373084 261410 373148
rect 264973 373146 265020 373148
rect 264928 373144 265020 373146
rect 264928 373088 264978 373144
rect 264928 373086 265020 373088
rect 264973 373084 265020 373086
rect 265084 373084 265090 373148
rect 300853 373146 300900 373148
rect 300808 373144 300900 373146
rect 300808 373088 300858 373144
rect 300808 373086 300900 373088
rect 300853 373084 300900 373086
rect 300964 373084 300970 373148
rect 261293 373083 261359 373084
rect 264973 373083 265039 373084
rect 300853 373083 300919 373084
rect 58525 372874 58591 372877
rect 60733 372874 60799 372877
rect 58525 372872 60799 372874
rect 58525 372816 58530 372872
rect 58586 372816 60738 372872
rect 60794 372816 60799 372872
rect 58525 372814 60799 372816
rect 58525 372811 58591 372814
rect 60733 372811 60799 372814
rect 57278 372676 57284 372740
rect 57348 372738 57354 372740
rect 58617 372738 58683 372741
rect 57348 372736 58683 372738
rect 57348 372680 58622 372736
rect 58678 372680 58683 372736
rect 57348 372678 58683 372680
rect 57348 372676 57354 372678
rect 58617 372675 58683 372678
rect 216990 372676 216996 372740
rect 217060 372738 217066 372740
rect 219249 372738 219315 372741
rect 217060 372736 219315 372738
rect 217060 372680 219254 372736
rect 219310 372680 219315 372736
rect 217060 372678 219315 372680
rect 217060 372676 217066 372678
rect 219249 372675 219315 372678
rect 252553 372738 252619 372741
rect 252870 372738 252876 372740
rect 252553 372736 252876 372738
rect 252553 372680 252558 372736
rect 252614 372680 252876 372736
rect 252553 372678 252876 372680
rect 252553 372675 252619 372678
rect 252870 372676 252876 372678
rect 252940 372676 252946 372740
rect 362902 372676 362908 372740
rect 362972 372738 362978 372740
rect 364241 372738 364307 372741
rect 362972 372736 364307 372738
rect 362972 372680 364246 372736
rect 364302 372680 364307 372736
rect 362972 372678 364307 372680
rect 362972 372676 362978 372678
rect 364241 372675 364307 372678
rect 371141 372738 371207 372741
rect 376886 372738 376892 372740
rect 371141 372736 376892 372738
rect 371141 372680 371146 372736
rect 371202 372680 376892 372736
rect 371141 372678 376892 372680
rect 371141 372675 371207 372678
rect 376886 372676 376892 372678
rect 376956 372676 376962 372740
rect 77201 372604 77267 372605
rect 81985 372604 82051 372605
rect 84745 372604 84811 372605
rect 86769 372604 86835 372605
rect 88057 372604 88123 372605
rect 89345 372604 89411 372605
rect 77150 372602 77156 372604
rect 77110 372542 77156 372602
rect 77220 372600 77267 372604
rect 81934 372602 81940 372604
rect 77262 372544 77267 372600
rect 77150 372540 77156 372542
rect 77220 372540 77267 372544
rect 81894 372542 81940 372602
rect 82004 372600 82051 372604
rect 84694 372602 84700 372604
rect 82046 372544 82051 372600
rect 81934 372540 81940 372542
rect 82004 372540 82051 372544
rect 84654 372542 84700 372602
rect 84764 372600 84811 372604
rect 86718 372602 86724 372604
rect 84806 372544 84811 372600
rect 84694 372540 84700 372542
rect 84764 372540 84811 372544
rect 86678 372542 86724 372602
rect 86788 372600 86835 372604
rect 88006 372602 88012 372604
rect 86830 372544 86835 372600
rect 86718 372540 86724 372542
rect 86788 372540 86835 372544
rect 87966 372542 88012 372602
rect 88076 372600 88123 372604
rect 89294 372602 89300 372604
rect 88118 372544 88123 372600
rect 88006 372540 88012 372542
rect 88076 372540 88123 372544
rect 89254 372542 89300 372602
rect 89364 372600 89411 372604
rect 89406 372544 89411 372600
rect 89294 372540 89300 372542
rect 89364 372540 89411 372544
rect 90030 372540 90036 372604
rect 90100 372602 90106 372604
rect 90725 372602 90791 372605
rect 90100 372600 90791 372602
rect 90100 372544 90730 372600
rect 90786 372544 90791 372600
rect 90100 372542 90791 372544
rect 90100 372540 90106 372542
rect 77201 372539 77267 372540
rect 81985 372539 82051 372540
rect 84745 372539 84811 372540
rect 86769 372539 86835 372540
rect 88057 372539 88123 372540
rect 89345 372539 89411 372540
rect 90725 372539 90791 372542
rect 91502 372540 91508 372604
rect 91572 372602 91578 372604
rect 92197 372602 92263 372605
rect 91572 372600 92263 372602
rect 91572 372544 92202 372600
rect 92258 372544 92263 372600
rect 91572 372542 92263 372544
rect 91572 372540 91578 372542
rect 92197 372539 92263 372542
rect 93342 372540 93348 372604
rect 93412 372602 93418 372604
rect 93577 372602 93643 372605
rect 102041 372604 102107 372605
rect 112897 372604 112963 372605
rect 101990 372602 101996 372604
rect 93412 372600 93643 372602
rect 93412 372544 93582 372600
rect 93638 372544 93643 372600
rect 93412 372542 93643 372544
rect 101950 372542 101996 372602
rect 102060 372600 102107 372604
rect 112846 372602 112852 372604
rect 102102 372544 102107 372600
rect 93412 372540 93418 372542
rect 93577 372539 93643 372542
rect 101990 372540 101996 372542
rect 102060 372540 102107 372544
rect 112806 372542 112852 372602
rect 112916 372600 112963 372604
rect 112958 372544 112963 372600
rect 112846 372540 112852 372542
rect 112916 372540 112963 372544
rect 102041 372539 102107 372540
rect 112897 372539 112963 372540
rect 114461 372604 114527 372605
rect 238109 372604 238175 372605
rect 239305 372604 239371 372605
rect 240409 372604 240475 372605
rect 241697 372604 241763 372605
rect 114461 372600 114508 372604
rect 114572 372602 114578 372604
rect 114461 372544 114466 372600
rect 114461 372540 114508 372544
rect 114572 372542 114618 372602
rect 238109 372600 238156 372604
rect 238220 372602 238226 372604
rect 239254 372602 239260 372604
rect 238109 372544 238114 372600
rect 114572 372540 114578 372542
rect 238109 372540 238156 372544
rect 238220 372542 238266 372602
rect 239214 372542 239260 372602
rect 239324 372600 239371 372604
rect 240358 372602 240364 372604
rect 239366 372544 239371 372600
rect 238220 372540 238226 372542
rect 239254 372540 239260 372542
rect 239324 372540 239371 372544
rect 240318 372542 240364 372602
rect 240428 372600 240475 372604
rect 241646 372602 241652 372604
rect 240470 372544 240475 372600
rect 240358 372540 240364 372542
rect 240428 372540 240475 372544
rect 241606 372542 241652 372602
rect 241716 372600 241763 372604
rect 241758 372544 241763 372600
rect 241646 372540 241652 372542
rect 241716 372540 241763 372544
rect 114461 372539 114527 372540
rect 238109 372539 238175 372540
rect 239305 372539 239371 372540
rect 240409 372539 240475 372540
rect 241697 372539 241763 372540
rect 244273 372602 244339 372605
rect 248413 372604 248479 372605
rect 244774 372602 244780 372604
rect 244273 372600 244780 372602
rect 244273 372544 244278 372600
rect 244334 372544 244780 372600
rect 244273 372542 244780 372544
rect 244273 372539 244339 372542
rect 244774 372540 244780 372542
rect 244844 372540 244850 372604
rect 248413 372600 248460 372604
rect 248524 372602 248530 372604
rect 251173 372602 251239 372605
rect 259453 372604 259519 372605
rect 262213 372604 262279 372605
rect 266353 372604 266419 372605
rect 251766 372602 251772 372604
rect 248413 372544 248418 372600
rect 248413 372540 248460 372544
rect 248524 372542 248570 372602
rect 251173 372600 251772 372602
rect 251173 372544 251178 372600
rect 251234 372544 251772 372600
rect 251173 372542 251772 372544
rect 248524 372540 248530 372542
rect 248413 372539 248479 372540
rect 251173 372539 251239 372542
rect 251766 372540 251772 372542
rect 251836 372540 251842 372604
rect 259453 372602 259500 372604
rect 259408 372600 259500 372602
rect 259408 372544 259458 372600
rect 259408 372542 259500 372544
rect 259453 372540 259500 372542
rect 259564 372540 259570 372604
rect 262213 372602 262260 372604
rect 262168 372600 262260 372602
rect 262168 372544 262218 372600
rect 262168 372542 262260 372544
rect 262213 372540 262260 372542
rect 262324 372540 262330 372604
rect 266302 372540 266308 372604
rect 266372 372602 266419 372604
rect 271873 372602 271939 372605
rect 272558 372602 272564 372604
rect 266372 372600 266464 372602
rect 266414 372544 266464 372600
rect 266372 372542 266464 372544
rect 271873 372600 272564 372602
rect 271873 372544 271878 372600
rect 271934 372544 272564 372600
rect 271873 372542 272564 372544
rect 266372 372540 266419 372542
rect 259453 372539 259519 372540
rect 262213 372539 262279 372540
rect 266353 372539 266419 372540
rect 271873 372539 271939 372542
rect 272558 372540 272564 372542
rect 272628 372540 272634 372604
rect 310513 372602 310579 372605
rect 310646 372602 310652 372604
rect 310513 372600 310652 372602
rect 310513 372544 310518 372600
rect 310574 372544 310652 372600
rect 310513 372542 310652 372544
rect 310513 372539 310579 372542
rect 310646 372540 310652 372542
rect 310716 372540 310722 372604
rect 314653 372602 314719 372605
rect 322933 372604 322999 372605
rect 400213 372604 400279 372605
rect 315062 372602 315068 372604
rect 314653 372600 315068 372602
rect 314653 372544 314658 372600
rect 314714 372544 315068 372600
rect 314653 372542 315068 372544
rect 314653 372539 314719 372542
rect 315062 372540 315068 372542
rect 315132 372540 315138 372604
rect 322933 372602 322980 372604
rect 322888 372600 322980 372602
rect 322888 372544 322938 372600
rect 322888 372542 322980 372544
rect 322933 372540 322980 372542
rect 323044 372540 323050 372604
rect 400213 372602 400260 372604
rect 400168 372600 400260 372602
rect 400168 372544 400218 372600
rect 400168 372542 400260 372544
rect 400213 372540 400260 372542
rect 400324 372540 400330 372604
rect 402881 372602 402947 372605
rect 403566 372602 403572 372604
rect 402881 372600 403572 372602
rect 402881 372544 402886 372600
rect 402942 372544 403572 372600
rect 402881 372542 403572 372544
rect 322933 372539 322999 372540
rect 400213 372539 400279 372540
rect 402881 372539 402947 372542
rect 403566 372540 403572 372542
rect 403636 372540 403642 372604
rect 78489 372468 78555 372469
rect 79961 372468 80027 372469
rect 78438 372466 78444 372468
rect 78398 372406 78444 372466
rect 78508 372464 78555 372468
rect 79910 372466 79916 372468
rect 78550 372408 78555 372464
rect 78438 372404 78444 372406
rect 78508 372404 78555 372408
rect 79870 372406 79916 372466
rect 79980 372464 80027 372468
rect 80022 372408 80027 372464
rect 79910 372404 79916 372406
rect 79980 372404 80027 372408
rect 78489 372403 78555 372404
rect 79961 372403 80027 372404
rect 80145 372466 80211 372469
rect 80462 372466 80468 372468
rect 80145 372464 80468 372466
rect 80145 372408 80150 372464
rect 80206 372408 80468 372464
rect 80145 372406 80468 372408
rect 80145 372403 80211 372406
rect 80462 372404 80468 372406
rect 80532 372404 80538 372468
rect 84510 372404 84516 372468
rect 84580 372466 84586 372468
rect 85481 372466 85547 372469
rect 84580 372464 85547 372466
rect 84580 372408 85486 372464
rect 85542 372408 85547 372464
rect 84580 372406 85547 372408
rect 84580 372404 84586 372406
rect 85481 372403 85547 372406
rect 118182 372404 118188 372468
rect 118252 372466 118258 372468
rect 215201 372466 215267 372469
rect 277526 372466 277532 372468
rect 118252 372464 277532 372466
rect 118252 372408 215206 372464
rect 215262 372408 277532 372464
rect 118252 372406 277532 372408
rect 118252 372404 118258 372406
rect 215201 372403 215267 372406
rect 277526 372404 277532 372406
rect 277596 372466 277602 372468
rect 278681 372466 278747 372469
rect 277596 372464 278747 372466
rect 277596 372408 278686 372464
rect 278742 372408 278747 372464
rect 277596 372406 278747 372408
rect 277596 372404 277602 372406
rect 278681 372403 278747 372406
rect 313273 372466 313339 372469
rect 313406 372466 313412 372468
rect 313273 372464 313412 372466
rect 313273 372408 313278 372464
rect 313334 372408 313412 372464
rect 313273 372406 313412 372408
rect 313273 372403 313339 372406
rect 313406 372404 313412 372406
rect 313476 372404 313482 372468
rect 376886 372404 376892 372468
rect 376956 372466 376962 372468
rect 433558 372466 433564 372468
rect 376956 372406 433564 372466
rect 376956 372404 376962 372406
rect 433558 372404 433564 372406
rect 433628 372404 433634 372468
rect 208117 372330 208183 372333
rect 218145 372330 218211 372333
rect 262857 372330 262923 372333
rect 200070 372328 262923 372330
rect 200070 372272 208122 372328
rect 208178 372272 218150 372328
rect 218206 372272 262862 372328
rect 262918 372272 262923 372328
rect 200070 372270 262923 372272
rect 104617 372196 104683 372197
rect 104566 372194 104572 372196
rect 104526 372134 104572 372194
rect 104636 372192 104683 372196
rect 104678 372136 104683 372192
rect 104566 372132 104572 372134
rect 104636 372132 104683 372136
rect 109534 372132 109540 372196
rect 109604 372194 109610 372196
rect 200070 372194 200130 372270
rect 208117 372267 208183 372270
rect 218145 372267 218211 372270
rect 262857 372267 262923 372270
rect 276933 372332 276999 372333
rect 276933 372328 276980 372332
rect 277044 372330 277050 372332
rect 304993 372330 305059 372333
rect 305310 372330 305316 372332
rect 276933 372272 276938 372328
rect 276933 372268 276980 372272
rect 277044 372270 277090 372330
rect 304993 372328 305316 372330
rect 304993 372272 304998 372328
rect 305054 372272 305316 372328
rect 304993 372270 305316 372272
rect 277044 372268 277050 372270
rect 276933 372267 276999 372268
rect 304993 372267 305059 372270
rect 305310 372268 305316 372270
rect 305380 372268 305386 372332
rect 371233 372330 371299 372333
rect 438894 372330 438900 372332
rect 371233 372328 438900 372330
rect 371233 372272 371238 372328
rect 371294 372272 438900 372328
rect 371233 372270 438900 372272
rect 371233 372267 371299 372270
rect 438894 372268 438900 372270
rect 438964 372268 438970 372332
rect 470593 372330 470659 372333
rect 470726 372330 470732 372332
rect 470593 372328 470732 372330
rect 470593 372272 470598 372328
rect 470654 372272 470732 372328
rect 470593 372270 470732 372272
rect 470593 372267 470659 372270
rect 470726 372268 470732 372270
rect 470796 372268 470802 372332
rect 109604 372134 200130 372194
rect 209497 372194 209563 372197
rect 222009 372194 222075 372197
rect 270493 372194 270559 372197
rect 209497 372192 270559 372194
rect 209497 372136 209502 372192
rect 209558 372136 222014 372192
rect 222070 372136 270498 372192
rect 270554 372136 270559 372192
rect 209497 372134 270559 372136
rect 109604 372132 109610 372134
rect 104617 372131 104683 372132
rect 209497 372131 209563 372134
rect 222009 372131 222075 372134
rect 270493 372131 270559 372134
rect 396073 372194 396139 372197
rect 503161 372196 503227 372197
rect 503529 372196 503595 372197
rect 396206 372194 396212 372196
rect 396073 372192 396212 372194
rect 396073 372136 396078 372192
rect 396134 372136 396212 372192
rect 396073 372134 396212 372136
rect 396073 372131 396139 372134
rect 396206 372132 396212 372134
rect 396276 372132 396282 372196
rect 503110 372194 503116 372196
rect 503070 372134 503116 372194
rect 503180 372192 503227 372196
rect 503478 372194 503484 372196
rect 503222 372136 503227 372192
rect 503110 372132 503116 372134
rect 503180 372132 503227 372136
rect 503438 372134 503484 372194
rect 503548 372192 503595 372196
rect 503590 372136 503595 372192
rect 503478 372132 503484 372134
rect 503548 372132 503595 372136
rect 503161 372131 503227 372132
rect 503529 372131 503595 372132
rect 113214 371996 113220 372060
rect 113284 372058 113290 372060
rect 214925 372058 214991 372061
rect 219525 372058 219591 372061
rect 397453 372060 397519 372061
rect 273294 372058 273300 372060
rect 113284 372056 273300 372058
rect 113284 372000 214930 372056
rect 214986 372000 219530 372056
rect 219586 372000 273300 372056
rect 113284 371998 273300 372000
rect 113284 371996 113290 371998
rect 214925 371995 214991 371998
rect 219525 371995 219591 371998
rect 273294 371996 273300 371998
rect 273364 371996 273370 372060
rect 397453 372058 397500 372060
rect 397408 372056 397500 372058
rect 397408 372000 397458 372056
rect 397408 371998 397500 372000
rect 397453 371996 397500 371998
rect 397564 371996 397570 372060
rect 404353 372058 404419 372061
rect 404854 372058 404860 372060
rect 404353 372056 404860 372058
rect 404353 372000 404358 372056
rect 404414 372000 404860 372056
rect 404353 371998 404860 372000
rect 397453 371995 397519 371996
rect 404353 371995 404419 371998
rect 404854 371996 404860 371998
rect 404924 371996 404930 372060
rect 407113 372058 407179 372061
rect 422293 372060 422359 372061
rect 407246 372058 407252 372060
rect 407113 372056 407252 372058
rect 407113 372000 407118 372056
rect 407174 372000 407252 372056
rect 407113 371998 407252 372000
rect 407113 371995 407179 371998
rect 407246 371996 407252 371998
rect 407316 371996 407322 372060
rect 422293 372056 422340 372060
rect 422404 372058 422410 372060
rect 422293 372000 422298 372056
rect 422293 371996 422340 372000
rect 422404 371998 422450 372058
rect 422404 371996 422410 371998
rect 422293 371995 422359 371996
rect 76598 371860 76604 371924
rect 76668 371922 76674 371924
rect 77017 371922 77083 371925
rect 76668 371920 77083 371922
rect 76668 371864 77022 371920
rect 77078 371864 77083 371920
rect 76668 371862 77083 371864
rect 76668 371860 76674 371862
rect 77017 371859 77083 371862
rect 108982 371860 108988 371924
rect 109052 371922 109058 371924
rect 209589 371922 209655 371925
rect 221917 371922 221983 371925
rect 270217 371922 270283 371925
rect 109052 371920 209655 371922
rect 109052 371864 209594 371920
rect 209650 371864 209655 371920
rect 109052 371862 209655 371864
rect 109052 371860 109058 371862
rect 209589 371859 209655 371862
rect 215250 371920 270283 371922
rect 215250 371864 221922 371920
rect 221978 371864 270222 371920
rect 270278 371864 270283 371920
rect 215250 371862 270283 371864
rect 115790 371724 115796 371788
rect 115860 371786 115866 371788
rect 211705 371786 211771 371789
rect 215250 371786 215310 371862
rect 221917 371859 221983 371862
rect 270217 371859 270283 371862
rect 377397 371922 377463 371925
rect 377806 371922 377812 371924
rect 377397 371920 377812 371922
rect 377397 371864 377402 371920
rect 377458 371864 377812 371920
rect 377397 371862 377812 371864
rect 377397 371859 377463 371862
rect 377806 371860 377812 371862
rect 377876 371922 377882 371924
rect 438342 371922 438348 371924
rect 377876 371862 438348 371922
rect 377876 371860 377882 371862
rect 438342 371860 438348 371862
rect 438412 371860 438418 371924
rect 483013 371922 483079 371925
rect 483238 371922 483244 371924
rect 483013 371920 483244 371922
rect 483013 371864 483018 371920
rect 483074 371864 483244 371920
rect 483013 371862 483244 371864
rect 483013 371859 483079 371862
rect 483238 371860 483244 371862
rect 483308 371860 483314 371924
rect 115860 371784 215310 371786
rect 115860 371728 211710 371784
rect 211766 371728 215310 371784
rect 115860 371726 215310 371728
rect 245653 371786 245719 371789
rect 245878 371786 245884 371788
rect 245653 371784 245884 371786
rect 245653 371728 245658 371784
rect 245714 371728 245884 371784
rect 245653 371726 245884 371728
rect 115860 371724 115866 371726
rect 211705 371723 211771 371726
rect 245653 371723 245719 371726
rect 245878 371724 245884 371726
rect 245948 371724 245954 371788
rect 273437 371786 273503 371789
rect 273662 371786 273668 371788
rect 273437 371784 273668 371786
rect 273437 371728 273442 371784
rect 273498 371728 273668 371784
rect 273437 371726 273668 371728
rect 273437 371723 273503 371726
rect 273662 371724 273668 371726
rect 273732 371724 273738 371788
rect 317413 371786 317479 371789
rect 317822 371786 317828 371788
rect 317413 371784 317828 371786
rect 317413 371728 317418 371784
rect 317474 371728 317828 371784
rect 317413 371726 317828 371728
rect 317413 371723 317479 371726
rect 317822 371724 317828 371726
rect 317892 371724 317898 371788
rect 401593 371786 401659 371789
rect 402278 371786 402284 371788
rect 401593 371784 402284 371786
rect 401593 371728 401598 371784
rect 401654 371728 402284 371784
rect 401593 371726 402284 371728
rect 401593 371723 401659 371726
rect 402278 371724 402284 371726
rect 402348 371724 402354 371788
rect 409873 371786 409939 371789
rect 410006 371786 410012 371788
rect 409873 371784 410012 371786
rect 409873 371728 409878 371784
rect 409934 371728 410012 371784
rect 409873 371726 410012 371728
rect 409873 371723 409939 371726
rect 410006 371724 410012 371726
rect 410076 371724 410082 371788
rect 95233 371652 95299 371653
rect 95182 371650 95188 371652
rect 95142 371590 95188 371650
rect 95252 371648 95299 371652
rect 95294 371592 95299 371648
rect 95182 371588 95188 371590
rect 95252 371588 95299 371592
rect 98126 371588 98132 371652
rect 98196 371650 98202 371652
rect 99281 371650 99347 371653
rect 98196 371648 99347 371650
rect 98196 371592 99286 371648
rect 99342 371592 99347 371648
rect 98196 371590 99347 371592
rect 98196 371588 98202 371590
rect 95233 371587 95299 371588
rect 99281 371587 99347 371590
rect 99966 371588 99972 371652
rect 100036 371650 100042 371652
rect 100477 371650 100543 371653
rect 100036 371648 100543 371650
rect 100036 371592 100482 371648
rect 100538 371592 100543 371648
rect 100036 371590 100543 371592
rect 100036 371588 100042 371590
rect 100477 371587 100543 371590
rect 105302 371588 105308 371652
rect 105372 371650 105378 371652
rect 106089 371650 106155 371653
rect 105372 371648 106155 371650
rect 105372 371592 106094 371648
rect 106150 371592 106155 371648
rect 105372 371590 106155 371592
rect 105372 371588 105378 371590
rect 106089 371587 106155 371590
rect 182817 371650 182883 371653
rect 182950 371650 182956 371652
rect 182817 371648 182956 371650
rect 182817 371592 182822 371648
rect 182878 371592 182956 371648
rect 182817 371590 182956 371592
rect 182817 371587 182883 371590
rect 182950 371588 182956 371590
rect 183020 371588 183026 371652
rect 183318 371588 183324 371652
rect 183388 371650 183394 371652
rect 183461 371650 183527 371653
rect 183388 371648 183527 371650
rect 183388 371592 183466 371648
rect 183522 371592 183527 371648
rect 183388 371590 183527 371592
rect 183388 371588 183394 371590
rect 183461 371587 183527 371590
rect 209589 371650 209655 371653
rect 217542 371650 217548 371652
rect 209589 371648 217548 371650
rect 209589 371592 209594 371648
rect 209650 371592 217548 371648
rect 209589 371590 217548 371592
rect 209589 371587 209655 371590
rect 217542 371588 217548 371590
rect 217612 371650 217618 371652
rect 262765 371650 262831 371653
rect 217612 371648 262831 371650
rect 217612 371592 262770 371648
rect 262826 371592 262831 371648
rect 217612 371590 262831 371592
rect 217612 371588 217618 371590
rect 262765 371587 262831 371590
rect 398833 371650 398899 371653
rect 411253 371652 411319 371653
rect 398966 371650 398972 371652
rect 398833 371648 398972 371650
rect 398833 371592 398838 371648
rect 398894 371592 398972 371648
rect 398833 371590 398972 371592
rect 398833 371587 398899 371590
rect 398966 371588 398972 371590
rect 399036 371588 399042 371652
rect 411253 371650 411300 371652
rect 411208 371648 411300 371650
rect 411208 371592 411258 371648
rect 411208 371590 411300 371592
rect 411253 371588 411300 371590
rect 411364 371588 411370 371652
rect 465073 371650 465139 371653
rect 465390 371650 465396 371652
rect 465073 371648 465396 371650
rect 465073 371592 465078 371648
rect 465134 371592 465396 371648
rect 465073 371590 465396 371592
rect 411253 371587 411319 371588
rect 465073 371587 465139 371590
rect 465390 371588 465396 371590
rect 465460 371588 465466 371652
rect -960 371228 480 371468
rect 97574 371452 97580 371516
rect 97644 371514 97650 371516
rect 97717 371514 97783 371517
rect 97644 371512 97783 371514
rect 97644 371456 97722 371512
rect 97778 371456 97783 371512
rect 97644 371454 97783 371456
rect 97644 371452 97650 371454
rect 97717 371451 97783 371454
rect 100702 371452 100708 371516
rect 100772 371514 100778 371516
rect 101121 371514 101187 371517
rect 100772 371512 101187 371514
rect 100772 371456 101126 371512
rect 101182 371456 101187 371512
rect 100772 371454 101187 371456
rect 100772 371452 100778 371454
rect 101121 371451 101187 371454
rect 111742 371452 111748 371516
rect 111812 371514 111818 371516
rect 209497 371514 209563 371517
rect 276013 371514 276079 371517
rect 111812 371512 209563 371514
rect 111812 371456 209502 371512
rect 209558 371456 209563 371512
rect 111812 371454 209563 371456
rect 111812 371452 111818 371454
rect 209497 371451 209563 371454
rect 219390 371512 276079 371514
rect 219390 371456 276018 371512
rect 276074 371456 276079 371512
rect 219390 371454 276079 371456
rect 55673 371378 55739 371381
rect 107561 371380 107627 371381
rect 57094 371378 57100 371380
rect 55673 371376 57100 371378
rect 55673 371320 55678 371376
rect 55734 371320 57100 371376
rect 55673 371318 57100 371320
rect 55673 371315 55739 371318
rect 57094 371316 57100 371318
rect 57164 371316 57170 371380
rect 102726 371316 102732 371380
rect 102796 371316 102802 371380
rect 107510 371378 107516 371380
rect 107470 371318 107516 371378
rect 107580 371376 107627 371380
rect 107622 371320 107627 371376
rect 107510 371316 107516 371318
rect 107580 371316 107627 371320
rect 117078 371316 117084 371380
rect 117148 371378 117154 371380
rect 216581 371378 216647 371381
rect 219390 371378 219450 371454
rect 276013 371451 276079 371454
rect 277669 371514 277735 371517
rect 278262 371514 278268 371516
rect 277669 371512 278268 371514
rect 277669 371456 277674 371512
rect 277730 371456 278268 371512
rect 277669 371454 278268 371456
rect 277669 371451 277735 371454
rect 278262 371452 278268 371454
rect 278332 371452 278338 371516
rect 411345 371514 411411 371517
rect 411846 371514 411852 371516
rect 411345 371512 411852 371514
rect 411345 371456 411350 371512
rect 411406 371456 411852 371512
rect 411345 371454 411852 371456
rect 411345 371451 411411 371454
rect 411846 371452 411852 371454
rect 411916 371452 411922 371516
rect 418245 371514 418311 371517
rect 418838 371514 418844 371516
rect 418245 371512 418844 371514
rect 418245 371456 418250 371512
rect 418306 371456 418844 371512
rect 418245 371454 418844 371456
rect 418245 371451 418311 371454
rect 418838 371452 418844 371454
rect 418908 371452 418914 371516
rect 421005 371514 421071 371517
rect 421230 371514 421236 371516
rect 421005 371512 421236 371514
rect 421005 371456 421010 371512
rect 421066 371456 421236 371512
rect 421005 371454 421236 371456
rect 421005 371451 421071 371454
rect 421230 371452 421236 371454
rect 421300 371452 421306 371516
rect 423673 371514 423739 371517
rect 426433 371516 426499 371517
rect 423990 371514 423996 371516
rect 423673 371512 423996 371514
rect 423673 371456 423678 371512
rect 423734 371456 423996 371512
rect 423673 371454 423996 371456
rect 423673 371451 423739 371454
rect 423990 371452 423996 371454
rect 424060 371452 424066 371516
rect 426382 371452 426388 371516
rect 426452 371514 426499 371516
rect 430665 371514 430731 371517
rect 431166 371514 431172 371516
rect 426452 371512 426544 371514
rect 426494 371456 426544 371512
rect 426452 371454 426544 371456
rect 430665 371512 431172 371514
rect 430665 371456 430670 371512
rect 430726 371456 431172 371512
rect 430665 371454 431172 371456
rect 426452 371452 426499 371454
rect 426433 371451 426499 371452
rect 430665 371451 430731 371454
rect 431166 371452 431172 371454
rect 431236 371452 431242 371516
rect 117148 371376 219450 371378
rect 117148 371320 216586 371376
rect 216642 371320 219450 371376
rect 117148 371318 219450 371320
rect 247033 371378 247099 371381
rect 247902 371378 247908 371380
rect 247033 371376 247908 371378
rect 247033 371320 247038 371376
rect 247094 371320 247908 371376
rect 247033 371318 247908 371320
rect 117148 371316 117154 371318
rect 102734 371242 102794 371316
rect 107561 371315 107627 371316
rect 216581 371315 216647 371318
rect 247033 371315 247099 371318
rect 247902 371316 247908 371318
rect 247972 371316 247978 371380
rect 252553 371378 252619 371381
rect 253606 371378 253612 371380
rect 252553 371376 253612 371378
rect 252553 371320 252558 371376
rect 252614 371320 253612 371376
rect 252553 371318 253612 371320
rect 252553 371315 252619 371318
rect 253606 371316 253612 371318
rect 253676 371316 253682 371380
rect 258165 371378 258231 371381
rect 258390 371378 258396 371380
rect 258165 371376 258396 371378
rect 258165 371320 258170 371376
rect 258226 371320 258396 371376
rect 258165 371318 258396 371320
rect 258165 371315 258231 371318
rect 258390 371316 258396 371318
rect 258460 371316 258466 371380
rect 260833 371378 260899 371381
rect 263593 371380 263659 371381
rect 260966 371378 260972 371380
rect 260833 371376 260972 371378
rect 260833 371320 260838 371376
rect 260894 371320 260972 371376
rect 260833 371318 260972 371320
rect 260833 371315 260899 371318
rect 260966 371316 260972 371318
rect 261036 371316 261042 371380
rect 263542 371316 263548 371380
rect 263612 371378 263659 371380
rect 264973 371378 265039 371381
rect 265750 371378 265756 371380
rect 263612 371376 263704 371378
rect 263654 371320 263704 371376
rect 263612 371318 263704 371320
rect 264973 371376 265756 371378
rect 264973 371320 264978 371376
rect 265034 371320 265756 371376
rect 264973 371318 265756 371320
rect 263612 371316 263659 371318
rect 263593 371315 263659 371316
rect 264973 371315 265039 371318
rect 265750 371316 265756 371318
rect 265820 371316 265826 371380
rect 266353 371378 266419 371381
rect 267733 371380 267799 371381
rect 267038 371378 267044 371380
rect 266353 371376 267044 371378
rect 266353 371320 266358 371376
rect 266414 371320 267044 371376
rect 266353 371318 267044 371320
rect 266353 371315 266419 371318
rect 267038 371316 267044 371318
rect 267108 371316 267114 371380
rect 267733 371376 267780 371380
rect 267844 371378 267850 371380
rect 270493 371378 270559 371381
rect 270902 371378 270908 371380
rect 267733 371320 267738 371376
rect 267733 371316 267780 371320
rect 267844 371318 267890 371378
rect 270493 371376 270908 371378
rect 270493 371320 270498 371376
rect 270554 371320 270908 371376
rect 270493 371318 270908 371320
rect 267844 371316 267850 371318
rect 267733 371315 267799 371316
rect 270493 371315 270559 371318
rect 270902 371316 270908 371318
rect 270972 371316 270978 371380
rect 273253 371378 273319 371381
rect 273846 371378 273852 371380
rect 273253 371376 273852 371378
rect 273253 371320 273258 371376
rect 273314 371320 273852 371376
rect 273253 371318 273852 371320
rect 273253 371315 273319 371318
rect 273846 371316 273852 371318
rect 273916 371316 273922 371380
rect 276013 371378 276079 371381
rect 276238 371378 276244 371380
rect 276013 371376 276244 371378
rect 276013 371320 276018 371376
rect 276074 371320 276244 371376
rect 276013 371318 276244 371320
rect 276013 371315 276079 371318
rect 276238 371316 276244 371318
rect 276308 371316 276314 371380
rect 280153 371378 280219 371381
rect 280286 371378 280292 371380
rect 280153 371376 280292 371378
rect 280153 371320 280158 371376
rect 280214 371320 280292 371376
rect 280153 371318 280292 371320
rect 280153 371315 280219 371318
rect 280286 371316 280292 371318
rect 280356 371316 280362 371380
rect 282913 371378 282979 371381
rect 283782 371378 283788 371380
rect 282913 371376 283788 371378
rect 282913 371320 282918 371376
rect 282974 371320 283788 371376
rect 282913 371318 283788 371320
rect 282913 371315 282979 371318
rect 283782 371316 283788 371318
rect 283852 371316 283858 371380
rect 285673 371378 285739 371381
rect 285806 371378 285812 371380
rect 285673 371376 285812 371378
rect 285673 371320 285678 371376
rect 285734 371320 285812 371376
rect 285673 371318 285812 371320
rect 285673 371315 285739 371318
rect 285806 371316 285812 371318
rect 285876 371316 285882 371380
rect 287329 371378 287395 371381
rect 287646 371378 287652 371380
rect 287329 371376 287652 371378
rect 287329 371320 287334 371376
rect 287390 371320 287652 371376
rect 287329 371318 287652 371320
rect 287329 371315 287395 371318
rect 287646 371316 287652 371318
rect 287716 371316 287722 371380
rect 289813 371378 289879 371381
rect 290590 371378 290596 371380
rect 289813 371376 290596 371378
rect 289813 371320 289818 371376
rect 289874 371320 290596 371376
rect 289813 371318 290596 371320
rect 289813 371315 289879 371318
rect 290590 371316 290596 371318
rect 290660 371316 290666 371380
rect 292573 371378 292639 371381
rect 295333 371380 295399 371381
rect 298093 371380 298159 371381
rect 292798 371378 292804 371380
rect 292573 371376 292804 371378
rect 292573 371320 292578 371376
rect 292634 371320 292804 371376
rect 292573 371318 292804 371320
rect 292573 371315 292639 371318
rect 292798 371316 292804 371318
rect 292868 371316 292874 371380
rect 295333 371378 295380 371380
rect 295288 371376 295380 371378
rect 295288 371320 295338 371376
rect 295288 371318 295380 371320
rect 295333 371316 295380 371318
rect 295444 371316 295450 371380
rect 298093 371378 298140 371380
rect 298048 371376 298140 371378
rect 298048 371320 298098 371376
rect 298048 371318 298140 371320
rect 298093 371316 298140 371318
rect 298204 371316 298210 371380
rect 302233 371378 302299 371381
rect 302918 371378 302924 371380
rect 302233 371376 302924 371378
rect 302233 371320 302238 371376
rect 302294 371320 302924 371376
rect 302233 371318 302924 371320
rect 295333 371315 295399 371316
rect 298093 371315 298159 371316
rect 302233 371315 302299 371318
rect 302918 371316 302924 371318
rect 302988 371316 302994 371380
rect 307753 371378 307819 371381
rect 308622 371378 308628 371380
rect 307753 371376 308628 371378
rect 307753 371320 307758 371376
rect 307814 371320 308628 371376
rect 307753 371318 308628 371320
rect 307753 371315 307819 371318
rect 308622 371316 308628 371318
rect 308692 371316 308698 371380
rect 326153 371378 326219 371381
rect 326654 371378 326660 371380
rect 326153 371376 326660 371378
rect 326153 371320 326158 371376
rect 326214 371320 326660 371376
rect 326153 371318 326660 371320
rect 326153 371315 326219 371318
rect 326654 371316 326660 371318
rect 326724 371316 326730 371380
rect 342897 371378 342963 371381
rect 343357 371380 343423 371381
rect 343030 371378 343036 371380
rect 342897 371376 343036 371378
rect 342897 371320 342902 371376
rect 342958 371320 343036 371376
rect 342897 371318 343036 371320
rect 342897 371315 342963 371318
rect 343030 371316 343036 371318
rect 343100 371316 343106 371380
rect 343357 371376 343404 371380
rect 343468 371378 343474 371380
rect 396073 371378 396139 371381
rect 402973 371380 403039 371381
rect 396574 371378 396580 371380
rect 343357 371320 343362 371376
rect 343357 371316 343404 371320
rect 343468 371318 343514 371378
rect 396073 371376 396580 371378
rect 396073 371320 396078 371376
rect 396134 371320 396580 371376
rect 396073 371318 396580 371320
rect 343468 371316 343474 371318
rect 343357 371315 343423 371316
rect 396073 371315 396139 371318
rect 396574 371316 396580 371318
rect 396644 371316 396650 371380
rect 402973 371376 403020 371380
rect 403084 371378 403090 371380
rect 412633 371378 412699 371381
rect 412766 371378 412772 371380
rect 402973 371320 402978 371376
rect 402973 371316 403020 371320
rect 403084 371318 403130 371378
rect 412633 371376 412772 371378
rect 412633 371320 412638 371376
rect 412694 371320 412772 371376
rect 412633 371318 412772 371320
rect 403084 371316 403090 371318
rect 402973 371315 403039 371316
rect 412633 371315 412699 371318
rect 412766 371316 412772 371318
rect 412836 371316 412842 371380
rect 413185 371378 413251 371381
rect 414013 371380 414079 371381
rect 413686 371378 413692 371380
rect 413185 371376 413692 371378
rect 413185 371320 413190 371376
rect 413246 371320 413692 371376
rect 413185 371318 413692 371320
rect 413185 371315 413251 371318
rect 413686 371316 413692 371318
rect 413756 371316 413762 371380
rect 414013 371378 414060 371380
rect 413968 371376 414060 371378
rect 413968 371320 414018 371376
rect 413968 371318 414060 371320
rect 414013 371316 414060 371318
rect 414124 371316 414130 371380
rect 415393 371378 415459 371381
rect 416773 371380 416839 371381
rect 418153 371380 418219 371381
rect 415526 371378 415532 371380
rect 415393 371376 415532 371378
rect 415393 371320 415398 371376
rect 415454 371320 415532 371376
rect 415393 371318 415532 371320
rect 414013 371315 414079 371316
rect 415393 371315 415459 371318
rect 415526 371316 415532 371318
rect 415596 371316 415602 371380
rect 416773 371378 416820 371380
rect 416728 371376 416820 371378
rect 416728 371320 416778 371376
rect 416728 371318 416820 371320
rect 416773 371316 416820 371318
rect 416884 371316 416890 371380
rect 418102 371316 418108 371380
rect 418172 371378 418219 371380
rect 419533 371378 419599 371381
rect 420310 371378 420316 371380
rect 418172 371376 418264 371378
rect 418214 371320 418264 371376
rect 418172 371318 418264 371320
rect 419533 371376 420316 371378
rect 419533 371320 419538 371376
rect 419594 371320 420316 371376
rect 419533 371318 420316 371320
rect 418172 371316 418219 371318
rect 416773 371315 416839 371316
rect 418153 371315 418219 371316
rect 419533 371315 419599 371318
rect 420310 371316 420316 371318
rect 420380 371316 420386 371380
rect 420913 371378 420979 371381
rect 421046 371378 421052 371380
rect 420913 371376 421052 371378
rect 420913 371320 420918 371376
rect 420974 371320 421052 371376
rect 420913 371318 421052 371320
rect 420913 371315 420979 371318
rect 421046 371316 421052 371318
rect 421116 371316 421122 371380
rect 425053 371378 425119 371381
rect 425646 371378 425652 371380
rect 425053 371376 425652 371378
rect 425053 371320 425058 371376
rect 425114 371320 425652 371376
rect 425053 371318 425652 371320
rect 425053 371315 425119 371318
rect 425646 371316 425652 371318
rect 425716 371316 425722 371380
rect 427813 371378 427879 371381
rect 428590 371378 428596 371380
rect 427813 371376 428596 371378
rect 427813 371320 427818 371376
rect 427874 371320 428596 371376
rect 427813 371318 428596 371320
rect 427813 371315 427879 371318
rect 428590 371316 428596 371318
rect 428660 371316 428666 371380
rect 429193 371378 429259 371381
rect 430573 371380 430639 371381
rect 429326 371378 429332 371380
rect 429193 371376 429332 371378
rect 429193 371320 429198 371376
rect 429254 371320 429332 371376
rect 429193 371318 429332 371320
rect 429193 371315 429259 371318
rect 429326 371316 429332 371318
rect 429396 371316 429402 371380
rect 430573 371378 430620 371380
rect 430528 371376 430620 371378
rect 430528 371320 430578 371376
rect 430528 371318 430620 371320
rect 430573 371316 430620 371318
rect 430684 371316 430690 371380
rect 431953 371378 432019 371381
rect 433333 371380 433399 371381
rect 432086 371378 432092 371380
rect 431953 371376 432092 371378
rect 431953 371320 431958 371376
rect 432014 371320 432092 371376
rect 431953 371318 432092 371320
rect 430573 371315 430639 371316
rect 431953 371315 432019 371318
rect 432086 371316 432092 371318
rect 432156 371316 432162 371380
rect 433333 371378 433380 371380
rect 433288 371376 433380 371378
rect 433288 371320 433338 371376
rect 433288 371318 433380 371320
rect 433333 371316 433380 371318
rect 433444 371316 433450 371380
rect 434713 371378 434779 371381
rect 434846 371378 434852 371380
rect 434713 371376 434852 371378
rect 434713 371320 434718 371376
rect 434774 371320 434852 371376
rect 434713 371318 434852 371320
rect 433333 371315 433399 371316
rect 434713 371315 434779 371318
rect 434846 371316 434852 371318
rect 434916 371316 434922 371380
rect 436093 371378 436159 371381
rect 458173 371380 458239 371381
rect 473353 371380 473419 371381
rect 436318 371378 436324 371380
rect 436093 371376 436324 371378
rect 436093 371320 436098 371376
rect 436154 371320 436324 371376
rect 436093 371318 436324 371320
rect 436093 371315 436159 371318
rect 436318 371316 436324 371318
rect 436388 371316 436394 371380
rect 458173 371378 458220 371380
rect 458128 371376 458220 371378
rect 458128 371320 458178 371376
rect 458128 371318 458220 371320
rect 458173 371316 458220 371318
rect 458284 371316 458290 371380
rect 473302 371316 473308 371380
rect 473372 371378 473419 371380
rect 474733 371378 474799 371381
rect 475326 371378 475332 371380
rect 473372 371376 473464 371378
rect 473414 371320 473464 371376
rect 473372 371318 473464 371320
rect 474733 371376 475332 371378
rect 474733 371320 474738 371376
rect 474794 371320 475332 371376
rect 474733 371318 475332 371320
rect 473372 371316 473419 371318
rect 458173 371315 458239 371316
rect 473353 371315 473419 371316
rect 474733 371315 474799 371318
rect 475326 371316 475332 371318
rect 475396 371316 475402 371380
rect 477493 371378 477559 371381
rect 480253 371380 480319 371381
rect 478086 371378 478092 371380
rect 477493 371376 478092 371378
rect 477493 371320 477498 371376
rect 477554 371320 478092 371376
rect 477493 371318 478092 371320
rect 477493 371315 477559 371318
rect 478086 371316 478092 371318
rect 478156 371316 478162 371380
rect 480253 371376 480300 371380
rect 480364 371378 480370 371380
rect 480253 371320 480258 371376
rect 480253 371316 480300 371320
rect 480364 371318 480410 371378
rect 480364 371316 480370 371318
rect 480253 371315 480319 371316
rect 215385 371242 215451 371245
rect 102734 371240 215451 371242
rect 102734 371184 215390 371240
rect 215446 371184 215451 371240
rect 102734 371182 215451 371184
rect 215385 371179 215451 371182
rect 359774 371180 359780 371244
rect 359844 371242 359850 371244
rect 467966 371242 467972 371244
rect 359844 371182 467972 371242
rect 359844 371180 359850 371182
rect 467966 371180 467972 371182
rect 468036 371180 468042 371244
rect 106406 371044 106412 371108
rect 106476 371106 106482 371108
rect 216990 371106 216996 371108
rect 106476 371046 216996 371106
rect 106476 371044 106482 371046
rect 216990 371044 216996 371046
rect 217060 371044 217066 371108
rect 95233 369746 95299 369749
rect 212625 369746 212691 369749
rect 95233 369744 212691 369746
rect 95233 369688 95238 369744
rect 95294 369688 212630 369744
rect 212686 369688 212691 369744
rect 95233 369686 212691 369688
rect 95233 369683 95299 369686
rect 212625 369683 212691 369686
rect 104617 369610 104683 369613
rect 215845 369610 215911 369613
rect 104617 369608 215911 369610
rect 104617 369552 104622 369608
rect 104678 369552 215850 369608
rect 215906 369552 215911 369608
rect 104617 369550 215911 369552
rect 104617 369547 104683 369550
rect 215845 369547 215911 369550
rect 212758 369140 212764 369204
rect 212828 369202 212834 369204
rect 213821 369202 213887 369205
rect 212828 369200 213887 369202
rect 212828 369144 213826 369200
rect 213882 369144 213887 369200
rect 212828 369142 213887 369144
rect 212828 369140 212834 369142
rect 213821 369139 213887 369142
rect 215518 369140 215524 369204
rect 215588 369202 215594 369204
rect 216581 369202 216647 369205
rect 215588 369200 216647 369202
rect 215588 369144 216586 369200
rect 216642 369144 216647 369200
rect 215588 369142 216647 369144
rect 215588 369140 215594 369142
rect 216581 369139 216647 369142
rect 376937 368524 377003 368525
rect 376886 368522 376892 368524
rect 376846 368462 376892 368522
rect 376956 368520 377003 368524
rect 376998 368464 377003 368520
rect 376886 368460 376892 368462
rect 376956 368460 377003 368464
rect 376937 368459 377003 368460
rect 214833 368386 214899 368389
rect 217358 368386 217364 368388
rect 214833 368384 217364 368386
rect 214833 368328 214838 368384
rect 214894 368328 217364 368384
rect 214833 368326 217364 368328
rect 214833 368323 214899 368326
rect 217358 368324 217364 368326
rect 217428 368386 217434 368388
rect 266353 368386 266419 368389
rect 217428 368384 266419 368386
rect 217428 368328 266358 368384
rect 266414 368328 266419 368384
rect 217428 368326 266419 368328
rect 217428 368324 217434 368326
rect 266353 368323 266419 368326
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 199510 357988 199516 358052
rect 199580 358050 199586 358052
rect 199745 358050 199811 358053
rect 359273 358050 359339 358053
rect 519353 358050 519419 358053
rect 199580 358048 519419 358050
rect 199580 357992 199750 358048
rect 199806 357992 359278 358048
rect 359334 357992 519358 358048
rect 519414 357992 519419 358048
rect 199580 357990 519419 357992
rect 199580 357988 199586 357990
rect 199745 357987 199811 357990
rect 359273 357987 359339 357990
rect 519353 357987 519419 357990
rect 178534 355268 178540 355332
rect 178604 355330 178610 355332
rect 179137 355330 179203 355333
rect 178604 355328 179203 355330
rect 178604 355272 179142 355328
rect 179198 355272 179203 355328
rect 178604 355270 179203 355272
rect 178604 355268 178610 355270
rect 179137 355267 179203 355270
rect 190862 355268 190868 355332
rect 190932 355330 190938 355332
rect 191465 355330 191531 355333
rect 190932 355328 191531 355330
rect 190932 355272 191470 355328
rect 191526 355272 191531 355328
rect 190932 355270 191531 355272
rect 190932 355268 190938 355270
rect 191465 355267 191531 355270
rect 338481 355060 338547 355061
rect 338430 355058 338436 355060
rect 338390 354998 338436 355058
rect 338500 355056 338547 355060
rect 338542 355000 338547 355056
rect 338430 354996 338436 354998
rect 338500 354996 338547 355000
rect 350942 354996 350948 355060
rect 351012 355058 351018 355060
rect 351729 355058 351795 355061
rect 351012 355056 351795 355058
rect 351012 355000 351734 355056
rect 351790 355000 351795 355056
rect 351012 354998 351795 355000
rect 351012 354996 351018 354998
rect 338481 354995 338547 354996
rect 351729 354995 351795 354998
rect 498510 354996 498516 355060
rect 498580 355058 498586 355060
rect 498837 355058 498903 355061
rect 498580 355056 498903 355058
rect 498580 355000 498842 355056
rect 498898 355000 498903 355056
rect 498580 354998 498903 355000
rect 498580 354996 498586 354998
rect 498837 354995 498903 354998
rect 499798 354860 499804 354924
rect 499868 354922 499874 354924
rect 500861 354922 500927 354925
rect 499868 354920 500927 354922
rect 499868 354864 500866 354920
rect 500922 354864 500927 354920
rect 499868 354862 500927 354864
rect 499868 354860 499874 354862
rect 500861 354859 500927 354862
rect 179689 354788 179755 354789
rect 339769 354788 339835 354789
rect 510889 354788 510955 354789
rect 179638 354786 179644 354788
rect 179598 354726 179644 354786
rect 179708 354784 179755 354788
rect 339718 354786 339724 354788
rect 179750 354728 179755 354784
rect 179638 354724 179644 354726
rect 179708 354724 179755 354728
rect 339678 354726 339724 354786
rect 339788 354784 339835 354788
rect 510838 354786 510844 354788
rect 339830 354728 339835 354784
rect 339718 354724 339724 354726
rect 339788 354724 339835 354728
rect 510798 354726 510844 354786
rect 510908 354784 510955 354788
rect 510950 354728 510955 354784
rect 510838 354724 510844 354726
rect 510908 354724 510955 354728
rect 179689 354723 179755 354724
rect 339769 354723 339835 354724
rect 510889 354723 510955 354724
rect 217358 353364 217364 353428
rect 217428 353426 217434 353428
rect 220997 353426 221063 353429
rect 217428 353424 221063 353426
rect 217428 353368 221002 353424
rect 221058 353368 221063 353424
rect 217428 353366 221063 353368
rect 217428 353364 217434 353366
rect 220997 353363 221063 353366
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect 198733 349618 198799 349621
rect 199009 349618 199075 349621
rect 358905 349618 358971 349621
rect 196558 349616 199075 349618
rect 196558 349560 198738 349616
rect 198794 349560 199014 349616
rect 199070 349560 199075 349616
rect 196558 349558 199075 349560
rect 196558 349190 196618 349558
rect 198733 349555 198799 349558
rect 199009 349555 199075 349558
rect 356562 349616 358971 349618
rect 356562 349560 358910 349616
rect 358966 349560 358971 349616
rect 356562 349558 358971 349560
rect 356562 349190 356622 349558
rect 358905 349555 358971 349558
rect 518893 349210 518959 349213
rect 516558 349208 518959 349210
rect 516558 349152 518898 349208
rect 518954 349152 518959 349208
rect 516558 349150 518959 349152
rect 518893 349147 518959 349150
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect 57145 307730 57211 307733
rect 57513 307730 57579 307733
rect 57145 307728 57579 307730
rect 57145 307672 57150 307728
rect 57206 307672 57518 307728
rect 57574 307672 57579 307728
rect 57145 307670 57579 307672
rect 57145 307667 57211 307670
rect 57513 307667 57579 307670
rect 216673 307730 216739 307733
rect 217777 307730 217843 307733
rect 216673 307728 217843 307730
rect 216673 307672 216678 307728
rect 216734 307672 217782 307728
rect 217838 307672 217843 307728
rect 216673 307670 217843 307672
rect 216673 307667 216739 307670
rect 217777 307667 217843 307670
rect 376845 307730 376911 307733
rect 377581 307730 377647 307733
rect 376845 307728 377647 307730
rect 376845 307672 376850 307728
rect 376906 307672 377586 307728
rect 377642 307672 377647 307728
rect 376845 307670 377647 307672
rect 376845 307667 376911 307670
rect 377581 307667 377647 307670
rect 57145 306914 57211 306917
rect 217777 306914 217843 306917
rect 219390 306914 220064 306924
rect 57145 306912 60062 306914
rect 57145 306856 57150 306912
rect 57206 306856 60062 306912
rect 57145 306854 60062 306856
rect 217777 306912 220064 306914
rect 217777 306856 217782 306912
rect 217838 306864 220064 306912
rect 376845 306914 376911 306917
rect 379470 306914 380052 306924
rect 376845 306912 380052 306914
rect 217838 306856 219450 306864
rect 217777 306854 219450 306856
rect 376845 306856 376850 306912
rect 376906 306864 380052 306912
rect 376906 306856 379530 306864
rect 376845 306854 379530 306856
rect 57145 306851 57211 306854
rect 217777 306851 217843 306854
rect 376845 306851 376911 306854
rect -960 306234 480 306324
rect -960 306174 674 306234
rect -960 306098 480 306174
rect 614 306098 674 306174
rect -960 306084 674 306098
rect 246 306038 674 306084
rect 246 305554 306 306038
rect 57881 305962 57947 305965
rect 217041 305962 217107 305965
rect 219390 305962 220064 305972
rect 57881 305960 60062 305962
rect 57881 305904 57886 305960
rect 57942 305904 60062 305960
rect 57881 305902 60062 305904
rect 217041 305960 220064 305962
rect 217041 305904 217046 305960
rect 217102 305912 220064 305960
rect 377489 305962 377555 305965
rect 379470 305962 380052 305972
rect 377489 305960 380052 305962
rect 217102 305904 219450 305912
rect 217041 305902 219450 305904
rect 377489 305904 377494 305960
rect 377550 305912 380052 305960
rect 377550 305904 379530 305912
rect 377489 305902 379530 305904
rect 57881 305899 57947 305902
rect 217041 305899 217107 305902
rect 377489 305899 377555 305902
rect 246 305494 6930 305554
rect 6870 305010 6930 305494
rect 54334 305010 54340 305012
rect 6870 304950 54340 305010
rect 54334 304948 54340 304950
rect 54404 304948 54410 305012
rect 56869 305010 56935 305013
rect 57881 305010 57947 305013
rect 56869 305008 57947 305010
rect 56869 304952 56874 305008
rect 56930 304952 57886 305008
rect 57942 304952 57947 305008
rect 56869 304950 57947 304952
rect 56869 304947 56935 304950
rect 57881 304947 57947 304950
rect 376937 305010 377003 305013
rect 377489 305010 377555 305013
rect 376937 305008 377555 305010
rect 376937 304952 376942 305008
rect 376998 304952 377494 305008
rect 377550 304952 377555 305008
rect 376937 304950 377555 304952
rect 376937 304947 377003 304950
rect 377489 304947 377555 304950
rect 216765 303786 216831 303789
rect 217685 303786 217751 303789
rect 219390 303786 220064 303796
rect 216765 303784 220064 303786
rect 57329 303650 57395 303653
rect 57697 303650 57763 303653
rect 60002 303650 60062 303766
rect 216765 303728 216770 303784
rect 216826 303728 217690 303784
rect 217746 303736 220064 303784
rect 377213 303786 377279 303789
rect 379470 303786 380052 303796
rect 377213 303784 380052 303786
rect 217746 303728 219450 303736
rect 216765 303726 219450 303728
rect 377213 303728 377218 303784
rect 377274 303736 380052 303784
rect 377274 303728 379530 303736
rect 377213 303726 379530 303728
rect 216765 303723 216831 303726
rect 217685 303723 217751 303726
rect 377213 303723 377279 303726
rect 57329 303648 60062 303650
rect 57329 303592 57334 303648
rect 57390 303592 57702 303648
rect 57758 303592 60062 303648
rect 57329 303590 60062 303592
rect 57329 303587 57395 303590
rect 57697 303587 57763 303590
rect 217225 302834 217291 302837
rect 219390 302834 220064 302844
rect 217225 302832 220064 302834
rect 57513 302290 57579 302293
rect 60002 302290 60062 302814
rect 217225 302776 217230 302832
rect 217286 302784 220064 302832
rect 376753 302834 376819 302837
rect 377581 302834 377647 302837
rect 379470 302834 380052 302844
rect 376753 302832 380052 302834
rect 217286 302776 219450 302784
rect 217225 302774 219450 302776
rect 376753 302776 376758 302832
rect 376814 302776 377586 302832
rect 377642 302784 380052 302832
rect 377642 302776 379530 302784
rect 376753 302774 379530 302776
rect 217225 302771 217291 302774
rect 376753 302771 376819 302774
rect 377581 302771 377647 302774
rect 57513 302288 60062 302290
rect 57513 302232 57518 302288
rect 57574 302232 60062 302288
rect 57513 302230 60062 302232
rect 57513 302227 57579 302230
rect 57605 301338 57671 301341
rect 57605 301336 60062 301338
rect 57605 301280 57610 301336
rect 57666 301280 60062 301336
rect 57605 301278 60062 301280
rect 57605 301275 57671 301278
rect 60002 301046 60062 301278
rect 217501 301066 217567 301069
rect 219390 301066 220064 301076
rect 217501 301064 220064 301066
rect 217501 301008 217506 301064
rect 217562 301016 220064 301064
rect 376753 301066 376819 301069
rect 377673 301066 377739 301069
rect 379470 301066 380052 301076
rect 376753 301064 380052 301066
rect 217562 301008 219450 301016
rect 217501 301006 219450 301008
rect 376753 301008 376758 301064
rect 376814 301008 377678 301064
rect 377734 301016 380052 301064
rect 377734 301008 379530 301016
rect 376753 301006 379530 301008
rect 217501 301003 217567 301006
rect 376753 301003 376819 301006
rect 377673 301003 377739 301006
rect 216949 299978 217015 299981
rect 217409 299978 217475 299981
rect 219390 299978 220064 299988
rect 216949 299976 220064 299978
rect 57421 299570 57487 299573
rect 60002 299570 60062 299958
rect 216949 299920 216954 299976
rect 217010 299920 217414 299976
rect 217470 299928 220064 299976
rect 377305 299978 377371 299981
rect 379470 299978 380052 299988
rect 377305 299976 380052 299978
rect 217470 299920 219450 299928
rect 216949 299918 219450 299920
rect 377305 299920 377310 299976
rect 377366 299928 380052 299976
rect 377366 299920 379530 299928
rect 377305 299918 379530 299920
rect 216949 299915 217015 299918
rect 217409 299915 217475 299918
rect 377305 299915 377371 299918
rect 57421 299568 60062 299570
rect 57421 299512 57426 299568
rect 57482 299512 60062 299568
rect 57421 299510 60062 299512
rect 57421 299507 57487 299510
rect 216857 299434 216923 299437
rect 217593 299434 217659 299437
rect 216857 299432 217659 299434
rect 216857 299376 216862 299432
rect 216918 299376 217598 299432
rect 217654 299376 217659 299432
rect 216857 299374 217659 299376
rect 216857 299371 216923 299374
rect 217593 299371 217659 299374
rect 583520 298604 584960 298844
rect 57421 298210 57487 298213
rect 217593 298210 217659 298213
rect 219390 298210 220064 298220
rect 57421 298208 60062 298210
rect 57421 298152 57426 298208
rect 57482 298152 60062 298208
rect 57421 298150 60062 298152
rect 217593 298208 220064 298210
rect 217593 298152 217598 298208
rect 217654 298160 220064 298208
rect 377765 298210 377831 298213
rect 379470 298210 380052 298220
rect 377765 298208 380052 298210
rect 217654 298152 219450 298160
rect 217593 298150 219450 298152
rect 377765 298152 377770 298208
rect 377826 298160 380052 298208
rect 377826 298152 379530 298160
rect 377765 298150 379530 298152
rect 57421 298147 57487 298150
rect 217593 298147 217659 298150
rect 377765 298147 377831 298150
rect -960 293028 480 293268
rect 198825 289778 198891 289781
rect 199653 289778 199719 289781
rect 359181 289778 359247 289781
rect 359549 289778 359615 289781
rect 196558 289776 199719 289778
rect 196558 289720 198830 289776
rect 198886 289720 199658 289776
rect 199714 289720 199719 289776
rect 196558 289718 199719 289720
rect 196558 289350 196618 289718
rect 198825 289715 198891 289718
rect 199653 289715 199719 289718
rect 356562 289776 359615 289778
rect 356562 289720 359186 289776
rect 359242 289720 359554 289776
rect 359610 289720 359615 289776
rect 356562 289718 359615 289720
rect 356562 289350 356622 289718
rect 359181 289715 359247 289718
rect 359549 289715 359615 289718
rect 519261 289370 519327 289373
rect 516558 289368 519327 289370
rect 516558 289312 519266 289368
rect 519322 289312 519327 289368
rect 516558 289310 519327 289312
rect 519261 289307 519327 289310
rect 358905 288418 358971 288421
rect 359273 288418 359339 288421
rect 358905 288416 359339 288418
rect 358905 288360 358910 288416
rect 358966 288360 359278 288416
rect 359334 288360 359339 288416
rect 358905 288358 359339 288360
rect 358905 288355 358971 288358
rect 359273 288355 359339 288358
rect 518985 288418 519051 288421
rect 519353 288418 519419 288421
rect 518985 288416 519419 288418
rect 518985 288360 518990 288416
rect 519046 288360 519358 288416
rect 519414 288360 519419 288416
rect 518985 288358 519419 288360
rect 518985 288355 519051 288358
rect 519353 288355 519419 288358
rect 199745 287738 199811 287741
rect 358905 287738 358971 287741
rect 196558 287736 199811 287738
rect 196558 287680 199750 287736
rect 199806 287680 199811 287736
rect 196558 287678 199811 287680
rect 356562 287736 358971 287738
rect 356562 287680 358910 287736
rect 358966 287680 358971 287736
rect 356562 287678 358971 287680
rect 199745 287675 199811 287678
rect 358905 287675 358971 287678
rect 516558 287194 516618 287718
rect 518985 287194 519051 287197
rect 516558 287192 519051 287194
rect 516558 287136 518990 287192
rect 519046 287136 519051 287192
rect 516558 287134 519051 287136
rect 518985 287131 519051 287134
rect 199469 286378 199535 286381
rect 358997 286378 359063 286381
rect 196558 286376 199535 286378
rect 196558 286320 199474 286376
rect 199530 286320 199535 286376
rect 196558 286318 199535 286320
rect 356562 286376 359063 286378
rect 356562 286320 359002 286376
rect 359058 286320 359063 286376
rect 356562 286318 359063 286320
rect 199469 286315 199535 286318
rect 358997 286315 359063 286318
rect 516558 285834 516618 286358
rect 519445 285834 519511 285837
rect 516558 285832 519511 285834
rect 516558 285776 519450 285832
rect 519506 285776 519511 285832
rect 516558 285774 519511 285776
rect 519445 285771 519511 285774
rect 583520 285276 584960 285516
rect 519077 285018 519143 285021
rect 519905 285018 519971 285021
rect 517102 285016 519971 285018
rect 517102 284960 519082 285016
rect 519138 284960 519910 285016
rect 519966 284960 519971 285016
rect 517102 284958 519971 284960
rect 517102 284892 517162 284958
rect 519077 284955 519143 284958
rect 519905 284955 519971 284958
rect 199009 284882 199075 284885
rect 359457 284882 359523 284885
rect 196558 284880 199075 284882
rect 196558 284824 199014 284880
rect 199070 284824 199075 284880
rect 196558 284822 199075 284824
rect 356562 284880 359523 284882
rect 356562 284824 359462 284880
rect 359518 284824 359523 284880
rect 516588 284832 517162 284892
rect 356562 284822 359523 284824
rect 199009 284819 199075 284822
rect 359457 284819 359523 284822
rect 519169 284202 519235 284205
rect 516558 284200 519235 284202
rect 516558 284144 519174 284200
rect 519230 284144 519235 284200
rect 516558 284142 519235 284144
rect 516558 283638 516618 284142
rect 519169 284139 519235 284142
rect 196558 283114 196618 283638
rect 198917 283114 198983 283117
rect 199561 283114 199627 283117
rect 196558 283112 199627 283114
rect 196558 283056 198922 283112
rect 198978 283056 199566 283112
rect 199622 283056 199627 283112
rect 196558 283054 199627 283056
rect 356562 283114 356622 283638
rect 359089 283114 359155 283117
rect 359365 283114 359431 283117
rect 356562 283112 359431 283114
rect 356562 283056 359094 283112
rect 359150 283056 359370 283112
rect 359426 283056 359431 283112
rect 356562 283054 359431 283056
rect 198917 283051 198983 283054
rect 199561 283051 199627 283054
rect 359089 283051 359155 283054
rect 359365 283051 359431 283054
rect -960 279972 480 280212
rect 58709 279986 58775 279989
rect 216673 279986 216739 279989
rect 219390 279986 220064 279996
rect 58709 279984 60062 279986
rect 58709 279928 58714 279984
rect 58770 279928 60062 279984
rect 58709 279926 60062 279928
rect 216673 279984 220064 279986
rect 216673 279928 216678 279984
rect 216734 279936 220064 279984
rect 377029 279986 377095 279989
rect 379470 279986 380052 279996
rect 377029 279984 380052 279986
rect 216734 279928 219450 279936
rect 216673 279926 219450 279928
rect 377029 279928 377034 279984
rect 377090 279936 380052 279984
rect 377090 279928 379530 279936
rect 377029 279926 379530 279928
rect 58709 279923 58775 279926
rect 216673 279923 216739 279926
rect 377029 279923 377095 279926
rect 57237 278762 57303 278765
rect 57881 278762 57947 278765
rect 57237 278760 60062 278762
rect 57237 278704 57242 278760
rect 57298 278704 57886 278760
rect 57942 278704 60062 278760
rect 57237 278702 60062 278704
rect 57237 278699 57303 278702
rect 57881 278699 57947 278702
rect 60002 278334 60062 278702
rect 216673 278354 216739 278357
rect 219390 278354 220064 278364
rect 216673 278352 220064 278354
rect 216673 278296 216678 278352
rect 216734 278304 220064 278352
rect 377397 278354 377463 278357
rect 379470 278354 380052 278364
rect 377397 278352 380052 278354
rect 216734 278296 219450 278304
rect 216673 278294 219450 278296
rect 377397 278296 377402 278352
rect 377458 278304 380052 278352
rect 377458 278296 379530 278304
rect 377397 278294 379530 278296
rect 216673 278291 216739 278294
rect 377397 278291 377463 278294
rect 58801 278082 58867 278085
rect 216857 278082 216923 278085
rect 219390 278082 220064 278092
rect 58801 278080 60062 278082
rect 58801 278024 58806 278080
rect 58862 278024 60062 278080
rect 58801 278022 60062 278024
rect 216857 278080 220064 278082
rect 216857 278024 216862 278080
rect 216918 278032 220064 278080
rect 377029 278082 377095 278085
rect 379470 278082 380052 278092
rect 377029 278080 380052 278082
rect 216918 278024 219450 278032
rect 216857 278022 219450 278024
rect 377029 278024 377034 278080
rect 377090 278032 380052 278080
rect 377090 278024 379530 278032
rect 377029 278022 379530 278024
rect 58801 278019 58867 278022
rect 216857 278019 216923 278022
rect 377029 278019 377095 278022
rect 57094 276116 57100 276180
rect 57164 276178 57170 276180
rect 59813 276178 59879 276181
rect 57164 276176 59879 276178
rect 57164 276120 59818 276176
rect 59874 276120 59879 276176
rect 57164 276118 59879 276120
rect 57164 276116 57170 276118
rect 59813 276115 59879 276118
rect 57278 275980 57284 276044
rect 57348 276042 57354 276044
rect 58525 276042 58591 276045
rect 57348 276040 58591 276042
rect 57348 275984 58530 276040
rect 58586 275984 58591 276040
rect 57348 275982 58591 275984
rect 57348 275980 57354 275982
rect 58525 275979 58591 275982
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 580349 272171 580415 272174
rect 583520 272084 584960 272174
rect 211521 270602 211587 270605
rect 216622 270602 216628 270604
rect 211521 270600 216628 270602
rect 211521 270544 211526 270600
rect 211582 270544 216628 270600
rect 211521 270542 216628 270544
rect 211521 270539 211587 270542
rect 216622 270540 216628 270542
rect 216692 270602 216698 270604
rect 217358 270602 217364 270604
rect 216692 270542 217364 270602
rect 216692 270540 216698 270542
rect 217358 270540 217364 270542
rect 217428 270540 217434 270604
rect 211613 270466 211679 270469
rect 211838 270466 211844 270468
rect 211613 270464 211844 270466
rect 211613 270408 211618 270464
rect 211674 270408 211844 270464
rect 211613 270406 211844 270408
rect 211613 270403 211679 270406
rect 211838 270404 211844 270406
rect 211908 270404 211914 270468
rect 218329 270466 218395 270469
rect 218830 270466 218836 270468
rect 218329 270464 218836 270466
rect 218329 270408 218334 270464
rect 218390 270408 218836 270464
rect 218329 270406 218836 270408
rect 218329 270403 218395 270406
rect 218830 270404 218836 270406
rect 218900 270404 218906 270468
rect 378174 270404 378180 270468
rect 378244 270466 378250 270468
rect 378501 270466 378567 270469
rect 378244 270464 378567 270466
rect 378244 270408 378506 270464
rect 378562 270408 378567 270464
rect 378244 270406 378567 270408
rect 378244 270404 378250 270406
rect 378501 270403 378567 270406
rect 377990 270268 377996 270332
rect 378060 270330 378066 270332
rect 379237 270330 379303 270333
rect 378060 270328 379303 270330
rect 378060 270272 379242 270328
rect 379298 270272 379303 270328
rect 378060 270270 379303 270272
rect 378060 270268 378066 270270
rect 379237 270267 379303 270270
rect 107561 269924 107627 269925
rect 110965 269924 111031 269925
rect 250713 269924 250779 269925
rect 107561 269920 107606 269924
rect 107670 269922 107676 269924
rect 107561 269864 107566 269920
rect 107561 269860 107606 269864
rect 107670 269862 107718 269922
rect 110965 269920 111006 269924
rect 111070 269922 111076 269924
rect 110965 269864 110970 269920
rect 107670 269860 107676 269862
rect 110965 269860 111006 269864
rect 111070 269862 111122 269922
rect 250713 269920 250742 269924
rect 250806 269922 250812 269924
rect 263501 269922 263567 269925
rect 266376 269922 266382 269924
rect 250713 269864 250718 269920
rect 111070 269860 111076 269862
rect 250713 269860 250742 269864
rect 250806 269862 250870 269922
rect 263501 269920 266382 269922
rect 263501 269864 263506 269920
rect 263562 269864 266382 269920
rect 263501 269862 266382 269864
rect 250806 269860 250812 269862
rect 107561 269859 107627 269860
rect 110965 269859 111031 269860
rect 250713 269859 250779 269860
rect 263501 269859 263567 269862
rect 266376 269860 266382 269862
rect 266446 269860 266452 269924
rect 108297 269788 108363 269789
rect 108280 269786 108286 269788
rect 108206 269726 108286 269786
rect 108350 269784 108363 269788
rect 108358 269728 108363 269784
rect 108280 269724 108286 269726
rect 108350 269724 108363 269728
rect 108297 269723 108363 269724
rect 133413 269788 133479 269789
rect 135897 269788 135963 269789
rect 138473 269788 138539 269789
rect 275737 269788 275803 269789
rect 280889 269788 280955 269789
rect 315849 269788 315915 269789
rect 418429 269788 418495 269789
rect 425237 269788 425303 269789
rect 133413 269784 133446 269788
rect 133510 269786 133516 269788
rect 135888 269786 135894 269788
rect 133413 269728 133418 269784
rect 133413 269724 133446 269728
rect 133510 269726 133570 269786
rect 135806 269726 135894 269786
rect 133510 269724 133516 269726
rect 135888 269724 135894 269726
rect 135958 269724 135964 269788
rect 138472 269724 138478 269788
rect 138542 269786 138548 269788
rect 138542 269726 138630 269786
rect 138542 269724 138548 269726
rect 216622 269724 216628 269788
rect 216692 269786 216698 269788
rect 274400 269786 274406 269788
rect 216692 269726 274406 269786
rect 216692 269724 216698 269726
rect 274400 269724 274406 269726
rect 274470 269724 274476 269788
rect 275737 269784 275766 269788
rect 275830 269786 275836 269788
rect 275737 269728 275742 269784
rect 275737 269724 275766 269728
rect 275830 269726 275894 269786
rect 280889 269784 280934 269788
rect 280998 269786 281004 269788
rect 280889 269728 280894 269784
rect 275830 269724 275836 269726
rect 280889 269724 280934 269728
rect 280998 269726 281046 269786
rect 315849 269784 315886 269788
rect 315950 269786 315956 269788
rect 315849 269728 315854 269784
rect 280998 269724 281004 269726
rect 315849 269724 315886 269728
rect 315950 269726 316006 269786
rect 418429 269784 418494 269788
rect 418429 269728 418434 269784
rect 418490 269728 418494 269784
rect 315950 269724 315956 269726
rect 418429 269724 418494 269728
rect 418558 269786 418564 269788
rect 418558 269726 418586 269786
rect 425237 269784 425294 269788
rect 425358 269786 425364 269788
rect 425237 269728 425242 269784
rect 418558 269724 418564 269726
rect 425237 269724 425294 269728
rect 425358 269726 425394 269786
rect 425358 269724 425364 269726
rect 133413 269723 133479 269724
rect 135897 269723 135963 269724
rect 138473 269723 138539 269724
rect 275737 269723 275803 269724
rect 280889 269723 280955 269724
rect 315849 269723 315915 269724
rect 418429 269723 418495 269724
rect 425237 269723 425303 269724
rect 83089 269652 83155 269653
rect 93577 269652 93643 269653
rect 94497 269652 94563 269653
rect 108665 269652 108731 269653
rect 140865 269652 140931 269653
rect 143533 269652 143599 269653
rect 83089 269648 83126 269652
rect 83190 269650 83196 269652
rect 83089 269592 83094 269648
rect 83089 269588 83126 269592
rect 83190 269590 83246 269650
rect 93577 269648 93598 269652
rect 93662 269650 93668 269652
rect 93577 269592 93582 269648
rect 83190 269588 83196 269590
rect 93577 269588 93598 269592
rect 93662 269590 93734 269650
rect 94497 269648 94550 269652
rect 94614 269650 94620 269652
rect 94497 269592 94502 269648
rect 93662 269588 93668 269590
rect 94497 269588 94550 269592
rect 94614 269590 94654 269650
rect 108665 269648 108694 269652
rect 108758 269650 108764 269652
rect 108665 269592 108670 269648
rect 94614 269588 94620 269590
rect 108665 269588 108694 269592
rect 108758 269590 108822 269650
rect 140865 269648 140926 269652
rect 140865 269592 140870 269648
rect 108758 269588 108764 269590
rect 140865 269588 140926 269592
rect 140990 269650 140996 269652
rect 143504 269650 143510 269652
rect 140990 269590 141022 269650
rect 143442 269590 143510 269650
rect 143574 269648 143599 269652
rect 143594 269592 143599 269648
rect 140990 269588 140996 269590
rect 143504 269588 143510 269590
rect 143574 269588 143599 269592
rect 83089 269587 83155 269588
rect 93577 269587 93643 269588
rect 94497 269587 94563 269588
rect 108665 269587 108731 269588
rect 140865 269587 140931 269588
rect 143533 269587 143599 269588
rect 145925 269652 145991 269653
rect 279141 269652 279207 269653
rect 283465 269652 283531 269653
rect 285949 269652 286015 269653
rect 288249 269652 288315 269653
rect 293401 269652 293467 269653
rect 308489 269652 308555 269653
rect 318425 269652 318491 269653
rect 423489 269652 423555 269653
rect 426433 269652 426499 269653
rect 433609 269652 433675 269653
rect 145925 269648 145958 269652
rect 146022 269650 146028 269652
rect 145925 269592 145930 269648
rect 145925 269588 145958 269592
rect 146022 269590 146082 269650
rect 279141 269648 279166 269652
rect 279230 269650 279236 269652
rect 279141 269592 279146 269648
rect 146022 269588 146028 269590
rect 279141 269588 279166 269592
rect 279230 269590 279298 269650
rect 283465 269648 283518 269652
rect 283582 269650 283588 269652
rect 283465 269592 283470 269648
rect 279230 269588 279236 269590
rect 283465 269588 283518 269592
rect 283582 269590 283622 269650
rect 285949 269648 285966 269652
rect 286030 269650 286036 269652
rect 285949 269592 285954 269648
rect 283582 269588 283588 269590
rect 285949 269588 285966 269592
rect 286030 269590 286106 269650
rect 288249 269648 288278 269652
rect 288342 269650 288348 269652
rect 288249 269592 288254 269648
rect 286030 269588 286036 269590
rect 288249 269588 288278 269592
rect 288342 269590 288406 269650
rect 293401 269648 293446 269652
rect 293510 269650 293516 269652
rect 293401 269592 293406 269648
rect 288342 269588 288348 269590
rect 293401 269588 293446 269592
rect 293510 269590 293558 269650
rect 308489 269648 308542 269652
rect 308606 269650 308612 269652
rect 308489 269592 308494 269648
rect 293510 269588 293516 269590
rect 308489 269588 308542 269592
rect 308606 269590 308646 269650
rect 318425 269648 318470 269652
rect 318534 269650 318540 269652
rect 318425 269592 318430 269648
rect 308606 269588 308612 269590
rect 318425 269588 318470 269592
rect 318534 269590 318582 269650
rect 423489 269648 423526 269652
rect 423590 269650 423596 269652
rect 426382 269650 426388 269652
rect 423489 269592 423494 269648
rect 318534 269588 318540 269590
rect 423489 269588 423526 269592
rect 423590 269590 423646 269650
rect 426342 269590 426388 269650
rect 426452 269648 426499 269652
rect 433584 269650 433590 269652
rect 426494 269592 426499 269648
rect 423590 269588 423596 269590
rect 426382 269588 426388 269590
rect 426452 269588 426499 269592
rect 433518 269590 433590 269650
rect 433654 269648 433675 269652
rect 433670 269592 433675 269648
rect 433584 269588 433590 269590
rect 433654 269588 433675 269592
rect 145925 269587 145991 269588
rect 279141 269587 279207 269588
rect 283465 269587 283531 269588
rect 285949 269587 286015 269588
rect 288249 269587 288315 269588
rect 293401 269587 293467 269588
rect 308489 269587 308555 269588
rect 318425 269587 318491 269588
rect 423489 269587 423555 269588
rect 426433 269587 426499 269588
rect 433609 269587 433675 269588
rect 453389 269652 453455 269653
rect 468477 269652 468543 269653
rect 480897 269652 480963 269653
rect 453389 269648 453446 269652
rect 453510 269650 453516 269652
rect 453389 269592 453394 269648
rect 453389 269588 453446 269592
rect 453510 269590 453546 269650
rect 468477 269648 468542 269652
rect 468477 269592 468482 269648
rect 468538 269592 468542 269648
rect 453510 269588 453516 269590
rect 468477 269588 468542 269592
rect 468606 269650 468612 269652
rect 468606 269590 468634 269650
rect 480897 269648 480918 269652
rect 480982 269650 480988 269652
rect 480897 269592 480902 269648
rect 468606 269588 468612 269590
rect 480897 269588 480918 269592
rect 480982 269590 481054 269650
rect 480982 269588 480988 269590
rect 453389 269587 453455 269588
rect 468477 269587 468543 269588
rect 480897 269587 480963 269588
rect 373901 269378 373967 269381
rect 376886 269378 376892 269380
rect 373901 269376 376892 269378
rect 373901 269320 373906 269376
rect 373962 269320 376892 269376
rect 373901 269318 376892 269320
rect 373901 269315 373967 269318
rect 376886 269316 376892 269318
rect 376956 269378 376962 269380
rect 377622 269378 377628 269380
rect 376956 269318 377628 269378
rect 376956 269316 376962 269318
rect 377622 269316 377628 269318
rect 377692 269316 377698 269380
rect 359406 269180 359412 269244
rect 359476 269242 359482 269244
rect 470910 269242 470916 269244
rect 359476 269182 470916 269242
rect 359476 269180 359482 269182
rect 470910 269180 470916 269182
rect 470980 269180 470986 269244
rect 57278 269044 57284 269108
rect 57348 269106 57354 269108
rect 60917 269106 60983 269109
rect 57348 269104 60983 269106
rect 57348 269048 60922 269104
rect 60978 269048 60983 269104
rect 57348 269046 60983 269048
rect 57348 269044 57354 269046
rect 60917 269043 60983 269046
rect 76005 269108 76071 269109
rect 77109 269108 77175 269109
rect 90725 269108 90791 269109
rect 95877 269108 95943 269109
rect 96061 269108 96127 269109
rect 98453 269108 98519 269109
rect 99373 269108 99439 269109
rect 76005 269104 76052 269108
rect 76116 269106 76122 269108
rect 76005 269048 76010 269104
rect 76005 269044 76052 269048
rect 76116 269046 76162 269106
rect 77109 269104 77156 269108
rect 77220 269106 77226 269108
rect 77109 269048 77114 269104
rect 76116 269044 76122 269046
rect 77109 269044 77156 269048
rect 77220 269046 77266 269106
rect 90725 269104 90772 269108
rect 90836 269106 90842 269108
rect 95877 269106 95924 269108
rect 90725 269048 90730 269104
rect 77220 269044 77226 269046
rect 90725 269044 90772 269048
rect 90836 269046 90882 269106
rect 95832 269104 95924 269106
rect 95832 269048 95882 269104
rect 95832 269046 95924 269048
rect 90836 269044 90842 269046
rect 95877 269044 95924 269046
rect 95988 269044 95994 269108
rect 96061 269104 96108 269108
rect 96172 269106 96178 269108
rect 96061 269048 96066 269104
rect 96061 269044 96108 269048
rect 96172 269046 96218 269106
rect 98453 269104 98500 269108
rect 98564 269106 98570 269108
rect 98453 269048 98458 269104
rect 96172 269044 96178 269046
rect 98453 269044 98500 269048
rect 98564 269046 98610 269106
rect 99373 269104 99420 269108
rect 99484 269106 99490 269108
rect 99373 269048 99378 269104
rect 98564 269044 98570 269046
rect 99373 269044 99420 269048
rect 99484 269046 99530 269106
rect 99484 269044 99490 269046
rect 212574 269044 212580 269108
rect 212644 269106 212650 269108
rect 213729 269106 213795 269109
rect 298461 269108 298527 269109
rect 300853 269108 300919 269109
rect 212644 269104 213795 269106
rect 212644 269048 213734 269104
rect 213790 269048 213795 269104
rect 212644 269046 213795 269048
rect 212644 269044 212650 269046
rect 76005 269043 76071 269044
rect 77109 269043 77175 269044
rect 90725 269043 90791 269044
rect 95877 269043 95943 269044
rect 96061 269043 96127 269044
rect 98453 269043 98519 269044
rect 99373 269043 99439 269044
rect 213729 269043 213795 269046
rect 217174 269044 217180 269108
rect 217244 269106 217250 269108
rect 217244 269046 296730 269106
rect 217244 269044 217250 269046
rect 60733 268970 60799 268973
rect 290917 268972 290983 268973
rect 295885 268972 295951 268973
rect 115790 268970 115796 268972
rect 60733 268968 115796 268970
rect 60733 268912 60738 268968
rect 60794 268912 115796 268968
rect 60733 268910 115796 268912
rect 60733 268907 60799 268910
rect 115790 268908 115796 268910
rect 115860 268908 115866 268972
rect 199326 268908 199332 268972
rect 199396 268970 199402 268972
rect 278446 268970 278452 268972
rect 199396 268910 278452 268970
rect 199396 268908 199402 268910
rect 278446 268908 278452 268910
rect 278516 268908 278522 268972
rect 290917 268968 290964 268972
rect 291028 268970 291034 268972
rect 290917 268912 290922 268968
rect 290917 268908 290964 268912
rect 291028 268910 291074 268970
rect 295885 268968 295932 268972
rect 295996 268970 296002 268972
rect 296670 268970 296730 269046
rect 298461 269104 298508 269108
rect 298572 269106 298578 269108
rect 298461 269048 298466 269104
rect 298461 269044 298508 269048
rect 298572 269046 298618 269106
rect 300853 269104 300900 269108
rect 300964 269106 300970 269108
rect 356789 269106 356855 269109
rect 485998 269106 486004 269108
rect 300853 269048 300858 269104
rect 298572 269044 298578 269046
rect 300853 269044 300900 269048
rect 300964 269046 301010 269106
rect 356789 269104 486004 269106
rect 356789 269048 356794 269104
rect 356850 269048 486004 269104
rect 356789 269046 486004 269048
rect 300964 269044 300970 269046
rect 298461 269043 298527 269044
rect 300853 269043 300919 269044
rect 356789 269043 356855 269046
rect 485998 269044 486004 269046
rect 486068 269044 486074 269108
rect 430941 268972 431007 268973
rect 433333 268972 433399 268973
rect 475837 268972 475903 268973
rect 478413 268972 478479 268973
rect 483381 268972 483447 268973
rect 305862 268970 305868 268972
rect 295885 268912 295890 268968
rect 291028 268908 291034 268910
rect 295885 268908 295932 268912
rect 295996 268910 296042 268970
rect 296670 268910 305868 268970
rect 295996 268908 296002 268910
rect 305862 268908 305868 268910
rect 305932 268908 305938 268972
rect 377254 268908 377260 268972
rect 377324 268970 377330 268972
rect 426014 268970 426020 268972
rect 377324 268910 426020 268970
rect 377324 268908 377330 268910
rect 426014 268908 426020 268910
rect 426084 268908 426090 268972
rect 430941 268968 430988 268972
rect 431052 268970 431058 268972
rect 430941 268912 430946 268968
rect 430941 268908 430988 268912
rect 431052 268910 431098 268970
rect 433333 268968 433380 268972
rect 433444 268970 433450 268972
rect 433333 268912 433338 268968
rect 431052 268908 431058 268910
rect 433333 268908 433380 268912
rect 433444 268910 433490 268970
rect 475837 268968 475884 268972
rect 475948 268970 475954 268972
rect 475837 268912 475842 268968
rect 433444 268908 433450 268910
rect 475837 268908 475884 268912
rect 475948 268910 475994 268970
rect 478413 268968 478460 268972
rect 478524 268970 478530 268972
rect 478413 268912 478418 268968
rect 475948 268908 475954 268910
rect 478413 268908 478460 268912
rect 478524 268910 478570 268970
rect 483381 268968 483428 268972
rect 483492 268970 483498 268972
rect 483381 268912 483386 268968
rect 478524 268908 478530 268910
rect 483381 268908 483428 268912
rect 483492 268910 483538 268970
rect 483492 268908 483498 268910
rect 290917 268907 290983 268908
rect 295885 268907 295951 268908
rect 430941 268907 431007 268908
rect 433333 268907 433399 268908
rect 475837 268907 475903 268908
rect 478413 268907 478479 268908
rect 483381 268907 483447 268908
rect 59813 268834 59879 268837
rect 61009 268834 61075 268837
rect 243077 268836 243143 268837
rect 117998 268834 118004 268836
rect 59813 268832 118004 268834
rect 59813 268776 59818 268832
rect 59874 268776 61014 268832
rect 61070 268776 118004 268832
rect 59813 268774 118004 268776
rect 59813 268771 59879 268774
rect 61009 268771 61075 268774
rect 117998 268772 118004 268774
rect 118068 268772 118074 268836
rect 243077 268832 243124 268836
rect 243188 268834 243194 268836
rect 243077 268776 243082 268832
rect 243077 268772 243124 268776
rect 243188 268774 243234 268834
rect 243188 268772 243194 268774
rect 257838 268772 257844 268836
rect 257908 268834 257914 268836
rect 258073 268834 258139 268837
rect 257908 268832 258139 268834
rect 257908 268776 258078 268832
rect 258134 268776 258139 268832
rect 257908 268774 258139 268776
rect 257908 268772 257914 268774
rect 243077 268771 243143 268772
rect 258073 268771 258139 268774
rect 261661 268836 261727 268837
rect 415853 268836 415919 268837
rect 421005 268836 421071 268837
rect 261661 268832 261708 268836
rect 261772 268834 261778 268836
rect 261661 268776 261666 268832
rect 261661 268772 261708 268776
rect 261772 268774 261818 268834
rect 261772 268772 261778 268774
rect 377622 268772 377628 268836
rect 377692 268834 377698 268836
rect 377692 268774 412650 268834
rect 377692 268772 377698 268774
rect 261661 268771 261727 268772
rect 60917 268698 60983 268701
rect 119102 268698 119108 268700
rect 60917 268696 119108 268698
rect 60917 268640 60922 268696
rect 60978 268640 119108 268696
rect 60917 268638 119108 268640
rect 60917 268635 60983 268638
rect 119102 268636 119108 268638
rect 119172 268636 119178 268700
rect 412590 268698 412650 268774
rect 415853 268832 415900 268836
rect 415964 268834 415970 268836
rect 415853 268776 415858 268832
rect 415853 268772 415900 268776
rect 415964 268774 416010 268834
rect 421005 268832 421052 268836
rect 421116 268834 421122 268836
rect 421005 268776 421010 268832
rect 415964 268772 415970 268774
rect 421005 268772 421052 268776
rect 421116 268774 421162 268834
rect 421116 268772 421122 268774
rect 415853 268771 415919 268772
rect 421005 268771 421071 268772
rect 423990 268698 423996 268700
rect 412590 268638 423996 268698
rect 423990 268636 423996 268638
rect 424060 268636 424066 268700
rect 47393 268562 47459 268565
rect 109718 268562 109724 268564
rect 47393 268560 109724 268562
rect 47393 268504 47398 268560
rect 47454 268504 109724 268560
rect 47393 268502 109724 268504
rect 47393 268499 47459 268502
rect 109718 268500 109724 268502
rect 109788 268500 109794 268564
rect 47301 268426 47367 268429
rect 111190 268426 111196 268428
rect 47301 268424 111196 268426
rect 47301 268368 47306 268424
rect 47362 268368 111196 268424
rect 47301 268366 111196 268368
rect 47301 268363 47367 268366
rect 111190 268364 111196 268366
rect 111260 268364 111266 268428
rect 85389 268156 85455 268157
rect 92381 268156 92447 268157
rect 85389 268152 85436 268156
rect 85500 268154 85506 268156
rect 85389 268096 85394 268152
rect 85389 268092 85436 268096
rect 85500 268094 85546 268154
rect 92381 268152 92428 268156
rect 92492 268154 92498 268156
rect 92381 268096 92386 268152
rect 85500 268092 85506 268094
rect 92381 268092 92428 268096
rect 92492 268094 92538 268154
rect 92492 268092 92498 268094
rect 103278 268092 103284 268156
rect 103348 268154 103354 268156
rect 103513 268154 103579 268157
rect 128353 268156 128419 268157
rect 153561 268156 153627 268157
rect 103348 268152 103579 268154
rect 103348 268096 103518 268152
rect 103574 268096 103579 268152
rect 103348 268094 103579 268096
rect 103348 268092 103354 268094
rect 85389 268091 85455 268092
rect 92381 268091 92447 268092
rect 103513 268091 103579 268094
rect 113582 268092 113588 268156
rect 113652 268092 113658 268156
rect 128302 268154 128308 268156
rect 128262 268094 128308 268154
rect 128372 268152 128419 268156
rect 153510 268154 153516 268156
rect 128414 268096 128419 268152
rect 128302 268092 128308 268094
rect 128372 268092 128419 268096
rect 153470 268094 153516 268154
rect 153580 268152 153627 268156
rect 153622 268096 153627 268152
rect 153510 268092 153516 268094
rect 153580 268092 153627 268096
rect 113265 268020 113331 268021
rect 113214 268018 113220 268020
rect 113174 267958 113220 268018
rect 113284 268016 113331 268020
rect 113326 267960 113331 268016
rect 113214 267956 113220 267958
rect 113284 267956 113331 267960
rect 113265 267955 113331 267956
rect 113590 267882 113650 268092
rect 128353 268091 128419 268092
rect 153561 268091 153627 268092
rect 265157 268156 265223 268157
rect 272149 268156 272215 268157
rect 398189 268156 398255 268157
rect 401685 268156 401751 268157
rect 416037 268156 416103 268157
rect 434253 268156 434319 268157
rect 455781 268156 455847 268157
rect 265157 268152 265204 268156
rect 265268 268154 265274 268156
rect 265157 268096 265162 268152
rect 265157 268092 265204 268096
rect 265268 268094 265314 268154
rect 272149 268152 272196 268156
rect 272260 268154 272266 268156
rect 272149 268096 272154 268152
rect 265268 268092 265274 268094
rect 272149 268092 272196 268096
rect 272260 268094 272306 268154
rect 398189 268152 398236 268156
rect 398300 268154 398306 268156
rect 398189 268096 398194 268152
rect 272260 268092 272266 268094
rect 398189 268092 398236 268096
rect 398300 268094 398346 268154
rect 401685 268152 401732 268156
rect 401796 268154 401802 268156
rect 401685 268096 401690 268152
rect 398300 268092 398306 268094
rect 401685 268092 401732 268096
rect 401796 268094 401842 268154
rect 416037 268152 416084 268156
rect 416148 268154 416154 268156
rect 416037 268096 416042 268152
rect 401796 268092 401802 268094
rect 416037 268092 416084 268096
rect 416148 268094 416194 268154
rect 434253 268152 434300 268156
rect 434364 268154 434370 268156
rect 434253 268096 434258 268152
rect 416148 268092 416154 268094
rect 434253 268092 434300 268096
rect 434364 268094 434410 268154
rect 455781 268152 455828 268156
rect 455892 268154 455898 268156
rect 455781 268096 455786 268152
rect 434364 268092 434370 268094
rect 455781 268092 455828 268096
rect 455892 268094 455938 268154
rect 455892 268092 455898 268094
rect 265157 268091 265223 268092
rect 272149 268091 272215 268092
rect 398189 268091 398255 268092
rect 401685 268091 401751 268092
rect 416037 268091 416103 268092
rect 434253 268091 434319 268092
rect 455781 268091 455847 268092
rect 113130 267822 113650 267882
rect 113130 267749 113190 267822
rect 83958 267684 83964 267748
rect 84028 267746 84034 267748
rect 84193 267746 84259 267749
rect 84028 267744 84259 267746
rect 84028 267688 84198 267744
rect 84254 267688 84259 267744
rect 84028 267686 84259 267688
rect 84028 267684 84034 267686
rect 84193 267683 84259 267686
rect 86953 267746 87019 267749
rect 102685 267748 102751 267749
rect 105261 267748 105327 267749
rect 106365 267748 106431 267749
rect 87454 267746 87460 267748
rect 86953 267744 87460 267746
rect 86953 267688 86958 267744
rect 87014 267688 87460 267744
rect 86953 267686 87460 267688
rect 86953 267683 87019 267686
rect 87454 267684 87460 267686
rect 87524 267684 87530 267748
rect 102685 267746 102732 267748
rect 102640 267744 102732 267746
rect 102640 267688 102690 267744
rect 102640 267686 102732 267688
rect 102685 267684 102732 267686
rect 102796 267684 102802 267748
rect 105261 267746 105308 267748
rect 105216 267744 105308 267746
rect 105216 267688 105266 267744
rect 105216 267686 105308 267688
rect 105261 267684 105308 267686
rect 105372 267684 105378 267748
rect 106365 267746 106412 267748
rect 106320 267744 106412 267746
rect 106320 267688 106370 267744
rect 106320 267686 106412 267688
rect 106365 267684 106412 267686
rect 106476 267684 106482 267748
rect 113130 267744 113239 267749
rect 117129 267748 117195 267749
rect 117078 267746 117084 267748
rect 113130 267688 113178 267744
rect 113234 267688 113239 267744
rect 113130 267686 113239 267688
rect 117038 267686 117084 267746
rect 117148 267744 117195 267748
rect 117190 267688 117195 267744
rect 102685 267683 102751 267684
rect 105261 267683 105327 267684
rect 106365 267683 106431 267684
rect 113173 267683 113239 267686
rect 117078 267684 117084 267686
rect 117148 267684 117195 267688
rect 117129 267683 117195 267684
rect 122833 267746 122899 267749
rect 123518 267746 123524 267748
rect 122833 267744 123524 267746
rect 122833 267688 122838 267744
rect 122894 267688 123524 267744
rect 122833 267686 123524 267688
rect 122833 267683 122899 267686
rect 123518 267684 123524 267686
rect 123588 267684 123594 267748
rect 129733 267746 129799 267749
rect 155953 267748 156019 267749
rect 158529 267748 158595 267749
rect 163497 267748 163563 267749
rect 130878 267746 130884 267748
rect 129733 267744 130884 267746
rect 129733 267688 129738 267744
rect 129794 267688 130884 267744
rect 129733 267686 130884 267688
rect 129733 267683 129799 267686
rect 130878 267684 130884 267686
rect 130948 267684 130954 267748
rect 155902 267746 155908 267748
rect 155862 267686 155908 267746
rect 155972 267744 156019 267748
rect 158478 267746 158484 267748
rect 156014 267688 156019 267744
rect 155902 267684 155908 267686
rect 155972 267684 156019 267688
rect 158438 267686 158484 267746
rect 158548 267744 158595 267748
rect 163446 267746 163452 267748
rect 158590 267688 158595 267744
rect 158478 267684 158484 267686
rect 158548 267684 158595 267688
rect 163406 267686 163452 267746
rect 163516 267744 163563 267748
rect 255773 267748 255839 267749
rect 255773 267746 255820 267748
rect 163558 267688 163563 267744
rect 163446 267684 163452 267686
rect 163516 267684 163563 267688
rect 255728 267744 255820 267746
rect 255728 267688 255778 267744
rect 255728 267686 255820 267688
rect 155953 267683 156019 267684
rect 158529 267683 158595 267684
rect 163497 267683 163563 267684
rect 255773 267684 255820 267686
rect 255884 267684 255890 267748
rect 260833 267746 260899 267749
rect 260966 267746 260972 267748
rect 260833 267744 260972 267746
rect 260833 267688 260838 267744
rect 260894 267688 260972 267744
rect 260833 267686 260972 267688
rect 255773 267683 255839 267684
rect 260833 267683 260899 267686
rect 260966 267684 260972 267686
rect 261036 267684 261042 267748
rect 263593 267746 263659 267749
rect 263726 267746 263732 267748
rect 263593 267744 263732 267746
rect 263593 267688 263598 267744
rect 263654 267688 263732 267744
rect 263593 267686 263732 267688
rect 263593 267683 263659 267686
rect 263726 267684 263732 267686
rect 263796 267684 263802 267748
rect 265801 267746 265867 267749
rect 265934 267746 265940 267748
rect 265801 267744 265940 267746
rect 265801 267688 265806 267744
rect 265862 267688 265940 267744
rect 265801 267686 265940 267688
rect 265801 267683 265867 267686
rect 265934 267684 265940 267686
rect 266004 267684 266010 267748
rect 267089 267746 267155 267749
rect 267590 267746 267596 267748
rect 267089 267744 267596 267746
rect 267089 267688 267094 267744
rect 267150 267688 267596 267744
rect 267089 267686 267596 267688
rect 267089 267683 267155 267686
rect 267590 267684 267596 267686
rect 267660 267684 267666 267748
rect 268193 267746 268259 267749
rect 270861 267748 270927 267749
rect 268326 267746 268332 267748
rect 268193 267744 268332 267746
rect 268193 267688 268198 267744
rect 268254 267688 268332 267744
rect 268193 267686 268332 267688
rect 268193 267683 268259 267686
rect 268326 267684 268332 267686
rect 268396 267684 268402 267748
rect 270861 267744 270908 267748
rect 270972 267746 270978 267748
rect 273253 267746 273319 267749
rect 273478 267746 273484 267748
rect 270861 267688 270866 267744
rect 270861 267684 270908 267688
rect 270972 267686 271018 267746
rect 273253 267744 273484 267746
rect 273253 267688 273258 267744
rect 273314 267688 273484 267744
rect 273253 267686 273484 267688
rect 270972 267684 270978 267686
rect 270861 267683 270927 267684
rect 273253 267683 273319 267686
rect 273478 267684 273484 267686
rect 273548 267684 273554 267748
rect 276013 267746 276079 267749
rect 276238 267746 276244 267748
rect 276013 267744 276244 267746
rect 276013 267688 276018 267744
rect 276074 267688 276244 267744
rect 276013 267686 276244 267688
rect 276013 267683 276079 267686
rect 276238 267684 276244 267686
rect 276308 267684 276314 267748
rect 302233 267746 302299 267749
rect 402973 267748 403039 267749
rect 414381 267748 414447 267749
rect 303470 267746 303476 267748
rect 302233 267744 303476 267746
rect 302233 267688 302238 267744
rect 302294 267688 303476 267744
rect 302233 267686 303476 267688
rect 302233 267683 302299 267686
rect 303470 267684 303476 267686
rect 303540 267684 303546 267748
rect 402973 267744 403020 267748
rect 403084 267746 403090 267748
rect 414381 267746 414428 267748
rect 402973 267688 402978 267744
rect 402973 267684 403020 267688
rect 403084 267686 403130 267746
rect 414336 267744 414428 267746
rect 414336 267688 414386 267744
rect 414336 267686 414428 267688
rect 403084 267684 403090 267686
rect 414381 267684 414428 267686
rect 414492 267684 414498 267748
rect 432137 267746 432203 267749
rect 435725 267748 435791 267749
rect 435909 267748 435975 267749
rect 432270 267746 432276 267748
rect 432137 267744 432276 267746
rect 432137 267688 432142 267744
rect 432198 267688 432276 267744
rect 432137 267686 432276 267688
rect 402973 267683 403039 267684
rect 414381 267683 414447 267684
rect 432137 267683 432203 267686
rect 432270 267684 432276 267686
rect 432340 267684 432346 267748
rect 435725 267746 435772 267748
rect 435680 267744 435772 267746
rect 435680 267688 435730 267744
rect 435680 267686 435772 267688
rect 435725 267684 435772 267686
rect 435836 267684 435842 267748
rect 435909 267744 435956 267748
rect 436020 267746 436026 267748
rect 445753 267746 445819 267749
rect 445886 267746 445892 267748
rect 435909 267688 435914 267744
rect 435909 267684 435956 267688
rect 436020 267686 436066 267746
rect 445753 267744 445892 267746
rect 445753 267688 445758 267744
rect 445814 267688 445892 267744
rect 445753 267686 445892 267688
rect 436020 267684 436026 267686
rect 435725 267683 435791 267684
rect 435909 267683 435975 267684
rect 445753 267683 445819 267686
rect 445886 267684 445892 267686
rect 445956 267684 445962 267748
rect 447133 267746 447199 267749
rect 448278 267746 448284 267748
rect 447133 267744 448284 267746
rect 447133 267688 447138 267744
rect 447194 267688 448284 267744
rect 447133 267686 448284 267688
rect 447133 267683 447199 267686
rect 448278 267684 448284 267686
rect 448348 267684 448354 267748
rect 449893 267746 449959 267749
rect 451038 267746 451044 267748
rect 449893 267744 451044 267746
rect 449893 267688 449898 267744
rect 449954 267688 451044 267744
rect 449893 267686 451044 267688
rect 449893 267683 449959 267686
rect 451038 267684 451044 267686
rect 451108 267684 451114 267748
rect 458173 267746 458239 267749
rect 473353 267748 473419 267749
rect 458398 267746 458404 267748
rect 458173 267744 458404 267746
rect 458173 267688 458178 267744
rect 458234 267688 458404 267744
rect 458173 267686 458404 267688
rect 458173 267683 458239 267686
rect 458398 267684 458404 267686
rect 458468 267684 458474 267748
rect 473302 267746 473308 267748
rect 473262 267686 473308 267746
rect 473372 267744 473419 267748
rect 473414 267688 473419 267744
rect 473302 267684 473308 267686
rect 473372 267684 473419 267688
rect 473353 267683 473419 267684
rect 46473 267610 46539 267613
rect 79542 267610 79548 267612
rect 46473 267608 79548 267610
rect 46473 267552 46478 267608
rect 46534 267552 79548 267608
rect 46473 267550 79548 267552
rect 46473 267547 46539 267550
rect 79542 267548 79548 267550
rect 79612 267548 79618 267612
rect 125593 267610 125659 267613
rect 125910 267610 125916 267612
rect 125593 267608 125916 267610
rect 125593 267552 125598 267608
rect 125654 267552 125916 267608
rect 125593 267550 125916 267552
rect 125593 267547 125659 267550
rect 125910 267548 125916 267550
rect 125980 267548 125986 267612
rect 150934 267548 150940 267612
rect 151004 267610 151010 267612
rect 198958 267610 198964 267612
rect 151004 267550 198964 267610
rect 151004 267548 151010 267550
rect 198958 267548 198964 267550
rect 199028 267548 199034 267612
rect 209405 267610 209471 267613
rect 323342 267610 323348 267612
rect 209405 267608 323348 267610
rect 209405 267552 209410 267608
rect 209466 267552 323348 267608
rect 209405 267550 323348 267552
rect 209405 267547 209471 267550
rect 323342 267548 323348 267550
rect 323412 267548 323418 267612
rect 378961 267610 379027 267613
rect 465942 267610 465948 267612
rect 378961 267608 465948 267610
rect 378961 267552 378966 267608
rect 379022 267552 465948 267608
rect 378961 267550 465948 267552
rect 378961 267547 379027 267550
rect 465942 267548 465948 267550
rect 466012 267548 466018 267612
rect 49049 267474 49115 267477
rect 81934 267474 81940 267476
rect 49049 267472 81940 267474
rect 49049 267416 49054 267472
rect 49110 267416 81940 267472
rect 49049 267414 81940 267416
rect 49049 267411 49115 267414
rect 81934 267412 81940 267414
rect 82004 267412 82010 267476
rect 117313 267474 117379 267477
rect 118366 267474 118372 267476
rect 117313 267472 118372 267474
rect 117313 267416 117318 267472
rect 117374 267416 118372 267472
rect 117313 267414 118372 267416
rect 117313 267411 117379 267414
rect 118366 267412 118372 267414
rect 118436 267412 118442 267476
rect 120073 267474 120139 267477
rect 160921 267476 160987 267477
rect 120758 267474 120764 267476
rect 120073 267472 120764 267474
rect 120073 267416 120078 267472
rect 120134 267416 120764 267472
rect 120073 267414 120764 267416
rect 120073 267411 120139 267414
rect 120758 267412 120764 267414
rect 120828 267412 120834 267476
rect 160870 267474 160876 267476
rect 160830 267414 160876 267474
rect 160940 267472 160987 267476
rect 160982 267416 160987 267472
rect 160870 267412 160876 267414
rect 160940 267412 160987 267416
rect 166022 267412 166028 267476
rect 166092 267474 166098 267476
rect 166165 267474 166231 267477
rect 166092 267472 166231 267474
rect 166092 267416 166170 267472
rect 166226 267416 166231 267472
rect 166092 267414 166231 267416
rect 166092 267412 166098 267414
rect 160921 267411 160987 267412
rect 166165 267411 166231 267414
rect 183461 267476 183527 267477
rect 183461 267472 183508 267476
rect 183572 267474 183578 267476
rect 209221 267474 209287 267477
rect 343449 267476 343515 267477
rect 320950 267474 320956 267476
rect 183461 267416 183466 267472
rect 183461 267412 183508 267416
rect 183572 267414 183618 267474
rect 209221 267472 320956 267474
rect 209221 267416 209226 267472
rect 209282 267416 320956 267472
rect 209221 267414 320956 267416
rect 183572 267412 183578 267414
rect 183461 267411 183527 267412
rect 209221 267411 209287 267414
rect 320950 267412 320956 267414
rect 321020 267412 321026 267476
rect 343398 267474 343404 267476
rect 343358 267414 343404 267474
rect 343468 267472 343515 267476
rect 343510 267416 343515 267472
rect 343398 267412 343404 267414
rect 343468 267412 343515 267416
rect 343449 267411 343515 267412
rect 374177 267474 374243 267477
rect 503529 267476 503595 267477
rect 460974 267474 460980 267476
rect 374177 267472 460980 267474
rect 374177 267416 374182 267472
rect 374238 267416 460980 267472
rect 374177 267414 460980 267416
rect 374177 267411 374243 267414
rect 460974 267412 460980 267414
rect 461044 267412 461050 267476
rect 503478 267474 503484 267476
rect 503438 267414 503484 267474
rect 503548 267472 503595 267476
rect 503590 267416 503595 267472
rect 503478 267412 503484 267414
rect 503548 267412 503595 267416
rect 503529 267411 503595 267412
rect 51349 267338 51415 267341
rect 52361 267338 52427 267341
rect 64873 267338 64939 267341
rect 115933 267340 115999 267341
rect 115933 267338 115980 267340
rect 51349 267336 64939 267338
rect -960 267052 480 267292
rect 51349 267280 51354 267336
rect 51410 267280 52366 267336
rect 52422 267280 64878 267336
rect 64934 267280 64939 267336
rect 51349 267278 64939 267280
rect 115888 267336 115980 267338
rect 115888 267280 115938 267336
rect 115888 267278 115980 267280
rect 51349 267275 51415 267278
rect 52361 267275 52427 267278
rect 64873 267275 64939 267278
rect 115933 267276 115980 267278
rect 116044 267276 116050 267340
rect 183134 267276 183140 267340
rect 183204 267338 183210 267340
rect 183277 267338 183343 267341
rect 183204 267336 183343 267338
rect 183204 267280 183282 267336
rect 183338 267280 183343 267336
rect 183204 267278 183343 267280
rect 183204 267276 183210 267278
rect 115933 267275 115999 267276
rect 183277 267275 183343 267278
rect 212073 267338 212139 267341
rect 313406 267338 313412 267340
rect 212073 267336 313412 267338
rect 212073 267280 212078 267336
rect 212134 267280 313412 267336
rect 212073 267278 313412 267280
rect 212073 267275 212139 267278
rect 313406 267276 313412 267278
rect 313476 267276 313482 267340
rect 343214 267276 343220 267340
rect 343284 267338 343290 267340
rect 343541 267338 343607 267341
rect 343284 267336 343607 267338
rect 343284 267280 343546 267336
rect 343602 267280 343607 267336
rect 343284 267278 343607 267280
rect 343284 267276 343290 267278
rect 343541 267275 343607 267278
rect 379462 267276 379468 267340
rect 379532 267338 379538 267340
rect 428222 267338 428228 267340
rect 379532 267278 428228 267338
rect 379532 267276 379538 267278
rect 428222 267276 428228 267278
rect 428292 267276 428298 267340
rect 437473 267338 437539 267341
rect 438526 267338 438532 267340
rect 437473 267336 438532 267338
rect 437473 267280 437478 267336
rect 437534 267280 438532 267336
rect 437473 267278 438532 267280
rect 437473 267275 437539 267278
rect 438526 267276 438532 267278
rect 438596 267276 438602 267340
rect 442993 267338 443059 267341
rect 443494 267338 443500 267340
rect 442993 267336 443500 267338
rect 442993 267280 442998 267336
rect 443054 267280 443500 267336
rect 442993 267278 443500 267280
rect 442993 267275 443059 267278
rect 443494 267276 443500 267278
rect 443564 267276 443570 267340
rect 503110 267276 503116 267340
rect 503180 267338 503186 267340
rect 503437 267338 503503 267341
rect 503180 267336 503503 267338
rect 503180 267280 503442 267336
rect 503498 267280 503503 267336
rect 503180 267278 503503 267280
rect 503180 267276 503186 267278
rect 503437 267275 503503 267278
rect 47853 267202 47919 267205
rect 59813 267202 59879 267205
rect 88333 267204 88399 267205
rect 88333 267202 88380 267204
rect 47853 267200 59879 267202
rect 47853 267144 47858 267200
rect 47914 267144 59818 267200
rect 59874 267144 59879 267200
rect 47853 267142 59879 267144
rect 88288 267200 88380 267202
rect 88288 267144 88338 267200
rect 88288 267142 88380 267144
rect 47853 267139 47919 267142
rect 59813 267139 59879 267142
rect 88333 267140 88380 267142
rect 88444 267140 88450 267204
rect 100753 267202 100819 267205
rect 101070 267202 101076 267204
rect 100753 267200 101076 267202
rect 100753 267144 100758 267200
rect 100814 267144 101076 267200
rect 100753 267142 101076 267144
rect 88333 267139 88399 267140
rect 100753 267139 100819 267142
rect 101070 267140 101076 267142
rect 101140 267140 101146 267204
rect 104893 267202 104959 267205
rect 105854 267202 105860 267204
rect 104893 267200 105860 267202
rect 104893 267144 104898 267200
rect 104954 267144 105860 267200
rect 104893 267142 105860 267144
rect 104893 267139 104959 267142
rect 105854 267140 105860 267142
rect 105924 267140 105930 267204
rect 216397 267202 216463 267205
rect 238150 267202 238156 267204
rect 216397 267200 238156 267202
rect 216397 267144 216402 267200
rect 216458 267144 238156 267200
rect 216397 267142 238156 267144
rect 216397 267139 216463 267142
rect 238150 267140 238156 267142
rect 238220 267140 238226 267204
rect 258257 267202 258323 267205
rect 269757 267204 269823 267205
rect 271229 267204 271295 267205
rect 258390 267202 258396 267204
rect 258257 267200 258396 267202
rect 258257 267144 258262 267200
rect 258318 267144 258396 267200
rect 258257 267142 258396 267144
rect 258257 267139 258323 267142
rect 258390 267140 258396 267142
rect 258460 267140 258466 267204
rect 269757 267200 269804 267204
rect 269868 267202 269874 267204
rect 269757 267144 269762 267200
rect 269757 267140 269804 267144
rect 269868 267142 269914 267202
rect 271229 267200 271276 267204
rect 271340 267202 271346 267204
rect 271229 267144 271234 267200
rect 269868 267140 269874 267142
rect 271229 267140 271276 267144
rect 271340 267142 271386 267202
rect 271340 267140 271346 267142
rect 276974 267140 276980 267204
rect 277044 267202 277050 267204
rect 277117 267202 277183 267205
rect 278129 267204 278195 267205
rect 278078 267202 278084 267204
rect 277044 267200 277183 267202
rect 277044 267144 277122 267200
rect 277178 267144 277183 267200
rect 277044 267142 277183 267144
rect 278038 267142 278084 267202
rect 278148 267200 278195 267204
rect 278190 267144 278195 267200
rect 277044 267140 277050 267142
rect 269757 267139 269823 267140
rect 271229 267139 271295 267140
rect 277117 267139 277183 267142
rect 278078 267140 278084 267142
rect 278148 267140 278195 267144
rect 278129 267139 278195 267140
rect 375189 267202 375255 267205
rect 397126 267202 397132 267204
rect 375189 267200 397132 267202
rect 375189 267144 375194 267200
rect 375250 267144 397132 267200
rect 375189 267142 397132 267144
rect 375189 267139 375255 267142
rect 397126 267140 397132 267142
rect 397196 267140 397202 267204
rect 440233 267202 440299 267205
rect 440918 267202 440924 267204
rect 440233 267200 440924 267202
rect 440233 267144 440238 267200
rect 440294 267144 440924 267200
rect 440233 267142 440924 267144
rect 440233 267139 440299 267142
rect 440918 267140 440924 267142
rect 440988 267140 440994 267204
rect 43529 267066 43595 267069
rect 58617 267066 58683 267069
rect 103830 267066 103836 267068
rect 43529 267064 103836 267066
rect 43529 267008 43534 267064
rect 43590 267008 58622 267064
rect 58678 267008 103836 267064
rect 43529 267006 103836 267008
rect 43529 267003 43595 267006
rect 58617 267003 58683 267006
rect 103830 267004 103836 267006
rect 103900 267004 103906 267068
rect 215109 267066 215175 267069
rect 236494 267066 236500 267068
rect 215109 267064 236500 267066
rect 215109 267008 215114 267064
rect 215170 267008 236500 267064
rect 215109 267006 236500 267008
rect 215109 267003 215175 267006
rect 236494 267004 236500 267006
rect 236564 267004 236570 267068
rect 255313 267066 255379 267069
rect 273253 267068 273319 267069
rect 256182 267066 256188 267068
rect 255313 267064 256188 267066
rect 255313 267008 255318 267064
rect 255374 267008 256188 267064
rect 255313 267006 256188 267008
rect 255313 267003 255379 267006
rect 256182 267004 256188 267006
rect 256252 267004 256258 267068
rect 273253 267066 273300 267068
rect 273208 267064 273300 267066
rect 273208 267008 273258 267064
rect 273208 267006 273300 267008
rect 273253 267004 273300 267006
rect 273364 267004 273370 267068
rect 379973 267066 380039 267069
rect 396206 267066 396212 267068
rect 379973 267064 396212 267066
rect 379973 267008 379978 267064
rect 380034 267008 396212 267064
rect 379973 267006 396212 267008
rect 273253 267003 273319 267004
rect 379973 267003 380039 267006
rect 396206 267004 396212 267006
rect 396276 267004 396282 267068
rect 407113 267066 407179 267069
rect 408166 267066 408172 267068
rect 407113 267064 408172 267066
rect 407113 267008 407118 267064
rect 407174 267008 408172 267064
rect 407113 267006 408172 267008
rect 407113 267003 407179 267006
rect 408166 267004 408172 267006
rect 408236 267004 408242 267068
rect 409873 267066 409939 267069
rect 410742 267066 410748 267068
rect 409873 267064 410748 267066
rect 409873 267008 409878 267064
rect 409934 267008 410748 267064
rect 409873 267006 410748 267008
rect 409873 267003 409939 267006
rect 410742 267004 410748 267006
rect 410812 267004 410818 267068
rect 412909 267066 412975 267069
rect 413686 267066 413692 267068
rect 412909 267064 413692 267066
rect 412909 267008 412914 267064
rect 412970 267008 413692 267064
rect 412909 267006 413692 267008
rect 412909 267003 412975 267006
rect 413686 267004 413692 267006
rect 413756 267004 413762 267068
rect 422569 267066 422635 267069
rect 422886 267066 422892 267068
rect 422569 267064 422892 267066
rect 422569 267008 422574 267064
rect 422630 267008 422892 267064
rect 422569 267006 422892 267008
rect 422569 267003 422635 267006
rect 422886 267004 422892 267006
rect 422956 267004 422962 267068
rect 77293 266930 77359 266933
rect 78254 266930 78260 266932
rect 77293 266928 78260 266930
rect 77293 266872 77298 266928
rect 77354 266872 78260 266928
rect 77293 266870 78260 266872
rect 77293 266867 77359 266870
rect 78254 266868 78260 266870
rect 78324 266868 78330 266932
rect 80053 266930 80119 266933
rect 80462 266930 80468 266932
rect 80053 266928 80468 266930
rect 80053 266872 80058 266928
rect 80114 266872 80468 266928
rect 80053 266870 80468 266872
rect 80053 266867 80119 266870
rect 80462 266868 80468 266870
rect 80532 266868 80538 266932
rect 216489 266930 216555 266933
rect 237046 266930 237052 266932
rect 216489 266928 237052 266930
rect 216489 266872 216494 266928
rect 216550 266872 237052 266928
rect 216489 266870 237052 266872
rect 216489 266867 216555 266870
rect 237046 266868 237052 266870
rect 237116 266868 237122 266932
rect 247033 266930 247099 266933
rect 248270 266930 248276 266932
rect 247033 266928 248276 266930
rect 247033 266872 247038 266928
rect 247094 266872 248276 266928
rect 247033 266870 248276 266872
rect 247033 266867 247099 266870
rect 248270 266868 248276 266870
rect 248340 266868 248346 266932
rect 252553 266930 252619 266933
rect 253606 266930 253612 266932
rect 252553 266928 253612 266930
rect 252553 266872 252558 266928
rect 252614 266872 253612 266928
rect 252553 266870 253612 266872
rect 252553 266867 252619 266870
rect 253606 266868 253612 266870
rect 253676 266868 253682 266932
rect 263593 266930 263659 266933
rect 263910 266930 263916 266932
rect 263593 266928 263916 266930
rect 263593 266872 263598 266928
rect 263654 266872 263916 266928
rect 263593 266870 263916 266872
rect 263593 266867 263659 266870
rect 263910 266868 263916 266870
rect 263980 266868 263986 266932
rect 267733 266930 267799 266933
rect 268694 266930 268700 266932
rect 267733 266928 268700 266930
rect 267733 266872 267738 266928
rect 267794 266872 268700 266928
rect 267733 266870 268700 266872
rect 267733 266867 267799 266870
rect 268694 266868 268700 266870
rect 268764 266868 268770 266932
rect 310513 266930 310579 266933
rect 311014 266930 311020 266932
rect 310513 266928 311020 266930
rect 310513 266872 310518 266928
rect 310574 266872 311020 266928
rect 310513 266870 311020 266872
rect 310513 266867 310579 266870
rect 311014 266868 311020 266870
rect 311084 266868 311090 266932
rect 373533 266930 373599 266933
rect 462630 266930 462636 266932
rect 373533 266928 462636 266930
rect 373533 266872 373538 266928
rect 373594 266872 462636 266928
rect 373533 266870 462636 266872
rect 373533 266867 373599 266870
rect 462630 266868 462636 266870
rect 462700 266868 462706 266932
rect 200757 266794 200823 266797
rect 326654 266794 326660 266796
rect 200757 266792 326660 266794
rect 200757 266736 200762 266792
rect 200818 266736 326660 266792
rect 200757 266734 326660 266736
rect 200757 266731 200823 266734
rect 326654 266732 326660 266734
rect 326724 266732 326730 266796
rect 91093 266658 91159 266661
rect 91318 266658 91324 266660
rect 91093 266656 91324 266658
rect 91093 266600 91098 266656
rect 91154 266600 91324 266656
rect 91093 266598 91324 266600
rect 91093 266595 91159 266598
rect 91318 266596 91324 266598
rect 91388 266596 91394 266660
rect 100753 266524 100819 266525
rect 100702 266460 100708 266524
rect 100772 266522 100819 266524
rect 100772 266520 100864 266522
rect 100814 266464 100864 266520
rect 100772 266462 100864 266464
rect 100772 266460 100819 266462
rect 244222 266460 244228 266524
rect 244292 266522 244298 266524
rect 244365 266522 244431 266525
rect 244292 266520 244431 266522
rect 244292 266464 244370 266520
rect 244426 266464 244431 266520
rect 244292 266462 244431 266464
rect 244292 266460 244298 266462
rect 100753 266459 100819 266460
rect 244365 266459 244431 266462
rect 251265 266522 251331 266525
rect 252318 266522 252324 266524
rect 251265 266520 252324 266522
rect 251265 266464 251270 266520
rect 251326 266464 252324 266520
rect 251265 266462 252324 266464
rect 251265 266459 251331 266462
rect 252318 266460 252324 266462
rect 252388 266460 252394 266524
rect 259545 266522 259611 266525
rect 260598 266522 260604 266524
rect 259545 266520 260604 266522
rect 259545 266464 259550 266520
rect 259606 266464 260604 266520
rect 259545 266462 260604 266464
rect 259545 266459 259611 266462
rect 260598 266460 260604 266462
rect 260668 266460 260674 266524
rect 411345 266522 411411 266525
rect 412398 266522 412404 266524
rect 411345 266520 412404 266522
rect 411345 266464 411350 266520
rect 411406 266464 412404 266520
rect 411345 266462 412404 266464
rect 411345 266459 411411 266462
rect 412398 266460 412404 266462
rect 412468 266460 412474 266524
rect 418245 266522 418311 266525
rect 419206 266522 419212 266524
rect 418245 266520 419212 266522
rect 418245 266464 418250 266520
rect 418306 266464 419212 266520
rect 418245 266462 419212 266464
rect 418245 266459 418311 266462
rect 419206 266460 419212 266462
rect 419276 266460 419282 266524
rect 59813 266386 59879 266389
rect 62113 266386 62179 266389
rect 59813 266384 62179 266386
rect 59813 266328 59818 266384
rect 59874 266328 62118 266384
rect 62174 266328 62179 266384
rect 59813 266326 62179 266328
rect 59813 266323 59879 266326
rect 62113 266323 62179 266326
rect 85573 266386 85639 266389
rect 86534 266386 86540 266388
rect 85573 266384 86540 266386
rect 85573 266328 85578 266384
rect 85634 266328 86540 266384
rect 85573 266326 86540 266328
rect 85573 266323 85639 266326
rect 86534 266324 86540 266326
rect 86604 266324 86610 266388
rect 88333 266386 88399 266389
rect 88742 266386 88748 266388
rect 88333 266384 88748 266386
rect 88333 266328 88338 266384
rect 88394 266328 88748 266384
rect 88333 266326 88748 266328
rect 88333 266323 88399 266326
rect 88742 266324 88748 266326
rect 88812 266324 88818 266388
rect 89713 266386 89779 266389
rect 90030 266386 90036 266388
rect 89713 266384 90036 266386
rect 89713 266328 89718 266384
rect 89774 266328 90036 266384
rect 89713 266326 90036 266328
rect 89713 266323 89779 266326
rect 90030 266324 90036 266326
rect 90100 266324 90106 266388
rect 92473 266386 92539 266389
rect 93342 266386 93348 266388
rect 92473 266384 93348 266386
rect 92473 266328 92478 266384
rect 92534 266328 93348 266384
rect 92473 266326 93348 266328
rect 92473 266323 92539 266326
rect 93342 266324 93348 266326
rect 93412 266324 93418 266388
rect 96613 266386 96679 266389
rect 97022 266386 97028 266388
rect 96613 266384 97028 266386
rect 96613 266328 96618 266384
rect 96674 266328 97028 266384
rect 96613 266326 97028 266328
rect 96613 266323 96679 266326
rect 97022 266324 97028 266326
rect 97092 266324 97098 266388
rect 97993 266386 98059 266389
rect 98126 266386 98132 266388
rect 97993 266384 98132 266386
rect 97993 266328 97998 266384
rect 98054 266328 98132 266384
rect 97993 266326 98132 266328
rect 97993 266323 98059 266326
rect 98126 266324 98132 266326
rect 98196 266324 98202 266388
rect 100845 266386 100911 266389
rect 101806 266386 101812 266388
rect 100845 266384 101812 266386
rect 100845 266328 100850 266384
rect 100906 266328 101812 266384
rect 100845 266326 101812 266328
rect 100845 266323 100911 266326
rect 101806 266324 101812 266326
rect 101876 266324 101882 266388
rect 111793 266386 111859 266389
rect 112110 266386 112116 266388
rect 111793 266384 112116 266386
rect 111793 266328 111798 266384
rect 111854 266328 112116 266384
rect 111793 266326 112116 266328
rect 111793 266323 111859 266326
rect 112110 266324 112116 266326
rect 112180 266324 112186 266388
rect 114502 266324 114508 266388
rect 114572 266324 114578 266388
rect 147673 266386 147739 266389
rect 148542 266386 148548 266388
rect 147673 266384 148548 266386
rect 147673 266328 147678 266384
rect 147734 266328 148548 266384
rect 147673 266326 148548 266328
rect 114510 266250 114570 266324
rect 147673 266323 147739 266326
rect 148542 266324 148548 266326
rect 148612 266324 148618 266388
rect 215569 266386 215635 266389
rect 216489 266386 216555 266389
rect 215569 266384 216555 266386
rect 215569 266328 215574 266384
rect 215630 266328 216494 266384
rect 216550 266328 216555 266384
rect 215569 266326 216555 266328
rect 215569 266323 215635 266326
rect 216489 266323 216555 266326
rect 244273 266386 244339 266389
rect 245326 266386 245332 266388
rect 244273 266384 245332 266386
rect 244273 266328 244278 266384
rect 244334 266328 245332 266384
rect 244273 266326 245332 266328
rect 244273 266323 244339 266326
rect 245326 266324 245332 266326
rect 245396 266324 245402 266388
rect 245653 266386 245719 266389
rect 246430 266386 246436 266388
rect 245653 266384 246436 266386
rect 245653 266328 245658 266384
rect 245714 266328 246436 266384
rect 245653 266326 246436 266328
rect 245653 266323 245719 266326
rect 246430 266324 246436 266326
rect 246500 266324 246506 266388
rect 247033 266386 247099 266389
rect 247718 266386 247724 266388
rect 247033 266384 247724 266386
rect 247033 266328 247038 266384
rect 247094 266328 247724 266384
rect 247033 266326 247724 266328
rect 247033 266323 247099 266326
rect 247718 266324 247724 266326
rect 247788 266324 247794 266388
rect 248505 266386 248571 266389
rect 248638 266386 248644 266388
rect 248505 266384 248644 266386
rect 248505 266328 248510 266384
rect 248566 266328 248644 266384
rect 248505 266326 248644 266328
rect 248505 266323 248571 266326
rect 248638 266324 248644 266326
rect 248708 266324 248714 266388
rect 249793 266386 249859 266389
rect 251173 266388 251239 266389
rect 250110 266386 250116 266388
rect 249793 266384 250116 266386
rect 249793 266328 249798 266384
rect 249854 266328 250116 266384
rect 249793 266326 250116 266328
rect 249793 266323 249859 266326
rect 250110 266324 250116 266326
rect 250180 266324 250186 266388
rect 251173 266386 251220 266388
rect 251128 266384 251220 266386
rect 251128 266328 251178 266384
rect 251128 266326 251220 266328
rect 251173 266324 251220 266326
rect 251284 266324 251290 266388
rect 252553 266386 252619 266389
rect 253422 266386 253428 266388
rect 252553 266384 253428 266386
rect 252553 266328 252558 266384
rect 252614 266328 253428 266384
rect 252553 266326 253428 266328
rect 251173 266323 251239 266324
rect 252553 266323 252619 266326
rect 253422 266324 253428 266326
rect 253492 266324 253498 266388
rect 253933 266386 253999 266389
rect 254526 266386 254532 266388
rect 253933 266384 254532 266386
rect 253933 266328 253938 266384
rect 253994 266328 254532 266384
rect 253933 266326 254532 266328
rect 253933 266323 253999 266326
rect 254526 266324 254532 266326
rect 254596 266324 254602 266388
rect 256693 266386 256759 266389
rect 259453 266388 259519 266389
rect 256918 266386 256924 266388
rect 256693 266384 256924 266386
rect 256693 266328 256698 266384
rect 256754 266328 256924 266384
rect 256693 266326 256924 266328
rect 256693 266323 256759 266326
rect 256918 266324 256924 266326
rect 256988 266324 256994 266388
rect 259453 266386 259500 266388
rect 259408 266384 259500 266386
rect 259408 266328 259458 266384
rect 259408 266326 259500 266328
rect 259453 266324 259500 266326
rect 259564 266324 259570 266388
rect 262213 266386 262279 266389
rect 262806 266386 262812 266388
rect 262213 266384 262812 266386
rect 262213 266328 262218 266384
rect 262274 266328 262812 266384
rect 262213 266326 262812 266328
rect 259453 266323 259519 266324
rect 262213 266323 262279 266326
rect 262806 266324 262812 266326
rect 262876 266324 262882 266388
rect 278998 266324 279004 266388
rect 279068 266386 279074 266388
rect 279969 266386 280035 266389
rect 279068 266384 280035 266386
rect 279068 266328 279974 266384
rect 280030 266328 280035 266384
rect 279068 266326 280035 266328
rect 279068 266324 279074 266326
rect 279969 266323 280035 266326
rect 374361 266386 374427 266389
rect 375189 266386 375255 266389
rect 374361 266384 375255 266386
rect 374361 266328 374366 266384
rect 374422 266328 375194 266384
rect 375250 266328 375255 266384
rect 374361 266326 375255 266328
rect 374361 266323 374427 266326
rect 375189 266323 375255 266326
rect 398833 266386 398899 266389
rect 399518 266386 399524 266388
rect 398833 266384 399524 266386
rect 398833 266328 398838 266384
rect 398894 266328 399524 266384
rect 398833 266326 399524 266328
rect 398833 266323 398899 266326
rect 399518 266324 399524 266326
rect 399588 266324 399594 266388
rect 400213 266386 400279 266389
rect 400438 266386 400444 266388
rect 400213 266384 400444 266386
rect 400213 266328 400218 266384
rect 400274 266328 400444 266384
rect 400213 266326 400444 266328
rect 400213 266323 400279 266326
rect 400438 266324 400444 266326
rect 400508 266324 400514 266388
rect 403157 266386 403223 266389
rect 404118 266386 404124 266388
rect 403157 266384 404124 266386
rect 403157 266328 403162 266384
rect 403218 266328 404124 266384
rect 403157 266326 404124 266328
rect 403157 266323 403223 266326
rect 404118 266324 404124 266326
rect 404188 266324 404194 266388
rect 404353 266386 404419 266389
rect 405038 266386 405044 266388
rect 404353 266384 405044 266386
rect 404353 266328 404358 266384
rect 404414 266328 405044 266384
rect 404353 266326 405044 266328
rect 404353 266323 404419 266326
rect 405038 266324 405044 266326
rect 405108 266324 405114 266388
rect 405733 266386 405799 266389
rect 406510 266386 406516 266388
rect 405733 266384 406516 266386
rect 405733 266328 405738 266384
rect 405794 266328 406516 266384
rect 405733 266326 406516 266328
rect 405733 266323 405799 266326
rect 406510 266324 406516 266326
rect 406580 266324 406586 266388
rect 407113 266386 407179 266389
rect 407614 266386 407620 266388
rect 407113 266384 407620 266386
rect 407113 266328 407118 266384
rect 407174 266328 407620 266384
rect 407113 266326 407620 266328
rect 407113 266323 407179 266326
rect 407614 266324 407620 266326
rect 407684 266324 407690 266388
rect 408493 266386 408559 266389
rect 408718 266386 408724 266388
rect 408493 266384 408724 266386
rect 408493 266328 408498 266384
rect 408554 266328 408724 266384
rect 408493 266326 408724 266328
rect 408493 266323 408559 266326
rect 408718 266324 408724 266326
rect 408788 266324 408794 266388
rect 409873 266386 409939 266389
rect 411253 266388 411319 266389
rect 410006 266386 410012 266388
rect 409873 266384 410012 266386
rect 409873 266328 409878 266384
rect 409934 266328 410012 266384
rect 409873 266326 410012 266328
rect 409873 266323 409939 266326
rect 410006 266324 410012 266326
rect 410076 266324 410082 266388
rect 411253 266386 411300 266388
rect 411208 266384 411300 266386
rect 411208 266328 411258 266384
rect 411208 266326 411300 266328
rect 411253 266324 411300 266326
rect 411364 266324 411370 266388
rect 412909 266386 412975 266389
rect 413318 266386 413324 266388
rect 412909 266384 413324 266386
rect 412909 266328 412914 266384
rect 412970 266328 413324 266384
rect 412909 266326 413324 266328
rect 411253 266323 411319 266324
rect 412909 266323 412975 266326
rect 413318 266324 413324 266326
rect 413388 266324 413394 266388
rect 416773 266386 416839 266389
rect 418153 266388 418219 266389
rect 416998 266386 417004 266388
rect 416773 266384 417004 266386
rect 416773 266328 416778 266384
rect 416834 266328 417004 266384
rect 416773 266326 417004 266328
rect 416773 266323 416839 266326
rect 416998 266324 417004 266326
rect 417068 266324 417074 266388
rect 418102 266324 418108 266388
rect 418172 266386 418219 266388
rect 419533 266386 419599 266389
rect 420678 266386 420684 266388
rect 418172 266384 418264 266386
rect 418214 266328 418264 266384
rect 418172 266326 418264 266328
rect 419533 266384 420684 266386
rect 419533 266328 419538 266384
rect 419594 266328 420684 266384
rect 419533 266326 420684 266328
rect 418172 266324 418219 266326
rect 418153 266323 418219 266324
rect 419533 266323 419599 266326
rect 420678 266324 420684 266326
rect 420748 266324 420754 266388
rect 420913 266386 420979 266389
rect 421782 266386 421788 266388
rect 420913 266384 421788 266386
rect 420913 266328 420918 266384
rect 420974 266328 421788 266384
rect 420913 266326 421788 266328
rect 420913 266323 420979 266326
rect 421782 266324 421788 266326
rect 421852 266324 421858 266388
rect 428774 266324 428780 266388
rect 428844 266386 428850 266388
rect 429101 266386 429167 266389
rect 428844 266384 429167 266386
rect 428844 266328 429106 266384
rect 429162 266328 429167 266384
rect 428844 266326 429167 266328
rect 428844 266324 428850 266326
rect 429101 266323 429167 266326
rect 429878 266324 429884 266388
rect 429948 266386 429954 266388
rect 430481 266386 430547 266389
rect 429948 266384 430547 266386
rect 429948 266328 430486 266384
rect 430542 266328 430547 266384
rect 429948 266326 430547 266328
rect 429948 266324 429954 266326
rect 430481 266323 430547 266326
rect 430665 266386 430731 266389
rect 431166 266386 431172 266388
rect 430665 266384 431172 266386
rect 430665 266328 430670 266384
rect 430726 266328 431172 266384
rect 430665 266326 431172 266328
rect 430665 266323 430731 266326
rect 431166 266324 431172 266326
rect 431236 266324 431242 266388
rect 436093 266386 436159 266389
rect 436870 266386 436876 266388
rect 436093 266384 436876 266386
rect 436093 266328 436098 266384
rect 436154 266328 436876 266384
rect 436093 266326 436876 266328
rect 436093 266323 436159 266326
rect 436870 266324 436876 266326
rect 436940 266324 436946 266388
rect 437473 266386 437539 266389
rect 438342 266386 438348 266388
rect 437473 266384 438348 266386
rect 437473 266328 437478 266384
rect 437534 266328 438348 266384
rect 437473 266326 438348 266328
rect 437473 266323 437539 266326
rect 438342 266324 438348 266326
rect 438412 266324 438418 266388
rect 438853 266386 438919 266389
rect 439078 266386 439084 266388
rect 438853 266384 439084 266386
rect 438853 266328 438858 266384
rect 438914 266328 439084 266384
rect 438853 266326 439084 266328
rect 438853 266323 438919 266326
rect 439078 266324 439084 266326
rect 439148 266324 439154 266388
rect 196750 266250 196756 266252
rect 114510 266190 196756 266250
rect 196750 266188 196756 266190
rect 196820 266188 196826 266252
rect 239254 266250 239260 266252
rect 229050 266190 239260 266250
rect 217542 265916 217548 265980
rect 217612 265978 217618 265980
rect 219617 265978 219683 265981
rect 220721 265978 220787 265981
rect 217612 265976 220787 265978
rect 217612 265920 219622 265976
rect 219678 265920 220726 265976
rect 220782 265920 220787 265976
rect 217612 265918 220787 265920
rect 217612 265916 217618 265918
rect 219617 265915 219683 265918
rect 220721 265915 220787 265918
rect 212073 265842 212139 265845
rect 229050 265842 229110 266190
rect 239254 266188 239260 266190
rect 239324 266188 239330 266252
rect 212073 265840 229110 265842
rect 212073 265784 212078 265840
rect 212134 265784 229110 265840
rect 212073 265782 229110 265784
rect 212073 265779 212139 265782
rect 212441 265706 212507 265709
rect 240542 265706 240548 265708
rect 212441 265704 240548 265706
rect 212441 265648 212446 265704
rect 212502 265648 240548 265704
rect 212441 265646 240548 265648
rect 212441 265643 212507 265646
rect 240542 265644 240548 265646
rect 240612 265644 240618 265708
rect 208945 265570 209011 265573
rect 212165 265570 212231 265573
rect 241646 265570 241652 265572
rect 208945 265568 241652 265570
rect 208945 265512 208950 265568
rect 209006 265512 212170 265568
rect 212226 265512 241652 265568
rect 208945 265510 241652 265512
rect 208945 265507 209011 265510
rect 212165 265507 212231 265510
rect 241646 265508 241652 265510
rect 241716 265508 241722 265572
rect 378961 265570 379027 265573
rect 427670 265570 427676 265572
rect 378961 265568 427676 265570
rect 378961 265512 378966 265568
rect 379022 265512 427676 265568
rect 378961 265510 427676 265512
rect 378961 265507 379027 265510
rect 427670 265508 427676 265510
rect 427740 265508 427746 265572
rect 371785 265298 371851 265301
rect 376477 265298 376543 265301
rect 388161 265298 388227 265301
rect 371785 265296 388227 265298
rect 371785 265240 371790 265296
rect 371846 265240 376482 265296
rect 376538 265240 388166 265296
rect 388222 265240 388227 265296
rect 371785 265238 388227 265240
rect 371785 265235 371851 265238
rect 376477 265235 376543 265238
rect 388161 265235 388227 265238
rect 210693 265162 210759 265165
rect 216397 265162 216463 265165
rect 210693 265160 216463 265162
rect 210693 265104 210698 265160
rect 210754 265104 216402 265160
rect 216458 265104 216463 265160
rect 210693 265102 216463 265104
rect 210693 265099 210759 265102
rect 216397 265099 216463 265102
rect 375373 265162 375439 265165
rect 375833 265162 375899 265165
rect 389173 265162 389239 265165
rect 375373 265160 389239 265162
rect 375373 265104 375378 265160
rect 375434 265104 375838 265160
rect 375894 265104 389178 265160
rect 389234 265104 389239 265160
rect 375373 265102 389239 265104
rect 375373 265099 375439 265102
rect 375833 265099 375899 265102
rect 389173 265099 389239 265102
rect 210969 265026 211035 265029
rect 212073 265026 212139 265029
rect 210969 265024 212139 265026
rect 210969 264968 210974 265024
rect 211030 264968 212078 265024
rect 212134 264968 212139 265024
rect 210969 264966 212139 264968
rect 210969 264963 211035 264966
rect 212073 264963 212139 264966
rect 212441 265026 212507 265029
rect 213085 265026 213151 265029
rect 212441 265024 213151 265026
rect 212441 264968 212446 265024
rect 212502 264968 213090 265024
rect 213146 264968 213151 265024
rect 212441 264966 213151 264968
rect 212441 264963 212507 264966
rect 213085 264963 213151 264966
rect 375465 265026 375531 265029
rect 375925 265026 375991 265029
rect 390553 265026 390619 265029
rect 375465 265024 390619 265026
rect 375465 264968 375470 265024
rect 375526 264968 375930 265024
rect 375986 264968 390558 265024
rect 390614 264968 390619 265024
rect 375465 264966 390619 264968
rect 375465 264963 375531 264966
rect 375925 264963 375991 264966
rect 390553 264963 390619 264966
rect 47894 264828 47900 264892
rect 47964 264890 47970 264892
rect 52729 264890 52795 264893
rect 53189 264890 53255 264893
rect 47964 264888 53255 264890
rect 47964 264832 52734 264888
rect 52790 264832 53194 264888
rect 53250 264832 53255 264888
rect 47964 264830 53255 264832
rect 47964 264828 47970 264830
rect 52729 264827 52795 264830
rect 53189 264827 53255 264830
rect 377806 263468 377812 263532
rect 377876 263530 377882 263532
rect 378041 263530 378107 263533
rect 377876 263528 378107 263530
rect 377876 263472 378046 263528
rect 378102 263472 378107 263528
rect 377876 263470 378107 263472
rect 377876 263468 377882 263470
rect 378041 263467 378107 263470
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect -960 254086 6930 254146
rect -960 253996 480 254086
rect 6870 254010 6930 254086
rect 53046 254010 53052 254012
rect 6870 253950 53052 254010
rect 53046 253948 53052 253950
rect 53116 253948 53122 254012
rect 215334 251092 215340 251156
rect 215404 251154 215410 251156
rect 216489 251154 216555 251157
rect 215404 251152 216555 251154
rect 215404 251096 216494 251152
rect 216550 251096 216555 251152
rect 215404 251094 216555 251096
rect 215404 251092 215410 251094
rect 216489 251091 216555 251094
rect 178534 249868 178540 249932
rect 178604 249930 178610 249932
rect 179321 249930 179387 249933
rect 178604 249928 179387 249930
rect 178604 249872 179326 249928
rect 179382 249872 179387 249928
rect 178604 249870 179387 249872
rect 178604 249868 178610 249870
rect 179321 249867 179387 249870
rect 179638 249868 179644 249932
rect 179708 249930 179714 249932
rect 180241 249930 180307 249933
rect 190913 249932 190979 249933
rect 338481 249932 338547 249933
rect 190862 249930 190868 249932
rect 179708 249928 180307 249930
rect 179708 249872 180246 249928
rect 180302 249872 180307 249928
rect 179708 249870 180307 249872
rect 190822 249870 190868 249930
rect 190932 249928 190979 249932
rect 338430 249930 338436 249932
rect 190974 249872 190979 249928
rect 179708 249868 179714 249870
rect 180241 249867 180307 249870
rect 190862 249868 190868 249870
rect 190932 249868 190979 249872
rect 338390 249870 338436 249930
rect 338500 249928 338547 249932
rect 338542 249872 338547 249928
rect 338430 249868 338436 249870
rect 338500 249868 338547 249872
rect 339718 249868 339724 249932
rect 339788 249930 339794 249932
rect 340229 249930 340295 249933
rect 350993 249932 351059 249933
rect 350942 249930 350948 249932
rect 339788 249928 340295 249930
rect 339788 249872 340234 249928
rect 340290 249872 340295 249928
rect 339788 249870 340295 249872
rect 350902 249870 350948 249930
rect 351012 249928 351059 249932
rect 351054 249872 351059 249928
rect 339788 249868 339794 249870
rect 190913 249867 190979 249868
rect 338481 249867 338547 249868
rect 340229 249867 340295 249870
rect 350942 249868 350948 249870
rect 351012 249868 351059 249872
rect 498510 249868 498516 249932
rect 498580 249930 498586 249932
rect 499021 249930 499087 249933
rect 498580 249928 499087 249930
rect 498580 249872 499026 249928
rect 499082 249872 499087 249928
rect 498580 249870 499087 249872
rect 498580 249868 498586 249870
rect 350993 249867 351059 249868
rect 499021 249867 499087 249870
rect 499798 249868 499804 249932
rect 499868 249930 499874 249932
rect 500401 249930 500467 249933
rect 510889 249932 510955 249933
rect 510838 249930 510844 249932
rect 499868 249928 500467 249930
rect 499868 249872 500406 249928
rect 500462 249872 500467 249928
rect 499868 249870 500467 249872
rect 510798 249870 510844 249930
rect 510908 249928 510955 249932
rect 510950 249872 510955 249928
rect 499868 249868 499874 249870
rect 500401 249867 500467 249870
rect 510838 249868 510844 249870
rect 510908 249868 510955 249872
rect 510889 249867 510955 249868
rect 583520 245428 584960 245668
rect 196604 244218 197186 244220
rect 198733 244218 198799 244221
rect 199193 244218 199259 244221
rect 518893 244218 518959 244221
rect 519353 244218 519419 244221
rect 196604 244216 199259 244218
rect 196604 244160 198738 244216
rect 198794 244160 199198 244216
rect 199254 244160 199259 244216
rect 516558 244216 519419 244218
rect 197126 244158 199259 244160
rect 198733 244155 198799 244158
rect 199193 244155 199259 244158
rect 356562 243810 356622 244190
rect 516558 244160 518898 244216
rect 518954 244160 519358 244216
rect 519414 244160 519419 244216
rect 516558 244158 519419 244160
rect 518893 244155 518959 244158
rect 519353 244155 519419 244158
rect 358813 243810 358879 243813
rect 359273 243810 359339 243813
rect 356562 243808 359339 243810
rect 356562 243752 358818 243808
rect 358874 243752 359278 243808
rect 359334 243752 359339 243808
rect 356562 243750 359339 243752
rect 358813 243747 358879 243750
rect 359273 243747 359339 243750
rect -960 240940 480 241180
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect 216673 202874 216739 202877
rect 216857 202874 216923 202877
rect 216673 202872 216923 202874
rect 216673 202816 216678 202872
rect 216734 202816 216862 202872
rect 216918 202816 216923 202872
rect 216673 202814 216923 202816
rect 216673 202811 216739 202814
rect 216857 202811 216923 202814
rect 376845 202874 376911 202877
rect 377489 202874 377555 202877
rect 376845 202872 377555 202874
rect 376845 202816 376850 202872
rect 376906 202816 377494 202872
rect 377550 202816 377555 202872
rect 376845 202814 377555 202816
rect 376845 202811 376911 202814
rect 377489 202811 377555 202814
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 57053 201922 57119 201925
rect 216857 201922 216923 201925
rect 219390 201922 220064 201924
rect 57053 201920 60062 201922
rect 57053 201864 57058 201920
rect 57114 201864 60062 201920
rect 57053 201862 60062 201864
rect 216857 201920 220064 201922
rect 216857 201864 216862 201920
rect 216918 201864 220064 201920
rect 377489 201922 377555 201925
rect 379470 201922 380052 201924
rect 377489 201920 380052 201922
rect 377489 201864 377494 201920
rect 377550 201864 380052 201920
rect 216857 201862 219450 201864
rect 377489 201862 379530 201864
rect 57053 201859 57119 201862
rect 216857 201859 216923 201862
rect 377489 201859 377555 201862
rect 56869 201378 56935 201381
rect 57145 201378 57211 201381
rect 56869 201376 60062 201378
rect 56869 201320 56874 201376
rect 56930 201320 57150 201376
rect 57206 201320 60062 201376
rect 56869 201318 60062 201320
rect 56869 201315 56935 201318
rect 57145 201315 57211 201318
rect 60002 200942 60062 201318
rect 217041 200970 217107 200973
rect 219390 200970 220064 200972
rect 217041 200968 220064 200970
rect 217041 200912 217046 200968
rect 217102 200912 220064 200968
rect 376937 200970 377003 200973
rect 379470 200970 380052 200972
rect 376937 200968 380052 200970
rect 376937 200912 376942 200968
rect 376998 200912 380052 200968
rect 217041 200910 219450 200912
rect 376937 200910 379530 200912
rect 217041 200907 217107 200910
rect 376937 200907 377003 200910
rect 56869 198794 56935 198797
rect 57329 198794 57395 198797
rect 217685 198794 217751 198797
rect 217961 198794 218027 198797
rect 219390 198794 220064 198796
rect 56869 198792 60062 198794
rect 56869 198736 56874 198792
rect 56930 198736 57334 198792
rect 57390 198736 60062 198792
rect 56869 198734 60062 198736
rect 217685 198792 220064 198794
rect 217685 198736 217690 198792
rect 217746 198736 217966 198792
rect 218022 198736 220064 198792
rect 377213 198794 377279 198797
rect 377857 198794 377923 198797
rect 379470 198794 380052 198796
rect 377213 198792 380052 198794
rect 377213 198736 377218 198792
rect 377274 198736 377862 198792
rect 377918 198736 380052 198792
rect 217685 198734 219450 198736
rect 377213 198734 379530 198736
rect 56869 198731 56935 198734
rect 57329 198731 57395 198734
rect 217685 198731 217751 198734
rect 217961 198731 218027 198734
rect 377213 198731 377279 198734
rect 377857 198731 377923 198734
rect 217225 197842 217291 197845
rect 219390 197842 220064 197844
rect 217225 197840 220064 197842
rect 57329 197434 57395 197437
rect 57513 197434 57579 197437
rect 60002 197434 60062 197814
rect 217225 197784 217230 197840
rect 217286 197784 220064 197840
rect 377581 197842 377647 197845
rect 379470 197842 380052 197844
rect 377581 197840 380052 197842
rect 377581 197784 377586 197840
rect 377642 197784 380052 197840
rect 217225 197782 219450 197784
rect 377581 197782 379530 197784
rect 217225 197779 217291 197782
rect 377581 197779 377647 197782
rect 57329 197432 60062 197434
rect 57329 197376 57334 197432
rect 57390 197376 57518 197432
rect 57574 197376 60062 197432
rect 57329 197374 60062 197376
rect 57329 197371 57395 197374
rect 57513 197371 57579 197374
rect 57697 196074 57763 196077
rect 217501 196074 217567 196077
rect 217685 196074 217751 196077
rect 219390 196074 220064 196076
rect 57697 196072 60062 196074
rect 57697 196016 57702 196072
rect 57758 196016 60062 196072
rect 57697 196014 60062 196016
rect 217501 196072 220064 196074
rect 217501 196016 217506 196072
rect 217562 196016 217690 196072
rect 217746 196016 220064 196072
rect 376753 196074 376819 196077
rect 377765 196074 377831 196077
rect 379470 196074 380052 196076
rect 376753 196072 380052 196074
rect 376753 196016 376758 196072
rect 376814 196016 377770 196072
rect 377826 196016 380052 196072
rect 217501 196014 219450 196016
rect 376753 196014 379530 196016
rect 57697 196011 57763 196014
rect 217501 196011 217567 196014
rect 217685 196011 217751 196014
rect 376753 196011 376819 196014
rect 377765 196011 377831 196014
rect 56961 195258 57027 195261
rect 57513 195258 57579 195261
rect 56961 195256 60062 195258
rect 56961 195200 56966 195256
rect 57022 195200 57518 195256
rect 57574 195200 60062 195256
rect 56961 195198 60062 195200
rect 56961 195195 57027 195198
rect 57513 195195 57579 195198
rect 60002 194958 60062 195198
rect 217409 194986 217475 194989
rect 219390 194986 220064 194988
rect 217409 194984 220064 194986
rect 217409 194928 217414 194984
rect 217470 194928 220064 194984
rect 377305 194986 377371 194989
rect 379470 194986 380052 194988
rect 377305 194984 380052 194986
rect 377305 194928 377310 194984
rect 377366 194928 380052 194984
rect 217409 194926 219450 194928
rect 377305 194926 379530 194928
rect 217409 194923 217475 194926
rect 377305 194923 377371 194926
rect 57421 193218 57487 193221
rect 217593 193218 217659 193221
rect 219390 193218 220064 193220
rect 57421 193216 60062 193218
rect 57421 193160 57426 193216
rect 57482 193160 60062 193216
rect 57421 193158 60062 193160
rect 217593 193216 220064 193218
rect 217593 193160 217598 193216
rect 217654 193160 220064 193216
rect 377673 193218 377739 193221
rect 379470 193218 380052 193220
rect 377673 193216 380052 193218
rect 377673 193160 377678 193216
rect 377734 193160 380052 193216
rect 217593 193158 219450 193160
rect 377673 193158 379530 193160
rect 57421 193155 57487 193158
rect 217593 193155 217659 193158
rect 377673 193155 377739 193158
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 358997 184922 359063 184925
rect 359549 184922 359615 184925
rect 518893 184922 518959 184925
rect 519261 184922 519327 184925
rect 356562 184920 359615 184922
rect 356562 184864 359002 184920
rect 359058 184864 359554 184920
rect 359610 184864 359615 184920
rect 356562 184862 359615 184864
rect 196604 184378 197186 184380
rect 198825 184378 198891 184381
rect 199377 184378 199443 184381
rect 196604 184376 199443 184378
rect 196604 184320 198830 184376
rect 198886 184320 199382 184376
rect 199438 184320 199443 184376
rect 356562 184350 356622 184862
rect 358997 184859 359063 184862
rect 359549 184859 359615 184862
rect 516558 184920 519327 184922
rect 516558 184864 518898 184920
rect 518954 184864 519266 184920
rect 519322 184864 519327 184920
rect 516558 184862 519327 184864
rect 516558 184350 516618 184862
rect 518893 184859 518959 184862
rect 519261 184859 519327 184862
rect 197126 184318 199443 184320
rect 198825 184315 198891 184318
rect 199377 184315 199443 184318
rect 196604 182746 197186 182748
rect 199285 182746 199351 182749
rect 358905 182746 358971 182749
rect 518985 182746 519051 182749
rect 520181 182746 520247 182749
rect 196604 182744 199351 182746
rect 196604 182688 199290 182744
rect 199346 182688 199351 182744
rect 197126 182686 199351 182688
rect 356562 182744 358971 182746
rect 356562 182688 358910 182744
rect 358966 182688 358971 182744
rect 356562 182686 358971 182688
rect 516558 182744 520247 182746
rect 516558 182688 518990 182744
rect 519046 182688 520186 182744
rect 520242 182688 520247 182744
rect 516558 182686 520247 182688
rect 199285 182683 199351 182686
rect 358905 182683 358971 182686
rect 518985 182683 519051 182686
rect 520181 182683 520247 182686
rect 196604 181386 197186 181388
rect 199101 181386 199167 181389
rect 359181 181386 359247 181389
rect 519261 181386 519327 181389
rect 196604 181384 199167 181386
rect 196604 181328 199106 181384
rect 199162 181328 199167 181384
rect 197126 181326 199167 181328
rect 356562 181384 359247 181386
rect 356562 181328 359186 181384
rect 359242 181328 359247 181384
rect 356562 181326 359247 181328
rect 516558 181384 519327 181386
rect 516558 181328 519266 181384
rect 519322 181328 519327 181384
rect 516558 181326 519327 181328
rect 199101 181323 199167 181326
rect 359181 181323 359247 181326
rect 519261 181323 519327 181326
rect 196558 179482 196618 179862
rect 198733 179482 198799 179485
rect 199009 179482 199075 179485
rect 196558 179480 199075 179482
rect 196558 179424 198738 179480
rect 198794 179424 199014 179480
rect 199070 179424 199075 179480
rect 196558 179422 199075 179424
rect 356562 179482 356622 179862
rect 358905 179482 358971 179485
rect 359457 179482 359523 179485
rect 356562 179480 359523 179482
rect 356562 179424 358910 179480
rect 358966 179424 359462 179480
rect 359518 179424 359523 179480
rect 356562 179422 359523 179424
rect 516558 179482 516618 179862
rect 519077 179482 519143 179485
rect 519445 179482 519511 179485
rect 516558 179480 519511 179482
rect 516558 179424 519082 179480
rect 519138 179424 519450 179480
rect 519506 179424 519511 179480
rect 516558 179422 519511 179424
rect 198733 179419 198799 179422
rect 199009 179419 199075 179422
rect 358905 179419 358971 179422
rect 359457 179419 359523 179422
rect 519077 179419 519143 179422
rect 519445 179419 519511 179422
rect 583520 179060 584960 179300
rect 519077 178802 519143 178805
rect 516558 178800 519143 178802
rect 516558 178744 519082 178800
rect 519138 178744 519143 178800
rect 516558 178742 519143 178744
rect 196604 178666 197186 178668
rect 198825 178666 198891 178669
rect 196604 178664 198891 178666
rect 196604 178608 198830 178664
rect 198886 178608 198891 178664
rect 516558 178638 516618 178742
rect 519077 178739 519143 178742
rect 197126 178606 198891 178608
rect 198825 178603 198891 178606
rect 356562 178122 356622 178638
rect 359089 178122 359155 178125
rect 359365 178122 359431 178125
rect 356562 178120 359431 178122
rect 356562 178064 359094 178120
rect 359150 178064 359370 178120
rect 359426 178064 359431 178120
rect 356562 178062 359431 178064
rect 359089 178059 359155 178062
rect 359365 178059 359431 178062
rect -960 175796 480 176036
rect 58341 175266 58407 175269
rect 58566 175266 58572 175268
rect 58341 175264 58572 175266
rect 58341 175208 58346 175264
rect 58402 175208 58572 175264
rect 58341 175206 58572 175208
rect 58341 175203 58407 175206
rect 58566 175204 58572 175206
rect 58636 175204 58642 175268
rect 58985 175266 59051 175269
rect 58985 175264 60062 175266
rect 58985 175208 58990 175264
rect 59046 175208 60062 175264
rect 58985 175206 60062 175208
rect 58985 175203 59051 175206
rect 60002 174966 60062 175206
rect 216673 174994 216739 174997
rect 219390 174994 220064 174996
rect 216673 174992 220064 174994
rect 216673 174936 216678 174992
rect 216734 174936 220064 174992
rect 376845 174994 376911 174997
rect 379470 174994 380052 174996
rect 376845 174992 380052 174994
rect 376845 174936 376850 174992
rect 376906 174936 380052 174992
rect 216673 174934 219450 174936
rect 376845 174934 379530 174936
rect 216673 174931 216739 174934
rect 376845 174931 376911 174934
rect 57881 173362 57947 173365
rect 59494 173362 60032 173364
rect 57881 173360 60032 173362
rect 57881 173304 57886 173360
rect 57942 173304 60032 173360
rect 216673 173362 216739 173365
rect 219390 173362 220064 173364
rect 216673 173360 220064 173362
rect 216673 173304 216678 173360
rect 216734 173304 220064 173360
rect 376845 173362 376911 173365
rect 379470 173362 380052 173364
rect 376845 173360 380052 173362
rect 376845 173304 376850 173360
rect 376906 173304 380052 173360
rect 57881 173302 59554 173304
rect 216673 173302 219450 173304
rect 376845 173302 379530 173304
rect 57881 173299 57947 173302
rect 216673 173299 216739 173302
rect 376845 173299 376911 173302
rect 57462 173028 57468 173092
rect 57532 173090 57538 173092
rect 217041 173090 217107 173093
rect 219390 173090 220064 173092
rect 57532 173030 60062 173090
rect 217041 173088 220064 173090
rect 217041 173032 217046 173088
rect 217102 173032 220064 173088
rect 376753 173090 376819 173093
rect 379470 173090 380052 173092
rect 376753 173088 380052 173090
rect 376753 173032 376758 173088
rect 376814 173032 380052 173088
rect 217041 173030 219450 173032
rect 376753 173030 379530 173032
rect 57532 173028 57538 173030
rect 217041 173027 217107 173030
rect 376753 173027 376819 173030
rect 583520 165732 584960 165972
rect 96061 164796 96127 164797
rect 140865 164796 140931 164797
rect 258441 164796 258507 164797
rect 96061 164792 96108 164796
rect 96172 164794 96178 164796
rect 96061 164736 96066 164792
rect 96061 164732 96108 164736
rect 96172 164734 96218 164794
rect 140865 164792 140926 164796
rect 140865 164736 140870 164792
rect 96172 164732 96178 164734
rect 140865 164732 140926 164736
rect 140990 164794 140996 164796
rect 140990 164734 141022 164794
rect 258441 164792 258494 164796
rect 258558 164794 258564 164796
rect 282177 164794 282243 164797
rect 425973 164796 426039 164797
rect 434345 164796 434411 164797
rect 450997 164796 451063 164797
rect 295888 164794 295894 164796
rect 258441 164736 258446 164792
rect 140990 164732 140996 164734
rect 258441 164732 258494 164736
rect 258558 164734 258598 164794
rect 282177 164792 295894 164794
rect 282177 164736 282182 164792
rect 282238 164736 295894 164792
rect 282177 164734 295894 164736
rect 258558 164732 258564 164734
rect 96061 164731 96127 164732
rect 140865 164731 140931 164732
rect 258441 164731 258507 164732
rect 282177 164731 282243 164734
rect 295888 164732 295894 164734
rect 295958 164732 295964 164796
rect 425968 164794 425974 164796
rect 425882 164734 425974 164794
rect 425968 164732 425974 164734
rect 426038 164732 426044 164796
rect 434345 164792 434406 164796
rect 434345 164736 434350 164792
rect 434345 164732 434406 164736
rect 434470 164794 434476 164796
rect 450992 164794 450998 164796
rect 434470 164734 434502 164794
rect 450906 164734 450998 164794
rect 434470 164732 434476 164734
rect 450992 164732 450998 164734
rect 451062 164732 451068 164796
rect 425973 164731 426039 164732
rect 434345 164731 434411 164732
rect 450997 164731 451063 164732
rect 103513 164660 103579 164661
rect 105905 164660 105971 164661
rect 117037 164660 117103 164661
rect 103513 164656 103526 164660
rect 103590 164658 103596 164660
rect 103513 164600 103518 164656
rect 103513 164596 103526 164600
rect 103590 164598 103670 164658
rect 105905 164656 105974 164660
rect 105905 164600 105910 164656
rect 105966 164600 105974 164656
rect 103590 164596 103596 164598
rect 105905 164596 105974 164600
rect 106038 164658 106044 164660
rect 116984 164658 116990 164660
rect 106038 164598 106062 164658
rect 116946 164598 116990 164658
rect 117054 164656 117103 164660
rect 117098 164600 117103 164656
rect 106038 164596 106044 164598
rect 116984 164596 116990 164598
rect 117054 164596 117103 164600
rect 103513 164595 103579 164596
rect 105905 164595 105971 164596
rect 117037 164595 117103 164596
rect 153377 164660 153443 164661
rect 163313 164660 163379 164661
rect 261017 164660 261083 164661
rect 153377 164656 153438 164660
rect 153377 164600 153382 164656
rect 153377 164596 153438 164600
rect 153502 164658 153508 164660
rect 153502 164598 153534 164658
rect 163313 164656 163366 164660
rect 163430 164658 163436 164660
rect 163313 164600 163318 164656
rect 153502 164596 153508 164598
rect 163313 164596 163366 164600
rect 163430 164598 163470 164658
rect 261017 164656 261078 164660
rect 261017 164600 261022 164656
rect 163430 164596 163436 164598
rect 261017 164596 261078 164600
rect 261142 164658 261148 164660
rect 261142 164598 261174 164658
rect 261142 164596 261148 164598
rect 275760 164596 275766 164660
rect 275830 164658 275836 164660
rect 276105 164658 276171 164661
rect 305913 164660 305979 164661
rect 318425 164660 318491 164661
rect 423489 164660 423555 164661
rect 436921 164660 436987 164661
rect 438025 164660 438091 164661
rect 480897 164660 480963 164661
rect 275830 164656 276171 164658
rect 275830 164600 276110 164656
rect 276166 164600 276171 164656
rect 275830 164598 276171 164600
rect 275830 164596 275836 164598
rect 153377 164595 153443 164596
rect 163313 164595 163379 164596
rect 261017 164595 261083 164596
rect 276105 164595 276171 164598
rect 288272 164596 288278 164660
rect 288342 164596 288348 164660
rect 305913 164656 305958 164660
rect 306022 164658 306028 164660
rect 305913 164600 305918 164656
rect 305913 164596 305958 164600
rect 306022 164598 306070 164658
rect 318425 164656 318470 164660
rect 318534 164658 318540 164660
rect 318425 164600 318430 164656
rect 306022 164596 306028 164598
rect 318425 164596 318470 164600
rect 318534 164598 318582 164658
rect 423489 164656 423526 164660
rect 423590 164658 423596 164660
rect 423489 164600 423494 164656
rect 318534 164596 318540 164598
rect 423489 164596 423526 164600
rect 423590 164598 423646 164658
rect 436921 164656 436990 164660
rect 436921 164600 436926 164656
rect 436982 164600 436990 164656
rect 423590 164596 423596 164598
rect 436921 164596 436990 164600
rect 437054 164658 437060 164660
rect 437054 164598 437078 164658
rect 438025 164656 438078 164660
rect 438142 164658 438148 164660
rect 438025 164600 438030 164656
rect 437054 164596 437060 164598
rect 438025 164596 438078 164600
rect 438142 164598 438182 164658
rect 480897 164656 480918 164660
rect 480982 164658 480988 164660
rect 480897 164600 480902 164656
rect 438142 164596 438148 164598
rect 480897 164596 480918 164600
rect 480982 164598 481054 164658
rect 480982 164596 480988 164598
rect 249149 164522 249215 164525
rect 262857 164522 262923 164525
rect 249149 164520 262923 164522
rect 249149 164464 249154 164520
rect 249210 164464 262862 164520
rect 262918 164464 262923 164520
rect 249149 164462 262923 164464
rect 249149 164459 249215 164462
rect 262857 164459 262923 164462
rect 55438 164324 55444 164388
rect 55508 164386 55514 164388
rect 138422 164386 138428 164388
rect 55508 164326 138428 164386
rect 55508 164324 55514 164326
rect 138422 164324 138428 164326
rect 138492 164324 138498 164388
rect 213126 164324 213132 164388
rect 213196 164386 213202 164388
rect 288280 164386 288340 164596
rect 305913 164595 305979 164596
rect 318425 164595 318491 164596
rect 423489 164595 423555 164596
rect 436921 164595 436987 164596
rect 438025 164595 438091 164596
rect 480897 164595 480963 164596
rect 213196 164326 288340 164386
rect 213196 164324 213202 164326
rect 98453 164252 98519 164253
rect 101029 164252 101095 164253
rect 108205 164252 108271 164253
rect 145925 164252 145991 164253
rect 148501 164252 148567 164253
rect 150893 164252 150959 164253
rect 98453 164248 98500 164252
rect 98564 164250 98570 164252
rect 98453 164192 98458 164248
rect 98453 164188 98500 164192
rect 98564 164190 98610 164250
rect 101029 164248 101076 164252
rect 101140 164250 101146 164252
rect 101029 164192 101034 164248
rect 98564 164188 98570 164190
rect 101029 164188 101076 164192
rect 101140 164190 101186 164250
rect 108205 164248 108252 164252
rect 108316 164250 108322 164252
rect 108205 164192 108210 164248
rect 101140 164188 101146 164190
rect 108205 164188 108252 164192
rect 108316 164190 108362 164250
rect 145925 164248 145972 164252
rect 146036 164250 146042 164252
rect 145925 164192 145930 164248
rect 108316 164188 108322 164190
rect 145925 164188 145972 164192
rect 146036 164190 146082 164250
rect 148501 164248 148548 164252
rect 148612 164250 148618 164252
rect 148501 164192 148506 164248
rect 146036 164188 146042 164190
rect 148501 164188 148548 164192
rect 148612 164190 148658 164250
rect 150893 164248 150940 164252
rect 151004 164250 151010 164252
rect 150893 164192 150898 164248
rect 148612 164188 148618 164190
rect 150893 164188 150940 164192
rect 151004 164190 151050 164250
rect 151004 164188 151010 164190
rect 210366 164188 210372 164252
rect 210436 164250 210442 164252
rect 249149 164250 249215 164253
rect 210436 164248 249215 164250
rect 210436 164192 249154 164248
rect 249210 164192 249215 164248
rect 210436 164190 249215 164192
rect 210436 164188 210442 164190
rect 98453 164187 98519 164188
rect 101029 164187 101095 164188
rect 108205 164187 108271 164188
rect 145925 164187 145991 164188
rect 148501 164187 148567 164188
rect 150893 164187 150959 164188
rect 249149 164187 249215 164190
rect 262857 164250 262923 164253
rect 282177 164250 282243 164253
rect 262857 164248 282243 164250
rect 262857 164192 262862 164248
rect 262918 164192 282182 164248
rect 282238 164192 282243 164248
rect 262857 164190 282243 164192
rect 262857 164187 262923 164190
rect 282177 164187 282243 164190
rect 298461 164252 298527 164253
rect 300853 164252 300919 164253
rect 298461 164248 298508 164252
rect 298572 164250 298578 164252
rect 298461 164192 298466 164248
rect 298461 164188 298508 164192
rect 298572 164190 298618 164250
rect 300853 164248 300900 164252
rect 300964 164250 300970 164252
rect 300853 164192 300858 164248
rect 298572 164188 298578 164190
rect 300853 164188 300900 164192
rect 300964 164190 301010 164250
rect 300964 164188 300970 164190
rect 377806 164188 377812 164252
rect 377876 164250 377882 164252
rect 378409 164250 378475 164253
rect 377876 164248 378475 164250
rect 377876 164192 378414 164248
rect 378470 164192 378475 164248
rect 377876 164190 378475 164192
rect 377876 164188 377882 164190
rect 298461 164187 298527 164188
rect 300853 164187 300919 164188
rect 378409 164187 378475 164190
rect 416037 164252 416103 164253
rect 421005 164252 421071 164253
rect 428181 164252 428247 164253
rect 430941 164252 431007 164253
rect 473445 164252 473511 164253
rect 475837 164252 475903 164253
rect 478413 164252 478479 164253
rect 416037 164248 416084 164252
rect 416148 164250 416154 164252
rect 416037 164192 416042 164248
rect 416037 164188 416084 164192
rect 416148 164190 416194 164250
rect 421005 164248 421052 164252
rect 421116 164250 421122 164252
rect 421005 164192 421010 164248
rect 416148 164188 416154 164190
rect 421005 164188 421052 164192
rect 421116 164190 421162 164250
rect 428181 164248 428228 164252
rect 428292 164250 428298 164252
rect 428181 164192 428186 164248
rect 421116 164188 421122 164190
rect 428181 164188 428228 164192
rect 428292 164190 428338 164250
rect 430941 164248 430988 164252
rect 431052 164250 431058 164252
rect 430941 164192 430946 164248
rect 428292 164188 428298 164190
rect 430941 164188 430988 164192
rect 431052 164190 431098 164250
rect 473445 164248 473492 164252
rect 473556 164250 473562 164252
rect 473445 164192 473450 164248
rect 431052 164188 431058 164190
rect 473445 164188 473492 164192
rect 473556 164190 473602 164250
rect 475837 164248 475884 164252
rect 475948 164250 475954 164252
rect 475837 164192 475842 164248
rect 473556 164188 473562 164190
rect 475837 164188 475884 164192
rect 475948 164190 475994 164250
rect 478413 164248 478460 164252
rect 478524 164250 478530 164252
rect 478413 164192 478418 164248
rect 475948 164188 475954 164190
rect 478413 164188 478460 164192
rect 478524 164190 478570 164250
rect 478524 164188 478530 164190
rect 416037 164187 416103 164188
rect 421005 164187 421071 164188
rect 428181 164187 428247 164188
rect 430941 164187 431007 164188
rect 473445 164187 473511 164188
rect 475837 164187 475903 164188
rect 478413 164187 478479 164188
rect 57646 164052 57652 164116
rect 57716 164114 57722 164116
rect 143574 164114 143580 164116
rect 57716 164054 143580 164114
rect 57716 164052 57722 164054
rect 143574 164052 143580 164054
rect 143644 164052 143650 164116
rect 202454 164052 202460 164116
rect 202524 164114 202530 164116
rect 323342 164114 323348 164116
rect 202524 164054 323348 164114
rect 202524 164052 202530 164054
rect 323342 164052 323348 164054
rect 323412 164052 323418 164116
rect 365345 164114 365411 164117
rect 485998 164114 486004 164116
rect 365345 164112 486004 164114
rect 365345 164056 365350 164112
rect 365406 164056 486004 164112
rect 365345 164054 486004 164056
rect 365345 164051 365411 164054
rect 485998 164052 486004 164054
rect 486068 164052 486074 164116
rect 203006 163916 203012 163980
rect 203076 163978 203082 163980
rect 311014 163978 311020 163980
rect 203076 163918 311020 163978
rect 203076 163916 203082 163918
rect 311014 163916 311020 163918
rect 311084 163916 311090 163980
rect 370773 163978 370839 163981
rect 483422 163978 483428 163980
rect 370773 163976 483428 163978
rect 370773 163920 370778 163976
rect 370834 163920 483428 163976
rect 370773 163918 483428 163920
rect 370773 163915 370839 163918
rect 483422 163916 483428 163918
rect 483492 163916 483498 163980
rect 206318 163780 206324 163844
rect 206388 163842 206394 163844
rect 313406 163842 313412 163844
rect 206388 163782 313412 163842
rect 206388 163780 206394 163782
rect 313406 163780 313412 163782
rect 313476 163780 313482 163844
rect 470358 163780 470364 163844
rect 470428 163842 470434 163844
rect 470593 163842 470659 163845
rect 470428 163840 470659 163842
rect 470428 163784 470598 163840
rect 470654 163784 470659 163840
rect 470428 163782 470659 163784
rect 470428 163780 470434 163782
rect 470593 163779 470659 163782
rect 207974 163644 207980 163708
rect 208044 163706 208050 163708
rect 315798 163706 315804 163708
rect 208044 163646 315804 163706
rect 208044 163644 208050 163646
rect 315798 163644 315804 163646
rect 315868 163644 315874 163708
rect 198038 163508 198044 163572
rect 198108 163570 198114 163572
rect 290958 163570 290964 163572
rect 198108 163510 290964 163570
rect 198108 163508 198114 163510
rect 290958 163508 290964 163510
rect 291028 163508 291034 163572
rect 196566 163372 196572 163436
rect 196636 163434 196642 163436
rect 270902 163434 270908 163436
rect 196636 163374 270908 163434
rect 196636 163372 196642 163374
rect 270902 163372 270908 163374
rect 270972 163372 270978 163436
rect 99373 163164 99439 163165
rect 113541 163164 113607 163165
rect 128353 163164 128419 163165
rect 235993 163164 236059 163165
rect 85430 163100 85436 163164
rect 85500 163100 85506 163164
rect 95918 163100 95924 163164
rect 95988 163100 95994 163164
rect 99373 163160 99420 163164
rect 99484 163162 99490 163164
rect 99373 163104 99378 163160
rect 99373 163100 99420 163104
rect 99484 163102 99530 163162
rect 113541 163160 113588 163164
rect 113652 163162 113658 163164
rect 128302 163162 128308 163164
rect 113541 163104 113546 163160
rect 99484 163100 99490 163102
rect 113541 163100 113588 163104
rect 113652 163102 113698 163162
rect 128262 163102 128308 163162
rect 128372 163160 128419 163164
rect 235942 163162 235948 163164
rect 128414 163104 128419 163160
rect 113652 163100 113658 163102
rect 128302 163100 128308 163102
rect 128372 163100 128419 163104
rect 235902 163102 235948 163162
rect 236012 163160 236059 163164
rect 236054 163104 236059 163160
rect 235942 163100 235948 163102
rect 236012 163100 236059 163104
rect 261702 163100 261708 163164
rect 261772 163100 261778 163164
rect 264973 163162 265039 163165
rect 265198 163162 265204 163164
rect 264973 163160 265204 163162
rect 264973 163104 264978 163160
rect 265034 163104 265204 163160
rect 264973 163102 265204 163104
rect -960 162740 480 162980
rect 54702 162692 54708 162756
rect 54772 162754 54778 162756
rect 55121 162754 55187 162757
rect 54772 162752 55187 162754
rect 54772 162696 55126 162752
rect 55182 162696 55187 162752
rect 54772 162694 55187 162696
rect 54772 162692 54778 162694
rect 55121 162691 55187 162694
rect 75913 162754 75979 162757
rect 76046 162754 76052 162756
rect 75913 162752 76052 162754
rect 75913 162696 75918 162752
rect 75974 162696 76052 162752
rect 75913 162694 76052 162696
rect 75913 162691 75979 162694
rect 76046 162692 76052 162694
rect 76116 162692 76122 162756
rect 77293 162754 77359 162757
rect 78254 162754 78260 162756
rect 77293 162752 78260 162754
rect 77293 162696 77298 162752
rect 77354 162696 78260 162752
rect 77293 162694 78260 162696
rect 77293 162691 77359 162694
rect 78254 162692 78260 162694
rect 78324 162692 78330 162756
rect 78673 162754 78739 162757
rect 79542 162754 79548 162756
rect 78673 162752 79548 162754
rect 78673 162696 78678 162752
rect 78734 162696 79548 162752
rect 78673 162694 79548 162696
rect 78673 162691 78739 162694
rect 79542 162692 79548 162694
rect 79612 162692 79618 162756
rect 80053 162754 80119 162757
rect 80462 162754 80468 162756
rect 80053 162752 80468 162754
rect 80053 162696 80058 162752
rect 80114 162696 80468 162752
rect 80053 162694 80468 162696
rect 80053 162691 80119 162694
rect 80462 162692 80468 162694
rect 80532 162692 80538 162756
rect 81433 162754 81499 162757
rect 81934 162754 81940 162756
rect 81433 162752 81940 162754
rect 81433 162696 81438 162752
rect 81494 162696 81940 162752
rect 81433 162694 81940 162696
rect 81433 162691 81499 162694
rect 81934 162692 81940 162694
rect 82004 162692 82010 162756
rect 82813 162754 82879 162757
rect 83038 162754 83044 162756
rect 82813 162752 83044 162754
rect 82813 162696 82818 162752
rect 82874 162696 83044 162752
rect 82813 162694 83044 162696
rect 82813 162691 82879 162694
rect 83038 162692 83044 162694
rect 83108 162692 83114 162756
rect 84193 162754 84259 162757
rect 85438 162754 85498 163100
rect 84193 162752 85498 162754
rect 84193 162696 84198 162752
rect 84254 162696 85498 162752
rect 84193 162694 85498 162696
rect 85573 162754 85639 162757
rect 86534 162754 86540 162756
rect 85573 162752 86540 162754
rect 85573 162696 85578 162752
rect 85634 162696 86540 162752
rect 85573 162694 86540 162696
rect 84193 162691 84259 162694
rect 85573 162691 85639 162694
rect 86534 162692 86540 162694
rect 86604 162692 86610 162756
rect 86953 162754 87019 162757
rect 87638 162754 87644 162756
rect 86953 162752 87644 162754
rect 86953 162696 86958 162752
rect 87014 162696 87644 162752
rect 86953 162694 87644 162696
rect 86953 162691 87019 162694
rect 87638 162692 87644 162694
rect 87708 162692 87714 162756
rect 88425 162754 88491 162757
rect 88742 162754 88748 162756
rect 88425 162752 88748 162754
rect 88425 162696 88430 162752
rect 88486 162696 88748 162752
rect 88425 162694 88748 162696
rect 88425 162691 88491 162694
rect 88742 162692 88748 162694
rect 88812 162692 88818 162756
rect 89805 162754 89871 162757
rect 90725 162756 90791 162757
rect 90030 162754 90036 162756
rect 89805 162752 90036 162754
rect 89805 162696 89810 162752
rect 89866 162696 90036 162752
rect 89805 162694 90036 162696
rect 89805 162691 89871 162694
rect 90030 162692 90036 162694
rect 90100 162692 90106 162756
rect 90725 162752 90772 162756
rect 90836 162754 90842 162756
rect 91185 162754 91251 162757
rect 91318 162754 91324 162756
rect 90725 162696 90730 162752
rect 90725 162692 90772 162696
rect 90836 162694 90882 162754
rect 91185 162752 91324 162754
rect 91185 162696 91190 162752
rect 91246 162696 91324 162752
rect 91185 162694 91324 162696
rect 90836 162692 90842 162694
rect 90725 162691 90791 162692
rect 91185 162691 91251 162694
rect 91318 162692 91324 162694
rect 91388 162692 91394 162756
rect 92473 162754 92539 162757
rect 93669 162756 93735 162757
rect 93342 162754 93348 162756
rect 92473 162752 93348 162754
rect 92473 162696 92478 162752
rect 92534 162696 93348 162752
rect 92473 162694 93348 162696
rect 92473 162691 92539 162694
rect 93342 162692 93348 162694
rect 93412 162692 93418 162756
rect 93669 162754 93716 162756
rect 93624 162752 93716 162754
rect 93624 162696 93674 162752
rect 93624 162694 93716 162696
rect 93669 162692 93716 162694
rect 93780 162692 93786 162756
rect 93853 162754 93919 162757
rect 94446 162754 94452 162756
rect 93853 162752 94452 162754
rect 93853 162696 93858 162752
rect 93914 162696 94452 162752
rect 93853 162694 94452 162696
rect 93669 162691 93735 162692
rect 93853 162691 93919 162694
rect 94446 162692 94452 162694
rect 94516 162692 94522 162756
rect 95233 162754 95299 162757
rect 95926 162754 95986 163100
rect 99373 163099 99439 163100
rect 113541 163099 113607 163100
rect 128353 163099 128419 163100
rect 235993 163099 236059 163100
rect 95233 162752 95986 162754
rect 95233 162696 95238 162752
rect 95294 162696 95986 162752
rect 95233 162694 95986 162696
rect 96889 162754 96955 162757
rect 97022 162754 97028 162756
rect 96889 162752 97028 162754
rect 96889 162696 96894 162752
rect 96950 162696 97028 162752
rect 96889 162694 97028 162696
rect 95233 162691 95299 162694
rect 96889 162691 96955 162694
rect 97022 162692 97028 162694
rect 97092 162692 97098 162756
rect 97993 162754 98059 162757
rect 100753 162756 100819 162757
rect 98126 162754 98132 162756
rect 97993 162752 98132 162754
rect 97993 162696 97998 162752
rect 98054 162696 98132 162752
rect 97993 162694 98132 162696
rect 97993 162691 98059 162694
rect 98126 162692 98132 162694
rect 98196 162692 98202 162756
rect 100702 162754 100708 162756
rect 100662 162694 100708 162754
rect 100772 162752 100819 162756
rect 100814 162696 100819 162752
rect 100702 162692 100708 162694
rect 100772 162692 100819 162696
rect 100753 162691 100819 162692
rect 102133 162754 102199 162757
rect 102726 162754 102732 162756
rect 102133 162752 102732 162754
rect 102133 162696 102138 162752
rect 102194 162696 102732 162752
rect 102133 162694 102732 162696
rect 102133 162691 102199 162694
rect 102726 162692 102732 162694
rect 102796 162692 102802 162756
rect 103513 162754 103579 162757
rect 103830 162754 103836 162756
rect 103513 162752 103836 162754
rect 103513 162696 103518 162752
rect 103574 162696 103836 162752
rect 103513 162694 103836 162696
rect 103513 162691 103579 162694
rect 103830 162692 103836 162694
rect 103900 162692 103906 162756
rect 104893 162754 104959 162757
rect 105302 162754 105308 162756
rect 104893 162752 105308 162754
rect 104893 162696 104898 162752
rect 104954 162696 105308 162752
rect 104893 162694 105308 162696
rect 104893 162691 104959 162694
rect 105302 162692 105308 162694
rect 105372 162692 105378 162756
rect 106273 162754 106339 162757
rect 106406 162754 106412 162756
rect 106273 162752 106412 162754
rect 106273 162696 106278 162752
rect 106334 162696 106412 162752
rect 106273 162694 106412 162696
rect 106273 162691 106339 162694
rect 106406 162692 106412 162694
rect 106476 162692 106482 162756
rect 107653 162754 107719 162757
rect 108614 162754 108620 162756
rect 107653 162752 108620 162754
rect 107653 162696 107658 162752
rect 107714 162696 108620 162752
rect 107653 162694 108620 162696
rect 107653 162691 107719 162694
rect 108614 162692 108620 162694
rect 108684 162692 108690 162756
rect 109033 162754 109099 162757
rect 109534 162754 109540 162756
rect 109033 162752 109540 162754
rect 109033 162696 109038 162752
rect 109094 162696 109540 162752
rect 109033 162694 109540 162696
rect 109033 162691 109099 162694
rect 109534 162692 109540 162694
rect 109604 162692 109610 162756
rect 110413 162754 110479 162757
rect 111190 162754 111196 162756
rect 110413 162752 111196 162754
rect 110413 162696 110418 162752
rect 110474 162696 111196 162752
rect 110413 162694 111196 162696
rect 110413 162691 110479 162694
rect 111190 162692 111196 162694
rect 111260 162692 111266 162756
rect 111793 162754 111859 162757
rect 112110 162754 112116 162756
rect 111793 162752 112116 162754
rect 111793 162696 111798 162752
rect 111854 162696 112116 162752
rect 111793 162694 112116 162696
rect 111793 162691 111859 162694
rect 112110 162692 112116 162694
rect 112180 162692 112186 162756
rect 113214 162692 113220 162756
rect 113284 162754 113290 162756
rect 114461 162754 114527 162757
rect 113284 162752 114527 162754
rect 113284 162696 114466 162752
rect 114522 162696 114527 162752
rect 113284 162694 114527 162696
rect 113284 162692 113290 162694
rect 114461 162691 114527 162694
rect 114737 162754 114803 162757
rect 115933 162756 115999 162757
rect 115790 162754 115796 162756
rect 114737 162752 115796 162754
rect 114737 162696 114742 162752
rect 114798 162696 115796 162752
rect 114737 162694 115796 162696
rect 114737 162691 114803 162694
rect 115790 162692 115796 162694
rect 115860 162692 115866 162756
rect 115933 162752 115980 162756
rect 116044 162754 116050 162756
rect 117313 162754 117379 162757
rect 118325 162756 118391 162757
rect 117998 162754 118004 162756
rect 115933 162696 115938 162752
rect 115933 162692 115980 162696
rect 116044 162694 116090 162754
rect 117313 162752 118004 162754
rect 117313 162696 117318 162752
rect 117374 162696 118004 162752
rect 117313 162694 118004 162696
rect 116044 162692 116050 162694
rect 115933 162691 115999 162692
rect 117313 162691 117379 162694
rect 117998 162692 118004 162694
rect 118068 162692 118074 162756
rect 118325 162752 118372 162756
rect 118436 162754 118442 162756
rect 118693 162754 118759 162757
rect 120717 162756 120783 162757
rect 119102 162754 119108 162756
rect 118325 162696 118330 162752
rect 118325 162692 118372 162696
rect 118436 162694 118482 162754
rect 118693 162752 119108 162754
rect 118693 162696 118698 162752
rect 118754 162696 119108 162752
rect 118693 162694 119108 162696
rect 118436 162692 118442 162694
rect 118325 162691 118391 162692
rect 118693 162691 118759 162694
rect 119102 162692 119108 162694
rect 119172 162692 119178 162756
rect 120717 162752 120764 162756
rect 120828 162754 120834 162756
rect 120717 162696 120722 162752
rect 120717 162692 120764 162696
rect 120828 162694 120874 162754
rect 120828 162692 120834 162694
rect 122598 162692 122604 162756
rect 122668 162754 122674 162756
rect 122833 162754 122899 162757
rect 122668 162752 122899 162754
rect 122668 162696 122838 162752
rect 122894 162696 122899 162752
rect 122668 162694 122899 162696
rect 122668 162692 122674 162694
rect 120717 162691 120783 162692
rect 122833 162691 122899 162694
rect 125869 162756 125935 162757
rect 130837 162756 130903 162757
rect 133413 162756 133479 162757
rect 183461 162756 183527 162757
rect 125869 162752 125916 162756
rect 125980 162754 125986 162756
rect 125869 162696 125874 162752
rect 125869 162692 125916 162696
rect 125980 162694 126026 162754
rect 130837 162752 130884 162756
rect 130948 162754 130954 162756
rect 130837 162696 130842 162752
rect 125980 162692 125986 162694
rect 130837 162692 130884 162696
rect 130948 162694 130994 162754
rect 133413 162752 133460 162756
rect 133524 162754 133530 162756
rect 133413 162696 133418 162752
rect 130948 162692 130954 162694
rect 133413 162692 133460 162696
rect 133524 162694 133570 162754
rect 183461 162752 183508 162756
rect 183572 162754 183578 162756
rect 236085 162754 236151 162757
rect 237046 162754 237052 162756
rect 183461 162696 183466 162752
rect 133524 162692 133530 162694
rect 183461 162692 183508 162696
rect 183572 162694 183618 162754
rect 236085 162752 237052 162754
rect 236085 162696 236090 162752
rect 236146 162696 237052 162752
rect 236085 162694 237052 162696
rect 183572 162692 183578 162694
rect 125869 162691 125935 162692
rect 130837 162691 130903 162692
rect 133413 162691 133479 162692
rect 183461 162691 183527 162692
rect 236085 162691 236151 162694
rect 237046 162692 237052 162694
rect 237116 162692 237122 162756
rect 237373 162754 237439 162757
rect 238150 162754 238156 162756
rect 237373 162752 238156 162754
rect 237373 162696 237378 162752
rect 237434 162696 238156 162752
rect 237373 162694 238156 162696
rect 237373 162691 237439 162694
rect 238150 162692 238156 162694
rect 238220 162692 238226 162756
rect 240133 162754 240199 162757
rect 240542 162754 240548 162756
rect 240133 162752 240548 162754
rect 240133 162696 240138 162752
rect 240194 162696 240548 162752
rect 240133 162694 240548 162696
rect 240133 162691 240199 162694
rect 240542 162692 240548 162694
rect 240612 162692 240618 162756
rect 241513 162754 241579 162757
rect 242893 162756 242959 162757
rect 244273 162756 244339 162757
rect 241646 162754 241652 162756
rect 241513 162752 241652 162754
rect 241513 162696 241518 162752
rect 241574 162696 241652 162752
rect 241513 162694 241652 162696
rect 241513 162691 241579 162694
rect 241646 162692 241652 162694
rect 241716 162692 241722 162756
rect 242893 162752 242940 162756
rect 243004 162754 243010 162756
rect 244222 162754 244228 162756
rect 242893 162696 242898 162752
rect 242893 162692 242940 162696
rect 243004 162694 243050 162754
rect 244182 162694 244228 162754
rect 244292 162752 244339 162756
rect 244334 162696 244339 162752
rect 243004 162692 243010 162694
rect 244222 162692 244228 162694
rect 244292 162692 244339 162696
rect 242893 162691 242959 162692
rect 244273 162691 244339 162692
rect 245653 162754 245719 162757
rect 246430 162754 246436 162756
rect 245653 162752 246436 162754
rect 245653 162696 245658 162752
rect 245714 162696 246436 162752
rect 245653 162694 246436 162696
rect 245653 162691 245719 162694
rect 246430 162692 246436 162694
rect 246500 162692 246506 162756
rect 247125 162754 247191 162757
rect 247718 162754 247724 162756
rect 247125 162752 247724 162754
rect 247125 162696 247130 162752
rect 247186 162696 247724 162752
rect 247125 162694 247724 162696
rect 247125 162691 247191 162694
rect 247718 162692 247724 162694
rect 247788 162692 247794 162756
rect 247861 162754 247927 162757
rect 248270 162754 248276 162756
rect 247861 162752 248276 162754
rect 247861 162696 247866 162752
rect 247922 162696 248276 162752
rect 247861 162694 248276 162696
rect 247861 162691 247927 162694
rect 248270 162692 248276 162694
rect 248340 162692 248346 162756
rect 248413 162754 248479 162757
rect 248638 162754 248644 162756
rect 248413 162752 248644 162754
rect 248413 162696 248418 162752
rect 248474 162696 248644 162752
rect 248413 162694 248644 162696
rect 248413 162691 248479 162694
rect 248638 162692 248644 162694
rect 248708 162692 248714 162756
rect 249793 162754 249859 162757
rect 251265 162756 251331 162757
rect 250110 162754 250116 162756
rect 249793 162752 250116 162754
rect 249793 162696 249798 162752
rect 249854 162696 250116 162752
rect 249793 162694 250116 162696
rect 249793 162691 249859 162694
rect 250110 162692 250116 162694
rect 250180 162692 250186 162756
rect 251214 162754 251220 162756
rect 251174 162694 251220 162754
rect 251284 162752 251331 162756
rect 251326 162696 251331 162752
rect 251214 162692 251220 162694
rect 251284 162692 251331 162696
rect 251265 162691 251331 162692
rect 252553 162754 252619 162757
rect 253422 162754 253428 162756
rect 252553 162752 253428 162754
rect 252553 162696 252558 162752
rect 252614 162696 253428 162752
rect 252553 162694 253428 162696
rect 252553 162691 252619 162694
rect 253422 162692 253428 162694
rect 253492 162692 253498 162756
rect 253933 162754 253999 162757
rect 254526 162754 254532 162756
rect 253933 162752 254532 162754
rect 253933 162696 253938 162752
rect 253994 162696 254532 162752
rect 253933 162694 254532 162696
rect 253933 162691 253999 162694
rect 254526 162692 254532 162694
rect 254596 162692 254602 162756
rect 255405 162754 255471 162757
rect 255957 162756 256023 162757
rect 255814 162754 255820 162756
rect 255405 162752 255820 162754
rect 255405 162696 255410 162752
rect 255466 162696 255820 162752
rect 255405 162694 255820 162696
rect 255405 162691 255471 162694
rect 255814 162692 255820 162694
rect 255884 162692 255890 162756
rect 255957 162752 256004 162756
rect 256068 162754 256074 162756
rect 256693 162754 256759 162757
rect 259545 162756 259611 162757
rect 256918 162754 256924 162756
rect 255957 162696 255962 162752
rect 255957 162692 256004 162696
rect 256068 162694 256114 162754
rect 256693 162752 256924 162754
rect 256693 162696 256698 162752
rect 256754 162696 256924 162752
rect 256693 162694 256924 162696
rect 256068 162692 256074 162694
rect 255957 162691 256023 162692
rect 256693 162691 256759 162694
rect 256918 162692 256924 162694
rect 256988 162692 256994 162756
rect 259494 162754 259500 162756
rect 259454 162694 259500 162754
rect 259564 162752 259611 162756
rect 259606 162696 259611 162752
rect 259494 162692 259500 162694
rect 259564 162692 259611 162696
rect 259545 162691 259611 162692
rect 260833 162754 260899 162757
rect 261710 162754 261770 163100
rect 264973 163099 265039 163102
rect 265198 163100 265204 163102
rect 265268 163100 265274 163164
rect 272190 163100 272196 163164
rect 272260 163100 272266 163164
rect 325918 163100 325924 163164
rect 325988 163100 325994 163164
rect 398230 163100 398236 163164
rect 398300 163100 398306 163164
rect 401593 163162 401659 163165
rect 455781 163164 455847 163165
rect 401726 163162 401732 163164
rect 401593 163160 401732 163162
rect 401593 163104 401598 163160
rect 401654 163104 401732 163160
rect 401593 163102 401732 163104
rect 260833 162752 261770 162754
rect 260833 162696 260838 162752
rect 260894 162696 261770 162752
rect 260833 162694 261770 162696
rect 262213 162754 262279 162757
rect 262806 162754 262812 162756
rect 262213 162752 262812 162754
rect 262213 162696 262218 162752
rect 262274 162696 262812 162752
rect 262213 162694 262812 162696
rect 260833 162691 260899 162694
rect 262213 162691 262279 162694
rect 262806 162692 262812 162694
rect 262876 162692 262882 162756
rect 263593 162754 263659 162757
rect 263910 162754 263916 162756
rect 263593 162752 263916 162754
rect 263593 162696 263598 162752
rect 263654 162696 263916 162752
rect 263593 162694 263916 162696
rect 263593 162691 263659 162694
rect 263910 162692 263916 162694
rect 263980 162692 263986 162756
rect 265433 162754 265499 162757
rect 266353 162756 266419 162757
rect 265934 162754 265940 162756
rect 265433 162752 265940 162754
rect 265433 162696 265438 162752
rect 265494 162696 265940 162752
rect 265433 162694 265940 162696
rect 265433 162691 265499 162694
rect 265934 162692 265940 162694
rect 266004 162692 266010 162756
rect 266302 162754 266308 162756
rect 266262 162694 266308 162754
rect 266372 162752 266419 162756
rect 267549 162756 267615 162757
rect 267549 162754 267596 162756
rect 266414 162696 266419 162752
rect 266302 162692 266308 162694
rect 266372 162692 266419 162696
rect 267504 162752 267596 162754
rect 267504 162696 267554 162752
rect 267504 162694 267596 162696
rect 266353 162691 266419 162692
rect 267549 162692 267596 162694
rect 267660 162692 267666 162756
rect 267733 162754 267799 162757
rect 268694 162754 268700 162756
rect 267733 162752 268700 162754
rect 267733 162696 267738 162752
rect 267794 162696 268700 162752
rect 267733 162694 268700 162696
rect 267549 162691 267615 162692
rect 267733 162691 267799 162694
rect 268694 162692 268700 162694
rect 268764 162692 268770 162756
rect 269113 162754 269179 162757
rect 269798 162754 269804 162756
rect 269113 162752 269804 162754
rect 269113 162696 269118 162752
rect 269174 162696 269804 162752
rect 269113 162694 269804 162696
rect 269113 162691 269179 162694
rect 269798 162692 269804 162694
rect 269868 162692 269874 162756
rect 270493 162754 270559 162757
rect 271086 162754 271092 162756
rect 270493 162752 271092 162754
rect 270493 162696 270498 162752
rect 270554 162696 271092 162752
rect 270493 162694 271092 162696
rect 270493 162691 270559 162694
rect 271086 162692 271092 162694
rect 271156 162692 271162 162756
rect 271873 162754 271939 162757
rect 272198 162754 272258 163100
rect 271873 162752 272258 162754
rect 271873 162696 271878 162752
rect 271934 162696 272258 162752
rect 271873 162694 272258 162696
rect 273253 162754 273319 162757
rect 274398 162754 274404 162756
rect 273253 162752 274404 162754
rect 273253 162696 273258 162752
rect 273314 162696 274404 162752
rect 273253 162694 274404 162696
rect 271873 162691 271939 162694
rect 273253 162691 273319 162694
rect 274398 162692 274404 162694
rect 274468 162692 274474 162756
rect 276013 162754 276079 162757
rect 278405 162756 278471 162757
rect 276974 162754 276980 162756
rect 276013 162752 276980 162754
rect 276013 162696 276018 162752
rect 276074 162696 276980 162752
rect 276013 162694 276980 162696
rect 276013 162691 276079 162694
rect 276974 162692 276980 162694
rect 277044 162692 277050 162756
rect 278405 162752 278452 162756
rect 278516 162754 278522 162756
rect 278405 162696 278410 162752
rect 278405 162692 278452 162696
rect 278516 162694 278562 162754
rect 278516 162692 278522 162694
rect 278998 162692 279004 162756
rect 279068 162754 279074 162756
rect 280061 162754 280127 162757
rect 279068 162752 280127 162754
rect 279068 162696 280066 162752
rect 280122 162696 280127 162752
rect 279068 162694 280127 162696
rect 279068 162692 279074 162694
rect 278405 162691 278471 162692
rect 280061 162691 280127 162694
rect 280797 162756 280863 162757
rect 283741 162756 283807 162757
rect 285949 162756 286015 162757
rect 293309 162756 293375 162757
rect 303429 162756 303495 162757
rect 308581 162756 308647 162757
rect 280797 162752 280844 162756
rect 280908 162754 280914 162756
rect 280797 162696 280802 162752
rect 280797 162692 280844 162696
rect 280908 162694 280954 162754
rect 283741 162752 283788 162756
rect 283852 162754 283858 162756
rect 283741 162696 283746 162752
rect 280908 162692 280914 162694
rect 283741 162692 283788 162696
rect 283852 162694 283898 162754
rect 285949 162752 285996 162756
rect 286060 162754 286066 162756
rect 285949 162696 285954 162752
rect 283852 162692 283858 162694
rect 285949 162692 285996 162696
rect 286060 162694 286106 162754
rect 293309 162752 293356 162756
rect 293420 162754 293426 162756
rect 293309 162696 293314 162752
rect 286060 162692 286066 162694
rect 293309 162692 293356 162696
rect 293420 162694 293466 162754
rect 303429 162752 303476 162756
rect 303540 162754 303546 162756
rect 303429 162696 303434 162752
rect 293420 162692 293426 162694
rect 303429 162692 303476 162696
rect 303540 162694 303586 162754
rect 308581 162752 308628 162756
rect 308692 162754 308698 162756
rect 325926 162754 325986 163100
rect 343449 162756 343515 162757
rect 396073 162756 396139 162757
rect 343398 162754 343404 162756
rect 308581 162696 308586 162752
rect 303540 162692 303546 162694
rect 308581 162692 308628 162696
rect 308692 162694 308738 162754
rect 315990 162694 325986 162754
rect 343358 162694 343404 162754
rect 343468 162752 343515 162756
rect 396022 162754 396028 162756
rect 343510 162696 343515 162752
rect 308692 162692 308698 162694
rect 280797 162691 280863 162692
rect 283741 162691 283807 162692
rect 285949 162691 286015 162692
rect 293309 162691 293375 162692
rect 303429 162691 303495 162692
rect 308581 162691 308647 162692
rect 49509 162618 49575 162621
rect 158478 162618 158484 162620
rect 49509 162616 158484 162618
rect 49509 162560 49514 162616
rect 49570 162560 158484 162616
rect 49509 162558 158484 162560
rect 49509 162555 49575 162558
rect 158478 162556 158484 162558
rect 158548 162556 158554 162620
rect 166022 162556 166028 162620
rect 166092 162618 166098 162620
rect 198774 162618 198780 162620
rect 166092 162558 198780 162618
rect 166092 162556 166098 162558
rect 198774 162556 198780 162558
rect 198844 162556 198850 162620
rect 214782 162556 214788 162620
rect 214852 162618 214858 162620
rect 259453 162618 259519 162621
rect 260598 162618 260604 162620
rect 214852 162558 258090 162618
rect 214852 162556 214858 162558
rect 53465 162482 53531 162485
rect 183185 162484 183251 162485
rect 155902 162482 155908 162484
rect 53465 162480 155908 162482
rect 53465 162424 53470 162480
rect 53526 162424 155908 162480
rect 53465 162422 155908 162424
rect 53465 162419 53531 162422
rect 155902 162420 155908 162422
rect 155972 162420 155978 162484
rect 183134 162482 183140 162484
rect 183094 162422 183140 162482
rect 183204 162480 183251 162484
rect 183246 162424 183251 162480
rect 183134 162420 183140 162422
rect 183204 162420 183251 162424
rect 203190 162420 203196 162484
rect 203260 162482 203266 162484
rect 251173 162482 251239 162485
rect 252318 162482 252324 162484
rect 203260 162422 251098 162482
rect 203260 162420 203266 162422
rect 183185 162419 183251 162420
rect 56317 162346 56383 162349
rect 136030 162346 136036 162348
rect 56317 162344 136036 162346
rect 56317 162288 56322 162344
rect 56378 162288 136036 162344
rect 56317 162286 136036 162288
rect 56317 162283 56383 162286
rect 136030 162284 136036 162286
rect 136100 162284 136106 162348
rect 214966 162284 214972 162348
rect 215036 162346 215042 162348
rect 250662 162346 250668 162348
rect 215036 162286 250668 162346
rect 215036 162284 215042 162286
rect 250662 162284 250668 162286
rect 250732 162284 250738 162348
rect 251038 162346 251098 162422
rect 251173 162480 252324 162482
rect 251173 162424 251178 162480
rect 251234 162424 252324 162480
rect 251173 162422 252324 162424
rect 251173 162419 251239 162422
rect 252318 162420 252324 162422
rect 252388 162420 252394 162484
rect 258030 162482 258090 162558
rect 259453 162616 260604 162618
rect 259453 162560 259458 162616
rect 259514 162560 260604 162616
rect 259453 162558 260604 162560
rect 259453 162555 259519 162558
rect 260598 162556 260604 162558
rect 260668 162556 260674 162620
rect 263542 162556 263548 162620
rect 263612 162618 263618 162620
rect 263685 162618 263751 162621
rect 263612 162616 263751 162618
rect 263612 162560 263690 162616
rect 263746 162560 263751 162616
rect 263612 162558 263751 162560
rect 263612 162556 263618 162558
rect 263685 162555 263751 162558
rect 268285 162620 268351 162621
rect 268285 162616 268332 162620
rect 268396 162618 268402 162620
rect 268285 162560 268290 162616
rect 268285 162556 268332 162560
rect 268396 162558 268442 162618
rect 268396 162556 268402 162558
rect 273294 162556 273300 162620
rect 273364 162618 273370 162620
rect 274541 162618 274607 162621
rect 273364 162616 274607 162618
rect 273364 162560 274546 162616
rect 274602 162560 274607 162616
rect 273364 162558 274607 162560
rect 273364 162556 273370 162558
rect 268285 162555 268351 162556
rect 274541 162555 274607 162558
rect 276238 162482 276244 162484
rect 258030 162422 276244 162482
rect 276238 162420 276244 162422
rect 276308 162420 276314 162484
rect 273437 162348 273503 162349
rect 253606 162346 253612 162348
rect 251038 162286 253612 162346
rect 253606 162284 253612 162286
rect 253676 162284 253682 162348
rect 273437 162344 273484 162348
rect 273548 162346 273554 162348
rect 273437 162288 273442 162344
rect 273437 162284 273484 162288
rect 273548 162286 273594 162346
rect 273548 162284 273554 162286
rect 273437 162283 273503 162284
rect 76005 162210 76071 162213
rect 88333 162212 88399 162213
rect 77150 162210 77156 162212
rect 76005 162208 77156 162210
rect 76005 162152 76010 162208
rect 76066 162152 77156 162208
rect 76005 162150 77156 162152
rect 76005 162147 76071 162150
rect 77150 162148 77156 162150
rect 77220 162148 77226 162212
rect 88333 162208 88380 162212
rect 88444 162210 88450 162212
rect 91093 162210 91159 162213
rect 91502 162210 91508 162212
rect 88333 162152 88338 162208
rect 88333 162148 88380 162152
rect 88444 162150 88490 162210
rect 91093 162208 91508 162210
rect 91093 162152 91098 162208
rect 91154 162152 91508 162208
rect 91093 162150 91508 162152
rect 88444 162148 88450 162150
rect 88333 162147 88399 162148
rect 91093 162147 91159 162150
rect 91502 162148 91508 162150
rect 91572 162148 91578 162212
rect 100845 162210 100911 162213
rect 101806 162210 101812 162212
rect 100845 162208 101812 162210
rect 100845 162152 100850 162208
rect 100906 162152 101812 162208
rect 100845 162150 101812 162152
rect 100845 162147 100911 162150
rect 101806 162148 101812 162150
rect 101876 162148 101882 162212
rect 106365 162210 106431 162213
rect 110965 162212 111031 162213
rect 107510 162210 107516 162212
rect 106365 162208 107516 162210
rect 106365 162152 106370 162208
rect 106426 162152 107516 162208
rect 106365 162150 107516 162152
rect 106365 162147 106431 162150
rect 107510 162148 107516 162150
rect 107580 162148 107586 162212
rect 110965 162208 111012 162212
rect 111076 162210 111082 162212
rect 244365 162210 244431 162213
rect 245326 162210 245332 162212
rect 110965 162152 110970 162208
rect 110965 162148 111012 162152
rect 111076 162150 111122 162210
rect 244365 162208 245332 162210
rect 244365 162152 244370 162208
rect 244426 162152 245332 162208
rect 244365 162150 245332 162152
rect 111076 162148 111082 162150
rect 110965 162147 111031 162148
rect 244365 162147 244431 162150
rect 245326 162148 245332 162150
rect 245396 162148 245402 162212
rect 258073 162210 258139 162213
rect 258390 162210 258396 162212
rect 258073 162208 258396 162210
rect 258073 162152 258078 162208
rect 258134 162152 258396 162208
rect 258073 162150 258396 162152
rect 258073 162147 258139 162150
rect 258390 162148 258396 162150
rect 258460 162148 258466 162212
rect 114502 162012 114508 162076
rect 114572 162074 114578 162076
rect 114645 162074 114711 162077
rect 196750 162074 196756 162076
rect 114572 162072 196756 162074
rect 114572 162016 114650 162072
rect 114706 162016 196756 162072
rect 114572 162014 196756 162016
rect 114572 162012 114578 162014
rect 114645 162011 114711 162014
rect 196750 162012 196756 162014
rect 196820 162012 196826 162076
rect 50613 161938 50679 161941
rect 160870 161938 160876 161940
rect 50613 161936 160876 161938
rect 50613 161880 50618 161936
rect 50674 161880 160876 161936
rect 50613 161878 160876 161880
rect 50613 161875 50679 161878
rect 160870 161876 160876 161878
rect 160940 161876 160946 161940
rect 200798 161876 200804 161940
rect 200868 161938 200874 161940
rect 315990 161938 316050 162694
rect 343398 162692 343404 162694
rect 343468 162692 343515 162696
rect 395982 162694 396028 162754
rect 396092 162752 396139 162756
rect 396134 162696 396139 162752
rect 396022 162692 396028 162694
rect 396092 162692 396139 162696
rect 343449 162691 343515 162692
rect 396073 162691 396139 162692
rect 397453 162754 397519 162757
rect 398238 162754 398298 163100
rect 401593 163099 401659 163102
rect 401726 163100 401732 163102
rect 401796 163100 401802 163164
rect 455781 163160 455828 163164
rect 455892 163162 455898 163164
rect 455781 163104 455786 163160
rect 455781 163100 455828 163104
rect 455892 163102 455938 163162
rect 455892 163100 455898 163102
rect 455781 163099 455847 163100
rect 418153 162892 418219 162893
rect 418102 162890 418108 162892
rect 418062 162830 418108 162890
rect 418172 162888 418219 162892
rect 418214 162832 418219 162888
rect 418102 162828 418108 162830
rect 418172 162828 418219 162832
rect 418153 162827 418219 162828
rect 397453 162752 398298 162754
rect 397453 162696 397458 162752
rect 397514 162696 398298 162752
rect 397453 162694 398298 162696
rect 398833 162754 398899 162757
rect 399518 162754 399524 162756
rect 398833 162752 399524 162754
rect 398833 162696 398838 162752
rect 398894 162696 399524 162752
rect 398833 162694 399524 162696
rect 397453 162691 397519 162694
rect 398833 162691 398899 162694
rect 399518 162692 399524 162694
rect 399588 162692 399594 162756
rect 400213 162754 400279 162757
rect 403065 162756 403131 162757
rect 400438 162754 400444 162756
rect 400213 162752 400444 162754
rect 400213 162696 400218 162752
rect 400274 162696 400444 162752
rect 400213 162694 400444 162696
rect 400213 162691 400279 162694
rect 400438 162692 400444 162694
rect 400508 162692 400514 162756
rect 403014 162754 403020 162756
rect 402974 162694 403020 162754
rect 403084 162752 403131 162756
rect 403126 162696 403131 162752
rect 403014 162692 403020 162694
rect 403084 162692 403131 162696
rect 403065 162691 403131 162692
rect 404353 162754 404419 162757
rect 405038 162754 405044 162756
rect 404353 162752 405044 162754
rect 404353 162696 404358 162752
rect 404414 162696 405044 162752
rect 404353 162694 405044 162696
rect 404353 162691 404419 162694
rect 405038 162692 405044 162694
rect 405108 162692 405114 162756
rect 405733 162754 405799 162757
rect 406510 162754 406516 162756
rect 405733 162752 406516 162754
rect 405733 162696 405738 162752
rect 405794 162696 406516 162752
rect 405733 162694 406516 162696
rect 405733 162691 405799 162694
rect 406510 162692 406516 162694
rect 406580 162692 406586 162756
rect 407205 162754 407271 162757
rect 408309 162756 408375 162757
rect 407614 162754 407620 162756
rect 407205 162752 407620 162754
rect 407205 162696 407210 162752
rect 407266 162696 407620 162752
rect 407205 162694 407620 162696
rect 407205 162691 407271 162694
rect 407614 162692 407620 162694
rect 407684 162692 407690 162756
rect 408309 162754 408356 162756
rect 408264 162752 408356 162754
rect 408264 162696 408314 162752
rect 408264 162694 408356 162696
rect 408309 162692 408356 162694
rect 408420 162692 408426 162756
rect 408493 162754 408559 162757
rect 409965 162756 410031 162757
rect 408718 162754 408724 162756
rect 408493 162752 408724 162754
rect 408493 162696 408498 162752
rect 408554 162696 408724 162752
rect 408493 162694 408724 162696
rect 408309 162691 408375 162692
rect 408493 162691 408559 162694
rect 408718 162692 408724 162694
rect 408788 162692 408794 162756
rect 409965 162752 410012 162756
rect 410076 162754 410082 162756
rect 410609 162754 410675 162757
rect 411345 162756 411411 162757
rect 410742 162754 410748 162756
rect 409965 162696 409970 162752
rect 409965 162692 410012 162696
rect 410076 162694 410122 162754
rect 410609 162752 410748 162754
rect 410609 162696 410614 162752
rect 410670 162696 410748 162752
rect 410609 162694 410748 162696
rect 410076 162692 410082 162694
rect 409965 162691 410031 162692
rect 410609 162691 410675 162694
rect 410742 162692 410748 162694
rect 410812 162692 410818 162756
rect 411294 162754 411300 162756
rect 411254 162694 411300 162754
rect 411364 162752 411411 162756
rect 411406 162696 411411 162752
rect 411294 162692 411300 162694
rect 411364 162692 411411 162696
rect 411345 162691 411411 162692
rect 412633 162754 412699 162757
rect 413645 162756 413711 162757
rect 413502 162754 413508 162756
rect 412633 162752 413508 162754
rect 412633 162696 412638 162752
rect 412694 162696 413508 162752
rect 412633 162694 413508 162696
rect 412633 162691 412699 162694
rect 413502 162692 413508 162694
rect 413572 162692 413578 162756
rect 413645 162752 413692 162756
rect 413756 162754 413762 162756
rect 414013 162754 414079 162757
rect 414606 162754 414612 162756
rect 413645 162696 413650 162752
rect 413645 162692 413692 162696
rect 413756 162694 413802 162754
rect 414013 162752 414612 162754
rect 414013 162696 414018 162752
rect 414074 162696 414612 162752
rect 414013 162694 414612 162696
rect 413756 162692 413762 162694
rect 413645 162691 413711 162692
rect 414013 162691 414079 162694
rect 414606 162692 414612 162694
rect 414676 162692 414682 162756
rect 415393 162754 415459 162757
rect 415526 162754 415532 162756
rect 415393 162752 415532 162754
rect 415393 162696 415398 162752
rect 415454 162696 415532 162752
rect 415393 162694 415532 162696
rect 415393 162691 415459 162694
rect 415526 162692 415532 162694
rect 415596 162692 415602 162756
rect 416773 162754 416839 162757
rect 416998 162754 417004 162756
rect 416773 162752 417004 162754
rect 416773 162696 416778 162752
rect 416834 162696 417004 162752
rect 416773 162694 417004 162696
rect 416773 162691 416839 162694
rect 416998 162692 417004 162694
rect 417068 162692 417074 162756
rect 418153 162754 418219 162757
rect 419206 162754 419212 162756
rect 418153 162752 419212 162754
rect 418153 162696 418158 162752
rect 418214 162696 419212 162752
rect 418153 162694 419212 162696
rect 418153 162691 418219 162694
rect 419206 162692 419212 162694
rect 419276 162692 419282 162756
rect 419533 162754 419599 162757
rect 420678 162754 420684 162756
rect 419533 162752 420684 162754
rect 419533 162696 419538 162752
rect 419594 162696 420684 162752
rect 419533 162694 420684 162696
rect 419533 162691 419599 162694
rect 420678 162692 420684 162694
rect 420748 162692 420754 162756
rect 420913 162754 420979 162757
rect 421782 162754 421788 162756
rect 420913 162752 421788 162754
rect 420913 162696 420918 162752
rect 420974 162696 421788 162752
rect 420913 162694 421788 162696
rect 420913 162691 420979 162694
rect 421782 162692 421788 162694
rect 421852 162692 421858 162756
rect 422293 162754 422359 162757
rect 422886 162754 422892 162756
rect 422293 162752 422892 162754
rect 422293 162696 422298 162752
rect 422354 162696 422892 162752
rect 422293 162694 422892 162696
rect 422293 162691 422359 162694
rect 422886 162692 422892 162694
rect 422956 162692 422962 162756
rect 423673 162754 423739 162757
rect 423990 162754 423996 162756
rect 423673 162752 423996 162754
rect 423673 162696 423678 162752
rect 423734 162696 423996 162752
rect 423673 162694 423996 162696
rect 423673 162691 423739 162694
rect 423990 162692 423996 162694
rect 424060 162692 424066 162756
rect 425053 162754 425119 162757
rect 426433 162756 426499 162757
rect 425278 162754 425284 162756
rect 425053 162752 425284 162754
rect 425053 162696 425058 162752
rect 425114 162696 425284 162752
rect 425053 162694 425284 162696
rect 425053 162691 425119 162694
rect 425278 162692 425284 162694
rect 425348 162692 425354 162756
rect 426382 162754 426388 162756
rect 426342 162694 426388 162754
rect 426452 162752 426499 162756
rect 426494 162696 426499 162752
rect 426382 162692 426388 162694
rect 426452 162692 426499 162696
rect 428774 162692 428780 162756
rect 428844 162754 428850 162756
rect 429101 162754 429167 162757
rect 428844 162752 429167 162754
rect 428844 162696 429106 162752
rect 429162 162696 429167 162752
rect 428844 162694 429167 162696
rect 428844 162692 428850 162694
rect 426433 162691 426499 162692
rect 429101 162691 429167 162694
rect 429285 162754 429351 162757
rect 429694 162754 429700 162756
rect 429285 162752 429700 162754
rect 429285 162696 429290 162752
rect 429346 162696 429700 162752
rect 429285 162694 429700 162696
rect 429285 162691 429351 162694
rect 429694 162692 429700 162694
rect 429764 162692 429770 162756
rect 430573 162754 430639 162757
rect 431166 162754 431172 162756
rect 430573 162752 431172 162754
rect 430573 162696 430578 162752
rect 430634 162696 431172 162752
rect 430573 162694 431172 162696
rect 430573 162691 430639 162694
rect 431166 162692 431172 162694
rect 431236 162692 431242 162756
rect 431718 162692 431724 162756
rect 431788 162754 431794 162756
rect 431953 162754 432019 162757
rect 431788 162752 432019 162754
rect 431788 162696 431958 162752
rect 432014 162696 432019 162752
rect 431788 162694 432019 162696
rect 431788 162692 431794 162694
rect 431953 162691 432019 162694
rect 433374 162692 433380 162756
rect 433444 162754 433450 162756
rect 434621 162754 434687 162757
rect 433444 162752 434687 162754
rect 433444 162696 434626 162752
rect 434682 162696 434687 162752
rect 433444 162694 434687 162696
rect 433444 162692 433450 162694
rect 434621 162691 434687 162694
rect 435357 162754 435423 162757
rect 435909 162756 435975 162757
rect 438485 162756 438551 162757
rect 439037 162756 439103 162757
rect 440877 162756 440943 162757
rect 443453 162756 443519 162757
rect 445845 162756 445911 162757
rect 448237 162756 448303 162757
rect 435766 162754 435772 162756
rect 435357 162752 435772 162754
rect 435357 162696 435362 162752
rect 435418 162696 435772 162752
rect 435357 162694 435772 162696
rect 435357 162691 435423 162694
rect 435766 162692 435772 162694
rect 435836 162692 435842 162756
rect 435909 162752 435956 162756
rect 436020 162754 436026 162756
rect 435909 162696 435914 162752
rect 435909 162692 435956 162696
rect 436020 162694 436066 162754
rect 438485 162752 438532 162756
rect 438596 162754 438602 162756
rect 438485 162696 438490 162752
rect 436020 162692 436026 162694
rect 438485 162692 438532 162696
rect 438596 162694 438642 162754
rect 439037 162752 439084 162756
rect 439148 162754 439154 162756
rect 439037 162696 439042 162752
rect 438596 162692 438602 162694
rect 439037 162692 439084 162696
rect 439148 162694 439194 162754
rect 440877 162752 440924 162756
rect 440988 162754 440994 162756
rect 440877 162696 440882 162752
rect 439148 162692 439154 162694
rect 440877 162692 440924 162696
rect 440988 162694 441034 162754
rect 443453 162752 443500 162756
rect 443564 162754 443570 162756
rect 443453 162696 443458 162752
rect 440988 162692 440994 162694
rect 443453 162692 443500 162696
rect 443564 162694 443610 162754
rect 445845 162752 445892 162756
rect 445956 162754 445962 162756
rect 445845 162696 445850 162752
rect 443564 162692 443570 162694
rect 445845 162692 445892 162696
rect 445956 162694 446002 162754
rect 448237 162752 448284 162756
rect 448348 162754 448354 162756
rect 453205 162754 453271 162757
rect 458357 162756 458423 162757
rect 453430 162754 453436 162756
rect 448237 162696 448242 162752
rect 445956 162692 445962 162694
rect 448237 162692 448284 162696
rect 448348 162694 448394 162754
rect 453205 162752 453436 162754
rect 453205 162696 453210 162752
rect 453266 162696 453436 162752
rect 453205 162694 453436 162696
rect 448348 162692 448354 162694
rect 435909 162691 435975 162692
rect 438485 162691 438551 162692
rect 439037 162691 439103 162692
rect 440877 162691 440943 162692
rect 443453 162691 443519 162692
rect 445845 162691 445911 162692
rect 448237 162691 448303 162692
rect 453205 162691 453271 162694
rect 453430 162692 453436 162694
rect 453500 162692 453506 162756
rect 458357 162752 458404 162756
rect 458468 162754 458474 162756
rect 458357 162696 458362 162752
rect 458357 162692 458404 162696
rect 458468 162694 458514 162754
rect 458468 162692 458474 162694
rect 503110 162692 503116 162756
rect 503180 162754 503186 162756
rect 503253 162754 503319 162757
rect 503180 162752 503319 162754
rect 503180 162696 503258 162752
rect 503314 162696 503319 162752
rect 503180 162694 503319 162696
rect 503180 162692 503186 162694
rect 458357 162691 458423 162692
rect 503253 162691 503319 162694
rect 320909 162620 320975 162621
rect 320909 162616 320956 162620
rect 321020 162618 321026 162620
rect 320909 162560 320914 162616
rect 320909 162556 320956 162560
rect 321020 162558 321066 162618
rect 321020 162556 321026 162558
rect 343214 162556 343220 162620
rect 343284 162618 343290 162620
rect 343357 162618 343423 162621
rect 343284 162616 343423 162618
rect 343284 162560 343362 162616
rect 343418 162560 343423 162616
rect 343284 162558 343423 162560
rect 343284 162556 343290 162558
rect 320909 162555 320975 162556
rect 343357 162555 343423 162558
rect 376201 162618 376267 162621
rect 465942 162618 465948 162620
rect 376201 162616 465948 162618
rect 376201 162560 376206 162616
rect 376262 162560 465948 162616
rect 376201 162558 465948 162560
rect 376201 162555 376267 162558
rect 465942 162556 465948 162558
rect 466012 162556 466018 162620
rect 503478 162556 503484 162620
rect 503548 162618 503554 162620
rect 503621 162618 503687 162621
rect 503548 162616 503687 162618
rect 503548 162560 503626 162616
rect 503682 162560 503687 162616
rect 503548 162558 503687 162560
rect 503548 162556 503554 162558
rect 503621 162555 503687 162558
rect 374729 162482 374795 162485
rect 462630 162482 462636 162484
rect 374729 162480 462636 162482
rect 374729 162424 374734 162480
rect 374790 162424 462636 162480
rect 374729 162422 462636 162424
rect 374729 162419 374795 162422
rect 462630 162420 462636 162422
rect 462700 162420 462706 162484
rect 379053 162346 379119 162349
rect 460974 162346 460980 162348
rect 379053 162344 460980 162346
rect 379053 162288 379058 162344
rect 379114 162288 460980 162344
rect 379053 162286 460980 162288
rect 379053 162283 379119 162286
rect 460974 162284 460980 162286
rect 461044 162284 461050 162348
rect 396165 162210 396231 162213
rect 397126 162210 397132 162212
rect 396165 162208 397132 162210
rect 396165 162152 396170 162208
rect 396226 162152 397132 162208
rect 396165 162150 397132 162152
rect 396165 162147 396231 162150
rect 397126 162148 397132 162150
rect 397196 162148 397202 162212
rect 402973 162210 403039 162213
rect 404118 162210 404124 162212
rect 402973 162208 404124 162210
rect 402973 162152 402978 162208
rect 403034 162152 404124 162208
rect 402973 162150 404124 162152
rect 402973 162147 403039 162150
rect 404118 162148 404124 162150
rect 404188 162148 404194 162212
rect 411253 162210 411319 162213
rect 418429 162212 418495 162213
rect 412398 162210 412404 162212
rect 411253 162208 412404 162210
rect 411253 162152 411258 162208
rect 411314 162152 412404 162208
rect 411253 162150 412404 162152
rect 411253 162147 411319 162150
rect 412398 162148 412404 162150
rect 412468 162148 412474 162212
rect 418429 162208 418476 162212
rect 418540 162210 418546 162212
rect 426525 162210 426591 162213
rect 433517 162212 433583 162213
rect 427670 162210 427676 162212
rect 418429 162152 418434 162208
rect 418429 162148 418476 162152
rect 418540 162150 418586 162210
rect 426525 162208 427676 162210
rect 426525 162152 426530 162208
rect 426586 162152 427676 162208
rect 426525 162150 427676 162152
rect 418540 162148 418546 162150
rect 418429 162147 418495 162148
rect 426525 162147 426591 162150
rect 427670 162148 427676 162150
rect 427740 162148 427746 162212
rect 433517 162208 433564 162212
rect 433628 162210 433634 162212
rect 433517 162152 433522 162208
rect 433517 162148 433564 162152
rect 433628 162150 433674 162210
rect 433628 162148 433634 162150
rect 433517 162147 433583 162148
rect 200868 161878 316050 161938
rect 378869 161938 378935 161941
rect 468518 161938 468524 161940
rect 378869 161936 468524 161938
rect 378869 161880 378874 161936
rect 378930 161880 468524 161936
rect 378869 161878 468524 161880
rect 200868 161876 200874 161878
rect 378869 161875 378935 161878
rect 468518 161876 468524 161878
rect 468588 161876 468594 161940
rect 84142 161468 84148 161532
rect 84212 161530 84218 161532
rect 84285 161530 84351 161533
rect 238753 161532 238819 161533
rect 84212 161528 84351 161530
rect 84212 161472 84290 161528
rect 84346 161472 84351 161528
rect 84212 161470 84351 161472
rect 84212 161468 84218 161470
rect 84285 161467 84351 161470
rect 238702 161468 238708 161532
rect 238772 161530 238819 161532
rect 238772 161528 238864 161530
rect 238814 161472 238864 161528
rect 238772 161470 238864 161472
rect 238772 161468 238819 161470
rect 277342 161468 277348 161532
rect 277412 161530 277418 161532
rect 278037 161530 278103 161533
rect 277412 161528 278103 161530
rect 277412 161472 278042 161528
rect 278098 161472 278103 161528
rect 277412 161470 278103 161472
rect 277412 161468 277418 161470
rect 238753 161467 238819 161468
rect 278037 161467 278103 161470
rect 55949 160170 56015 160173
rect 57646 160170 57652 160172
rect 55949 160168 57652 160170
rect 55949 160112 55954 160168
rect 56010 160112 57652 160168
rect 55949 160110 57652 160112
rect 55949 160107 56015 160110
rect 57646 160108 57652 160110
rect 57716 160108 57722 160172
rect 375465 158810 375531 158813
rect 377254 158810 377260 158812
rect 375465 158808 377260 158810
rect 375465 158752 375470 158808
rect 375526 158752 377260 158808
rect 375465 158750 377260 158752
rect 375465 158747 375531 158750
rect 377254 158748 377260 158750
rect 377324 158810 377330 158812
rect 378041 158810 378107 158813
rect 377324 158808 378107 158810
rect 377324 158752 378046 158808
rect 378102 158752 378107 158808
rect 377324 158750 378107 158752
rect 377324 158748 377330 158750
rect 378041 158747 378107 158750
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect -960 149774 674 149834
rect -960 149698 480 149774
rect 614 149698 674 149774
rect -960 149684 674 149698
rect 246 149638 674 149684
rect 246 149154 306 149638
rect 360694 149154 360700 149156
rect 246 149094 360700 149154
rect 360694 149092 360700 149094
rect 360764 149092 360770 149156
rect 278221 149018 278287 149021
rect 356789 149018 356855 149021
rect 278221 149016 356855 149018
rect 278221 148960 278226 149016
rect 278282 148960 356794 149016
rect 356850 148960 356855 149016
rect 278221 148958 356855 148960
rect 278221 148955 278287 148958
rect 356789 148955 356855 148958
rect 217358 148276 217364 148340
rect 217428 148338 217434 148340
rect 278221 148338 278287 148341
rect 217428 148336 278287 148338
rect 217428 148280 278226 148336
rect 278282 148280 278287 148336
rect 217428 148278 278287 148280
rect 217428 148276 217434 148278
rect 278221 148275 278287 148278
rect 217174 146372 217180 146436
rect 217244 146434 217250 146436
rect 276013 146434 276079 146437
rect 217244 146432 276079 146434
rect 217244 146376 276018 146432
rect 276074 146376 276079 146432
rect 217244 146374 276079 146376
rect 217244 146372 217250 146374
rect 276013 146371 276079 146374
rect 73797 146298 73863 146301
rect 100845 146298 100911 146301
rect 73797 146296 100911 146298
rect 73797 146240 73802 146296
rect 73858 146240 100850 146296
rect 100906 146240 100911 146296
rect 73797 146238 100911 146240
rect 73797 146235 73863 146238
rect 100845 146235 100911 146238
rect 214925 146298 214991 146301
rect 269113 146298 269179 146301
rect 214925 146296 269179 146298
rect 214925 146240 214930 146296
rect 214986 146240 269118 146296
rect 269174 146240 269179 146296
rect 214925 146238 269179 146240
rect 214925 146235 214991 146238
rect 269113 146235 269179 146238
rect 373901 146298 373967 146301
rect 376477 146298 376543 146301
rect 373901 146296 376543 146298
rect 373901 146240 373906 146296
rect 373962 146240 376482 146296
rect 376538 146240 376543 146296
rect 373901 146238 376543 146240
rect 373901 146235 373967 146238
rect 376477 146235 376543 146238
rect 377990 146236 377996 146300
rect 378060 146298 378066 146300
rect 425053 146298 425119 146301
rect 378060 146296 425119 146298
rect 378060 146240 425058 146296
rect 425114 146240 425119 146296
rect 378060 146238 425119 146240
rect 378060 146236 378066 146238
rect 425053 146235 425119 146238
rect 379697 146162 379763 146165
rect 415393 146162 415459 146165
rect 379697 146160 415459 146162
rect 379697 146104 379702 146160
rect 379758 146104 415398 146160
rect 415454 146104 415459 146160
rect 379697 146102 415459 146104
rect 379697 146099 379763 146102
rect 415393 146099 415459 146102
rect 510613 146162 510679 146165
rect 510838 146162 510844 146164
rect 510613 146160 510844 146162
rect 510613 146104 510618 146160
rect 510674 146104 510844 146160
rect 510613 146102 510844 146104
rect 510613 146099 510679 146102
rect 510838 146100 510844 146102
rect 510908 146100 510914 146164
rect 57462 145964 57468 146028
rect 57532 146026 57538 146028
rect 87597 146026 87663 146029
rect 57532 146024 87663 146026
rect 57532 145968 87602 146024
rect 87658 145968 87663 146024
rect 57532 145966 87663 145968
rect 57532 145964 57538 145966
rect 87597 145963 87663 145966
rect 217542 145964 217548 146028
rect 217612 146026 217618 146028
rect 217869 146026 217935 146029
rect 217612 146024 217935 146026
rect 217612 145968 217874 146024
rect 217930 145968 217935 146024
rect 217612 145966 217935 145968
rect 217612 145964 217618 145966
rect 217869 145963 217935 145966
rect 378869 146026 378935 146029
rect 412633 146026 412699 146029
rect 378869 146024 412699 146026
rect 378869 145968 378874 146024
rect 378930 145968 412638 146024
rect 412694 145968 412699 146024
rect 378869 145966 412699 145968
rect 378869 145963 378935 145966
rect 412633 145963 412699 145966
rect 58617 145890 58683 145893
rect 92473 145890 92539 145893
rect 58617 145888 92539 145890
rect 58617 145832 58622 145888
rect 58678 145832 92478 145888
rect 92534 145832 92539 145888
rect 58617 145830 92539 145832
rect 58617 145827 58683 145830
rect 92473 145827 92539 145830
rect 214557 145890 214623 145893
rect 237373 145890 237439 145893
rect 214557 145888 237439 145890
rect 214557 145832 214562 145888
rect 214618 145832 237378 145888
rect 237434 145832 237439 145888
rect 214557 145830 237439 145832
rect 214557 145827 214623 145830
rect 237373 145827 237439 145830
rect 54293 145754 54359 145757
rect 58525 145754 58591 145757
rect 102133 145754 102199 145757
rect 54293 145752 102199 145754
rect 54293 145696 54298 145752
rect 54354 145696 58530 145752
rect 58586 145696 102138 145752
rect 102194 145696 102199 145752
rect 54293 145694 102199 145696
rect 54293 145691 54359 145694
rect 58525 145691 58591 145694
rect 102133 145691 102199 145694
rect 214649 145754 214715 145757
rect 270493 145754 270559 145757
rect 214649 145752 270559 145754
rect 214649 145696 214654 145752
rect 214710 145696 270498 145752
rect 270554 145696 270559 145752
rect 214649 145694 270559 145696
rect 214649 145691 214715 145694
rect 270493 145691 270559 145694
rect 56409 145618 56475 145621
rect 100753 145618 100819 145621
rect 56409 145616 100819 145618
rect 56409 145560 56414 145616
rect 56470 145560 100758 145616
rect 100814 145560 100819 145616
rect 56409 145558 100819 145560
rect 56409 145555 56475 145558
rect 100753 145555 100819 145558
rect 215845 145618 215911 145621
rect 271873 145618 271939 145621
rect 215845 145616 271939 145618
rect 215845 145560 215850 145616
rect 215906 145560 271878 145616
rect 271934 145560 271939 145616
rect 215845 145558 271939 145560
rect 215845 145555 215911 145558
rect 271873 145555 271939 145558
rect 375925 145618 375991 145621
rect 376477 145618 376543 145621
rect 423673 145618 423739 145621
rect 375925 145616 423739 145618
rect 375925 145560 375930 145616
rect 375986 145560 376482 145616
rect 376538 145560 423678 145616
rect 423734 145560 423739 145616
rect 375925 145558 423739 145560
rect 375925 145555 375991 145558
rect 376477 145555 376543 145558
rect 423673 145555 423739 145558
rect 190862 145420 190868 145484
rect 190932 145482 190938 145484
rect 191741 145482 191807 145485
rect 190932 145480 191807 145482
rect 190932 145424 191746 145480
rect 191802 145424 191807 145480
rect 190932 145422 191807 145424
rect 190932 145420 190938 145422
rect 191741 145419 191807 145422
rect 178534 144876 178540 144940
rect 178604 144938 178610 144940
rect 179045 144938 179111 144941
rect 179689 144940 179755 144941
rect 338481 144940 338547 144941
rect 179638 144938 179644 144940
rect 178604 144936 179111 144938
rect 178604 144880 179050 144936
rect 179106 144880 179111 144936
rect 178604 144878 179111 144880
rect 179598 144878 179644 144938
rect 179708 144936 179755 144940
rect 338430 144938 338436 144940
rect 179750 144880 179755 144936
rect 178604 144876 178610 144878
rect 179045 144875 179111 144878
rect 179638 144876 179644 144878
rect 179708 144876 179755 144880
rect 338390 144878 338436 144938
rect 338500 144936 338547 144940
rect 338542 144880 338547 144936
rect 338430 144876 338436 144878
rect 338500 144876 338547 144880
rect 339718 144876 339724 144940
rect 339788 144938 339794 144940
rect 340229 144938 340295 144941
rect 339788 144936 340295 144938
rect 339788 144880 340234 144936
rect 340290 144880 340295 144936
rect 339788 144878 340295 144880
rect 339788 144876 339794 144878
rect 179689 144875 179755 144876
rect 338481 144875 338547 144876
rect 340229 144875 340295 144878
rect 350942 144876 350948 144940
rect 351012 144938 351018 144940
rect 351637 144938 351703 144941
rect 351012 144936 351703 144938
rect 351012 144880 351642 144936
rect 351698 144880 351703 144936
rect 351012 144878 351703 144880
rect 351012 144876 351018 144878
rect 351637 144875 351703 144878
rect 498510 144876 498516 144940
rect 498580 144938 498586 144940
rect 498653 144938 498719 144941
rect 499849 144940 499915 144941
rect 499798 144938 499804 144940
rect 498580 144936 498719 144938
rect 498580 144880 498658 144936
rect 498714 144880 498719 144936
rect 498580 144878 498719 144880
rect 499758 144878 499804 144938
rect 499868 144936 499915 144940
rect 499910 144880 499915 144936
rect 498580 144876 498586 144878
rect 498653 144875 498719 144878
rect 499798 144876 499804 144878
rect 499868 144876 499915 144880
rect 499849 144875 499915 144876
rect 47853 144802 47919 144805
rect 57094 144802 57100 144804
rect 47853 144800 57100 144802
rect 47853 144744 47858 144800
rect 47914 144744 57100 144800
rect 47853 144742 57100 144744
rect 47853 144739 47919 144742
rect 57094 144740 57100 144742
rect 57164 144802 57170 144804
rect 57462 144802 57468 144804
rect 57164 144742 57468 144802
rect 57164 144740 57170 144742
rect 57462 144740 57468 144742
rect 57532 144740 57538 144804
rect 372429 144122 372495 144125
rect 377949 144122 378015 144125
rect 372429 144120 378015 144122
rect 372429 144064 372434 144120
rect 372490 144064 377954 144120
rect 378010 144064 378015 144120
rect 372429 144062 378015 144064
rect 372429 144059 372495 144062
rect 377949 144059 378015 144062
rect 377438 143652 377444 143716
rect 377508 143714 377514 143716
rect 377949 143714 378015 143717
rect 377508 143712 378015 143714
rect 377508 143656 377954 143712
rect 378010 143656 378015 143712
rect 377508 143654 378015 143656
rect 377508 143652 377514 143654
rect 377949 143651 378015 143654
rect 57462 140796 57468 140860
rect 57532 140858 57538 140860
rect 59353 140858 59419 140861
rect 57532 140856 59419 140858
rect 57532 140800 59358 140856
rect 59414 140800 59419 140856
rect 57532 140798 59419 140800
rect 57532 140796 57538 140798
rect 59353 140795 59419 140798
rect 359273 139362 359339 139365
rect 519353 139362 519419 139365
rect 356562 139360 359339 139362
rect 356562 139304 359278 139360
rect 359334 139304 359339 139360
rect 356562 139302 359339 139304
rect 199193 139226 199259 139229
rect 197126 139224 199259 139226
rect 197126 139220 199198 139224
rect 196604 139168 199198 139220
rect 199254 139168 199259 139224
rect 356562 139190 356622 139302
rect 359273 139299 359339 139302
rect 516558 139360 519419 139362
rect 516558 139304 519358 139360
rect 519414 139304 519419 139360
rect 516558 139302 519419 139304
rect 516558 139190 516618 139302
rect 519353 139299 519419 139302
rect 583520 139212 584960 139452
rect 196604 139166 199259 139168
rect 196604 139160 197186 139166
rect 199193 139163 199259 139166
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 57053 97474 57119 97477
rect 57053 97472 60062 97474
rect 57053 97416 57058 97472
rect 57114 97416 60062 97472
rect 57053 97414 60062 97416
rect 57053 97411 57119 97414
rect 60002 96894 60062 97414
rect 216857 96930 216923 96933
rect 377489 96930 377555 96933
rect 216857 96928 219450 96930
rect 216857 96872 216862 96928
rect 216918 96924 219450 96928
rect 377489 96928 379530 96930
rect 216918 96872 220064 96924
rect 216857 96870 220064 96872
rect 216857 96867 216923 96870
rect 219390 96864 220064 96870
rect 377489 96872 377494 96928
rect 377550 96924 379530 96928
rect 377550 96872 380052 96924
rect 377489 96870 380052 96872
rect 377489 96867 377555 96870
rect 379470 96864 380052 96870
rect 57145 96522 57211 96525
rect 57145 96520 60062 96522
rect 57145 96464 57150 96520
rect 57206 96464 60062 96520
rect 57145 96462 60062 96464
rect 57145 96459 57211 96462
rect 60002 95942 60062 96462
rect 216949 95978 217015 95981
rect 376937 95978 377003 95981
rect 216949 95976 219450 95978
rect 216949 95920 216954 95976
rect 217010 95972 219450 95976
rect 376937 95976 379530 95978
rect 217010 95920 220064 95972
rect 216949 95918 220064 95920
rect 216949 95915 217015 95918
rect 219390 95912 220064 95918
rect 376937 95920 376942 95976
rect 376998 95972 379530 95976
rect 376998 95920 380052 95972
rect 376937 95918 380052 95920
rect 376937 95915 377003 95918
rect 379470 95912 380052 95918
rect 56869 93802 56935 93805
rect 217961 93802 218027 93805
rect 377857 93802 377923 93805
rect 56869 93800 60062 93802
rect 56869 93744 56874 93800
rect 56930 93744 60062 93800
rect 56869 93742 60062 93744
rect 217961 93800 219450 93802
rect 217961 93744 217966 93800
rect 218022 93796 219450 93800
rect 377857 93800 379530 93802
rect 218022 93744 220064 93796
rect 217961 93742 220064 93744
rect 56869 93739 56935 93742
rect 217961 93739 218027 93742
rect 219390 93736 220064 93742
rect 377857 93744 377862 93800
rect 377918 93796 379530 93800
rect 377918 93744 380052 93796
rect 377857 93742 380052 93744
rect 377857 93739 377923 93742
rect 379470 93736 380052 93742
rect 57329 93394 57395 93397
rect 57329 93392 60062 93394
rect 57329 93336 57334 93392
rect 57390 93336 60062 93392
rect 57329 93334 60062 93336
rect 57329 93331 57395 93334
rect 60002 92814 60062 93334
rect 217225 92850 217291 92853
rect 377581 92850 377647 92853
rect 217225 92848 219450 92850
rect 217225 92792 217230 92848
rect 217286 92844 219450 92848
rect 377581 92848 379530 92850
rect 217286 92792 220064 92844
rect 217225 92790 220064 92792
rect 217225 92787 217291 92790
rect 219390 92784 220064 92790
rect 377581 92792 377586 92848
rect 377642 92844 379530 92848
rect 377642 92792 380052 92844
rect 377581 92790 380052 92792
rect 377581 92787 377647 92790
rect 379470 92784 380052 92790
rect 57697 91082 57763 91085
rect 217685 91082 217751 91085
rect 377765 91082 377831 91085
rect 57697 91080 60062 91082
rect 57697 91024 57702 91080
rect 57758 91024 60062 91080
rect 57697 91022 60062 91024
rect 217685 91080 219450 91082
rect 217685 91024 217690 91080
rect 217746 91076 219450 91080
rect 377765 91080 379530 91082
rect 217746 91024 220064 91076
rect 217685 91022 220064 91024
rect 57697 91019 57763 91022
rect 217685 91019 217751 91022
rect 219390 91016 220064 91022
rect 377765 91024 377770 91080
rect 377826 91076 379530 91080
rect 377826 91024 380052 91076
rect 377765 91022 380052 91024
rect 377765 91019 377831 91022
rect 379470 91016 380052 91022
rect 57513 90538 57579 90541
rect 57513 90536 60062 90538
rect 57513 90480 57518 90536
rect 57574 90480 60062 90536
rect 57513 90478 60062 90480
rect 57513 90475 57579 90478
rect 60002 89958 60062 90478
rect 217409 89994 217475 89997
rect 377305 89994 377371 89997
rect 217409 89992 219450 89994
rect 217409 89936 217414 89992
rect 217470 89988 219450 89992
rect 377305 89992 379530 89994
rect 217470 89936 220064 89988
rect 217409 89934 220064 89936
rect 217409 89931 217475 89934
rect 219390 89928 220064 89934
rect 377305 89936 377310 89992
rect 377366 89988 379530 89992
rect 377366 89936 380052 89988
rect 377305 89934 380052 89936
rect 377305 89931 377371 89934
rect 379470 89928 380052 89934
rect 57421 88226 57487 88229
rect 217501 88226 217567 88229
rect 377673 88226 377739 88229
rect 57421 88224 60062 88226
rect 57421 88168 57426 88224
rect 57482 88168 60062 88224
rect 57421 88166 60062 88168
rect 217501 88224 219450 88226
rect 217501 88168 217506 88224
rect 217562 88220 219450 88224
rect 377673 88224 379530 88226
rect 217562 88168 220064 88220
rect 217501 88166 220064 88168
rect 57421 88163 57487 88166
rect 217501 88163 217567 88166
rect 219390 88160 220064 88166
rect 377673 88168 377678 88224
rect 377734 88220 379530 88224
rect 377734 88168 380052 88220
rect 377673 88166 380052 88168
rect 377673 88163 377739 88166
rect 379470 88160 380052 88166
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 358997 79930 359063 79933
rect 518893 79930 518959 79933
rect 520181 79930 520247 79933
rect 356562 79928 359063 79930
rect 356562 79872 359002 79928
rect 359058 79872 359063 79928
rect 356562 79870 359063 79872
rect 199377 79386 199443 79389
rect 197126 79384 199443 79386
rect 197126 79380 199382 79384
rect 196604 79328 199382 79380
rect 199438 79328 199443 79384
rect 356562 79350 356622 79870
rect 358997 79867 359063 79870
rect 516558 79928 520247 79930
rect 516558 79872 518898 79928
rect 518954 79872 520186 79928
rect 520242 79872 520247 79928
rect 516558 79870 520247 79872
rect 516558 79350 516618 79870
rect 518893 79867 518959 79870
rect 520181 79867 520247 79870
rect 196604 79326 199443 79328
rect 196604 79320 197186 79326
rect 199377 79323 199443 79326
rect 358813 78298 358879 78301
rect 518985 78298 519051 78301
rect 356562 78296 358879 78298
rect 356562 78240 358818 78296
rect 358874 78240 358879 78296
rect 356562 78238 358879 78240
rect 199285 77754 199351 77757
rect 197126 77752 199351 77754
rect 197126 77748 199290 77752
rect 196604 77696 199290 77748
rect 199346 77696 199351 77752
rect 356562 77718 356622 78238
rect 358813 78235 358879 78238
rect 516558 78296 519051 78298
rect 516558 78240 518990 78296
rect 519046 78240 519051 78296
rect 516558 78238 519051 78240
rect 516558 77718 516618 78238
rect 518985 78235 519051 78238
rect 196604 77694 199351 77696
rect 196604 77688 197186 77694
rect 199285 77691 199351 77694
rect 359181 76938 359247 76941
rect 356562 76936 359247 76938
rect 356562 76880 359186 76936
rect 359242 76880 359247 76936
rect 356562 76878 359247 76880
rect 199101 76394 199167 76397
rect 197126 76392 199167 76394
rect 197126 76388 199106 76392
rect 196604 76336 199106 76388
rect 199162 76336 199167 76392
rect 356562 76358 356622 76878
rect 359181 76875 359247 76878
rect 519261 76802 519327 76805
rect 516558 76800 519327 76802
rect 516558 76744 519266 76800
rect 519322 76744 519327 76800
rect 516558 76742 519327 76744
rect 516558 76358 516618 76742
rect 519261 76739 519327 76742
rect 196604 76334 199167 76336
rect 196604 76328 197186 76334
rect 199101 76331 199167 76334
rect 358905 75442 358971 75445
rect 519445 75442 519511 75445
rect 356562 75440 358971 75442
rect 356562 75384 358910 75440
rect 358966 75384 358971 75440
rect 356562 75382 358971 75384
rect 198733 74898 198799 74901
rect 197126 74896 198799 74898
rect 197126 74892 198738 74896
rect 196604 74840 198738 74892
rect 198794 74840 198799 74896
rect 356562 74862 356622 75382
rect 358905 75379 358971 75382
rect 516558 75440 519511 75442
rect 516558 75384 519450 75440
rect 519506 75384 519511 75440
rect 516558 75382 519511 75384
rect 516558 74862 516618 75382
rect 519445 75379 519511 75382
rect 196604 74838 198799 74840
rect 196604 74832 197186 74838
rect 198733 74835 198799 74838
rect 519077 74218 519143 74221
rect 516558 74216 519143 74218
rect 516558 74160 519082 74216
rect 519138 74160 519143 74216
rect 516558 74158 519143 74160
rect 359089 74082 359155 74085
rect 356562 74080 359155 74082
rect 356562 74024 359094 74080
rect 359150 74024 359155 74080
rect 356562 74022 359155 74024
rect 198825 73674 198891 73677
rect 197126 73672 198891 73674
rect 197126 73668 198830 73672
rect 196604 73616 198830 73668
rect 198886 73616 198891 73672
rect 356562 73638 356622 74022
rect 359089 74019 359155 74022
rect 516558 73638 516618 74158
rect 519077 74155 519143 74158
rect 196604 73614 198891 73616
rect 196604 73608 197186 73614
rect 198825 73611 198891 73614
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 57830 70348 57836 70412
rect 57900 70410 57906 70412
rect 57900 70350 60062 70410
rect 57900 70348 57906 70350
rect 60002 69966 60062 70350
rect 208894 69940 208900 70004
rect 208964 70002 208970 70004
rect 376937 70002 377003 70005
rect 208964 69996 219450 70002
rect 376937 70000 379530 70002
rect 208964 69942 220064 69996
rect 208964 69940 208970 69942
rect 219390 69936 220064 69942
rect 376937 69944 376942 70000
rect 376998 69996 379530 70000
rect 376998 69944 380052 69996
rect 376937 69942 380052 69944
rect 376937 69939 377003 69942
rect 379470 69936 380052 69942
rect 57881 68914 57947 68917
rect 57881 68912 60062 68914
rect 57881 68856 57886 68912
rect 57942 68856 60062 68912
rect 57881 68854 60062 68856
rect 57881 68851 57947 68854
rect 60002 68334 60062 68854
rect 216673 68370 216739 68373
rect 217961 68370 218027 68373
rect 376937 68370 377003 68373
rect 216673 68368 219450 68370
rect 216673 68312 216678 68368
rect 216734 68312 217966 68368
rect 218022 68364 219450 68368
rect 376937 68368 379530 68370
rect 218022 68312 220064 68364
rect 216673 68310 220064 68312
rect 216673 68307 216739 68310
rect 217961 68307 218027 68310
rect 219390 68304 220064 68310
rect 376937 68312 376942 68368
rect 376998 68364 379530 68368
rect 376998 68312 380052 68364
rect 376937 68310 380052 68312
rect 376937 68307 377003 68310
rect 379470 68304 380052 68310
rect 46790 67764 46796 67828
rect 46860 67826 46866 67828
rect 60002 67826 60062 68062
rect 206134 68036 206140 68100
rect 206204 68098 206210 68100
rect 377305 68098 377371 68101
rect 206204 68092 219450 68098
rect 377305 68096 379530 68098
rect 206204 68038 220064 68092
rect 206204 68036 206210 68038
rect 219390 68032 220064 68038
rect 377305 68040 377310 68096
rect 377366 68092 379530 68096
rect 377366 68040 380052 68092
rect 377305 68038 380052 68040
rect 377305 68035 377371 68038
rect 379470 68032 380052 68038
rect 46860 67766 60062 67826
rect 46860 67764 46866 67766
rect 218646 60556 218652 60620
rect 218716 60618 218722 60620
rect 218973 60618 219039 60621
rect 219249 60620 219315 60621
rect 219198 60618 219204 60620
rect 218716 60616 219039 60618
rect 218716 60560 218978 60616
rect 219034 60560 219039 60616
rect 218716 60558 219039 60560
rect 219158 60558 219204 60618
rect 219268 60616 219315 60620
rect 219310 60560 219315 60616
rect 218716 60556 218722 60558
rect 218973 60555 219039 60558
rect 219198 60556 219204 60558
rect 219268 60556 219315 60560
rect 219249 60555 219315 60556
rect 77109 59804 77175 59805
rect 83089 59804 83155 59805
rect 99465 59804 99531 59805
rect 77109 59800 77142 59804
rect 77206 59802 77212 59804
rect 77109 59744 77114 59800
rect 77109 59740 77142 59744
rect 77206 59742 77266 59802
rect 83089 59800 83126 59804
rect 83190 59802 83196 59804
rect 99440 59802 99446 59804
rect 83089 59744 83094 59800
rect 77206 59740 77212 59742
rect 83089 59740 83126 59744
rect 83190 59742 83246 59802
rect 99374 59742 99446 59802
rect 99510 59800 99531 59804
rect 99526 59744 99531 59800
rect 83190 59740 83196 59742
rect 99440 59740 99446 59742
rect 99510 59740 99531 59744
rect 77109 59739 77175 59740
rect 83089 59739 83155 59740
rect 99465 59739 99531 59740
rect 113541 59804 113607 59805
rect 120901 59804 120967 59805
rect 237097 59804 237163 59805
rect 255865 59804 255931 59805
rect 259453 59804 259519 59805
rect 113541 59800 113590 59804
rect 113654 59802 113660 59804
rect 113541 59744 113546 59800
rect 113541 59740 113590 59744
rect 113654 59742 113698 59802
rect 120901 59800 120934 59804
rect 120998 59802 121004 59804
rect 120901 59744 120906 59800
rect 113654 59740 113660 59742
rect 120901 59740 120934 59744
rect 120998 59742 121058 59802
rect 237097 59800 237142 59804
rect 237206 59802 237212 59804
rect 237097 59744 237102 59800
rect 120998 59740 121004 59742
rect 237097 59740 237142 59744
rect 237206 59742 237254 59802
rect 255865 59800 255910 59804
rect 255974 59802 255980 59804
rect 259440 59802 259446 59804
rect 255865 59744 255870 59800
rect 237206 59740 237212 59742
rect 255865 59740 255910 59744
rect 255974 59742 256022 59802
rect 259362 59742 259446 59802
rect 259510 59800 259519 59804
rect 259514 59744 259519 59800
rect 255974 59740 255980 59742
rect 259440 59740 259446 59742
rect 259510 59740 259519 59744
rect 113541 59739 113607 59740
rect 120901 59739 120967 59740
rect 237097 59739 237163 59740
rect 255865 59739 255931 59740
rect 259453 59739 259519 59740
rect 260649 59804 260715 59805
rect 261753 59804 261819 59805
rect 263869 59804 263935 59805
rect 396073 59804 396139 59805
rect 260649 59800 260670 59804
rect 260734 59802 260740 59804
rect 260649 59744 260654 59800
rect 260649 59740 260670 59744
rect 260734 59742 260806 59802
rect 260734 59740 260740 59742
rect 261752 59740 261758 59804
rect 261822 59802 261828 59804
rect 261822 59742 261910 59802
rect 263869 59800 263934 59804
rect 263869 59744 263874 59800
rect 263930 59744 263934 59800
rect 261822 59740 261828 59742
rect 263869 59740 263934 59744
rect 263998 59802 264004 59804
rect 396048 59802 396054 59804
rect 263998 59742 264026 59802
rect 395982 59742 396054 59802
rect 396118 59800 396139 59804
rect 396134 59744 396139 59800
rect 263998 59740 264004 59742
rect 396048 59740 396054 59742
rect 396118 59740 396139 59744
rect 260649 59739 260715 59740
rect 261753 59739 261819 59740
rect 263869 59739 263935 59740
rect 396073 59739 396139 59740
rect 397085 59804 397151 59805
rect 416957 59804 417023 59805
rect 418429 59804 418495 59805
rect 422845 59804 422911 59805
rect 423949 59804 424015 59805
rect 397085 59800 397142 59804
rect 397206 59802 397212 59804
rect 397085 59744 397090 59800
rect 397085 59740 397142 59744
rect 397206 59742 397242 59802
rect 416957 59800 416998 59804
rect 417062 59802 417068 59804
rect 416957 59744 416962 59800
rect 397206 59740 397212 59742
rect 416957 59740 416998 59744
rect 417062 59742 417114 59802
rect 418429 59800 418494 59804
rect 418429 59744 418434 59800
rect 418490 59744 418494 59800
rect 417062 59740 417068 59742
rect 418429 59740 418494 59744
rect 418558 59802 418564 59804
rect 422840 59802 422846 59804
rect 418558 59742 418586 59802
rect 422754 59742 422846 59802
rect 418558 59740 418564 59742
rect 422840 59740 422846 59742
rect 422910 59740 422916 59804
rect 423928 59802 423934 59804
rect 423858 59742 423934 59802
rect 423998 59800 424015 59804
rect 424010 59744 424015 59800
rect 423928 59740 423934 59742
rect 423998 59740 424015 59744
rect 397085 59739 397151 59740
rect 416957 59739 417023 59740
rect 418429 59739 418495 59740
rect 422845 59739 422911 59740
rect 423949 59739 424015 59740
rect 94497 59668 94563 59669
rect 102777 59668 102843 59669
rect 113265 59668 113331 59669
rect 116945 59668 117011 59669
rect 256969 59668 257035 59669
rect 258073 59668 258139 59669
rect 265249 59668 265315 59669
rect 315849 59668 315915 59669
rect 403065 59668 403131 59669
rect 404169 59668 404235 59669
rect 94497 59664 94550 59668
rect 94614 59666 94620 59668
rect 94497 59608 94502 59664
rect 94497 59604 94550 59608
rect 94614 59606 94654 59666
rect 102777 59664 102846 59668
rect 102777 59608 102782 59664
rect 102838 59608 102846 59664
rect 94614 59604 94620 59606
rect 102777 59604 102846 59608
rect 102910 59666 102916 59668
rect 102910 59606 102934 59666
rect 102910 59604 102916 59606
rect 105968 59604 105974 59668
rect 106038 59604 106044 59668
rect 113265 59664 113318 59668
rect 113382 59666 113388 59668
rect 113265 59608 113270 59664
rect 113265 59604 113318 59608
rect 113382 59606 113422 59666
rect 116945 59664 116990 59668
rect 117054 59666 117060 59668
rect 116945 59608 116950 59664
rect 113382 59604 113388 59606
rect 116945 59604 116990 59608
rect 117054 59606 117102 59666
rect 256969 59664 256998 59668
rect 257062 59666 257068 59668
rect 256969 59608 256974 59664
rect 117054 59604 117060 59606
rect 256969 59604 256998 59608
rect 257062 59606 257126 59666
rect 258073 59664 258086 59668
rect 258150 59666 258156 59668
rect 258073 59608 258078 59664
rect 257062 59604 257068 59606
rect 258073 59604 258086 59608
rect 258150 59606 258230 59666
rect 265249 59664 265294 59668
rect 265358 59666 265364 59668
rect 265249 59608 265254 59664
rect 258150 59604 258156 59606
rect 265249 59604 265294 59608
rect 265358 59606 265406 59666
rect 315849 59664 315886 59668
rect 315950 59666 315956 59668
rect 315849 59608 315854 59664
rect 265358 59604 265364 59606
rect 315849 59604 315886 59608
rect 315950 59606 316006 59666
rect 403065 59664 403126 59668
rect 403065 59608 403070 59664
rect 315950 59604 315956 59606
rect 403065 59604 403126 59608
rect 403190 59666 403196 59668
rect 403190 59606 403222 59666
rect 404169 59664 404214 59668
rect 404278 59666 404284 59668
rect 412541 59666 412607 59669
rect 423489 59668 423555 59669
rect 480897 59668 480963 59669
rect 413456 59666 413462 59668
rect 404169 59608 404174 59664
rect 403190 59604 403196 59606
rect 404169 59604 404214 59608
rect 404278 59606 404326 59666
rect 412541 59664 413462 59666
rect 412541 59608 412546 59664
rect 412602 59608 413462 59664
rect 412541 59606 413462 59608
rect 404278 59604 404284 59606
rect 94497 59603 94563 59604
rect 102777 59603 102843 59604
rect 46606 59468 46612 59532
rect 46676 59530 46682 59532
rect 105976 59530 106036 59604
rect 113265 59603 113331 59604
rect 116945 59603 117011 59604
rect 256969 59603 257035 59604
rect 258073 59603 258139 59604
rect 265249 59603 265315 59604
rect 315849 59603 315915 59604
rect 403065 59603 403131 59604
rect 404169 59603 404235 59604
rect 412541 59603 412607 59606
rect 413456 59604 413462 59606
rect 413526 59604 413532 59668
rect 423489 59664 423526 59668
rect 423590 59666 423596 59668
rect 423489 59608 423494 59664
rect 423489 59604 423526 59608
rect 423590 59606 423646 59666
rect 480897 59664 480918 59668
rect 480982 59666 480988 59668
rect 480897 59608 480902 59664
rect 423590 59604 423596 59606
rect 480897 59604 480918 59608
rect 480982 59606 481054 59666
rect 480982 59604 480988 59606
rect 423489 59603 423555 59604
rect 480897 59603 480963 59604
rect 46676 59470 106036 59530
rect 262765 59532 262831 59533
rect 418153 59532 418219 59533
rect 262765 59528 262812 59532
rect 262876 59530 262882 59532
rect 418102 59530 418108 59532
rect 262765 59472 262770 59528
rect 46676 59468 46682 59470
rect 262765 59468 262812 59472
rect 262876 59470 262922 59530
rect 418062 59470 418108 59530
rect 418172 59528 418219 59532
rect 418214 59472 418219 59528
rect 583520 59516 584960 59756
rect 262876 59468 262882 59470
rect 418102 59468 418108 59470
rect 418172 59468 418219 59472
rect 262765 59467 262831 59468
rect 418153 59467 418219 59468
rect 95877 59396 95943 59397
rect 98085 59396 98151 59397
rect 100753 59396 100819 59397
rect 95877 59392 95924 59396
rect 95988 59394 95994 59396
rect 95877 59336 95882 59392
rect 95877 59332 95924 59336
rect 95988 59334 96034 59394
rect 98085 59392 98132 59396
rect 98196 59394 98202 59396
rect 100702 59394 100708 59396
rect 98085 59336 98090 59392
rect 95988 59332 95994 59334
rect 98085 59332 98132 59336
rect 98196 59334 98242 59394
rect 100662 59334 100708 59394
rect 100772 59392 100819 59396
rect 100814 59336 100819 59392
rect 98196 59332 98202 59334
rect 100702 59332 100708 59334
rect 100772 59332 100819 59336
rect 95877 59331 95943 59332
rect 98085 59331 98151 59332
rect 100753 59331 100819 59332
rect 101765 59396 101831 59397
rect 420637 59396 420703 59397
rect 421741 59396 421807 59397
rect 425973 59396 426039 59397
rect 428181 59396 428247 59397
rect 453389 59396 453455 59397
rect 463509 59396 463575 59397
rect 101765 59392 101812 59396
rect 101876 59394 101882 59396
rect 101765 59336 101770 59392
rect 101765 59332 101812 59336
rect 101876 59334 101922 59394
rect 101876 59332 101882 59334
rect 197854 59332 197860 59396
rect 197924 59394 197930 59396
rect 263542 59394 263548 59396
rect 197924 59334 263548 59394
rect 197924 59332 197930 59334
rect 263542 59332 263548 59334
rect 263612 59332 263618 59396
rect 420637 59392 420684 59396
rect 420748 59394 420754 59396
rect 420637 59336 420642 59392
rect 420637 59332 420684 59336
rect 420748 59334 420794 59394
rect 421741 59392 421788 59396
rect 421852 59394 421858 59396
rect 421741 59336 421746 59392
rect 420748 59332 420754 59334
rect 421741 59332 421788 59336
rect 421852 59334 421898 59394
rect 425973 59392 426020 59396
rect 426084 59394 426090 59396
rect 425973 59336 425978 59392
rect 421852 59332 421858 59334
rect 425973 59332 426020 59336
rect 426084 59334 426130 59394
rect 428181 59392 428228 59396
rect 428292 59394 428298 59396
rect 428181 59336 428186 59392
rect 426084 59332 426090 59334
rect 428181 59332 428228 59336
rect 428292 59334 428338 59394
rect 453389 59392 453436 59396
rect 453500 59394 453506 59396
rect 453389 59336 453394 59392
rect 428292 59332 428298 59334
rect 453389 59332 453436 59336
rect 453500 59334 453546 59394
rect 463509 59392 463556 59396
rect 463620 59394 463626 59396
rect 463509 59336 463514 59392
rect 453500 59332 453506 59334
rect 463509 59332 463556 59336
rect 463620 59334 463666 59394
rect 463620 59332 463626 59334
rect 101765 59331 101831 59332
rect 420637 59331 420703 59332
rect 421741 59331 421807 59332
rect 425973 59331 426039 59332
rect 428181 59331 428247 59332
rect 453389 59331 453455 59332
rect 463509 59331 463575 59332
rect 148501 59260 148567 59261
rect 150893 59260 150959 59261
rect 295885 59260 295951 59261
rect 298461 59260 298527 59261
rect 303429 59260 303495 59261
rect 323301 59260 323367 59261
rect 485957 59260 486023 59261
rect 52126 59196 52132 59260
rect 52196 59258 52202 59260
rect 143574 59258 143580 59260
rect 52196 59198 143580 59258
rect 52196 59196 52202 59198
rect 143574 59196 143580 59198
rect 143644 59196 143650 59260
rect 148501 59256 148548 59260
rect 148612 59258 148618 59260
rect 148501 59200 148506 59256
rect 148501 59196 148548 59200
rect 148612 59198 148658 59258
rect 150893 59256 150940 59260
rect 151004 59258 151010 59260
rect 150893 59200 150898 59256
rect 148612 59196 148618 59198
rect 150893 59196 150940 59200
rect 151004 59198 151050 59258
rect 151004 59196 151010 59198
rect 202638 59196 202644 59260
rect 202708 59258 202714 59260
rect 285990 59258 285996 59260
rect 202708 59198 285996 59258
rect 202708 59196 202714 59198
rect 285990 59196 285996 59198
rect 286060 59196 286066 59260
rect 295885 59256 295932 59260
rect 295996 59258 296002 59260
rect 295885 59200 295890 59256
rect 295885 59196 295932 59200
rect 295996 59198 296042 59258
rect 298461 59256 298508 59260
rect 298572 59258 298578 59260
rect 298461 59200 298466 59256
rect 295996 59196 296002 59198
rect 298461 59196 298508 59200
rect 298572 59198 298618 59258
rect 303429 59256 303476 59260
rect 303540 59258 303546 59260
rect 303429 59200 303434 59256
rect 298572 59196 298578 59198
rect 303429 59196 303476 59200
rect 303540 59198 303586 59258
rect 323301 59256 323348 59260
rect 323412 59258 323418 59260
rect 323301 59200 323306 59256
rect 303540 59196 303546 59198
rect 323301 59196 323348 59200
rect 323412 59198 323458 59258
rect 323412 59196 323418 59198
rect 357934 59196 357940 59260
rect 358004 59258 358010 59260
rect 483422 59258 483428 59260
rect 358004 59198 483428 59258
rect 358004 59196 358010 59198
rect 483422 59196 483428 59198
rect 483492 59196 483498 59260
rect 485957 59256 486004 59260
rect 486068 59258 486074 59260
rect 485957 59200 485962 59256
rect 485957 59196 486004 59200
rect 486068 59198 486114 59258
rect 486068 59196 486074 59198
rect 148501 59195 148567 59196
rect 150893 59195 150959 59196
rect 295885 59195 295951 59196
rect 298461 59195 298527 59196
rect 303429 59195 303495 59196
rect 323301 59195 323367 59196
rect 485957 59195 486023 59196
rect 54886 59060 54892 59124
rect 54956 59122 54962 59124
rect 140814 59122 140820 59124
rect 54956 59062 140820 59122
rect 54956 59060 54962 59062
rect 140814 59060 140820 59062
rect 140884 59060 140890 59124
rect 198590 59060 198596 59124
rect 198660 59122 198666 59124
rect 280838 59122 280844 59124
rect 198660 59062 280844 59122
rect 198660 59060 198666 59062
rect 280838 59060 280844 59062
rect 280908 59060 280914 59124
rect 367686 59060 367692 59124
rect 367756 59122 367762 59124
rect 468518 59122 468524 59124
rect 367756 59062 468524 59122
rect 367756 59060 367762 59062
rect 468518 59060 468524 59062
rect 468588 59060 468594 59124
rect 53414 58924 53420 58988
rect 53484 58986 53490 58988
rect 138422 58986 138428 58988
rect 53484 58926 138428 58986
rect 53484 58924 53490 58926
rect 138422 58924 138428 58926
rect 138492 58924 138498 58988
rect 210734 58924 210740 58988
rect 210804 58986 210810 58988
rect 290958 58986 290964 58988
rect 210804 58926 290964 58986
rect 210804 58924 210810 58926
rect 290958 58924 290964 58926
rect 291028 58924 291034 58988
rect 374494 58924 374500 58988
rect 374564 58986 374570 58988
rect 473486 58986 473492 58988
rect 374564 58926 473492 58986
rect 374564 58924 374570 58926
rect 473486 58924 473492 58926
rect 473556 58924 473562 58988
rect 51942 58788 51948 58852
rect 52012 58850 52018 58852
rect 135846 58850 135852 58852
rect 52012 58790 135852 58850
rect 52012 58788 52018 58790
rect 135846 58788 135852 58790
rect 135916 58788 135922 58852
rect 201350 58788 201356 58852
rect 201420 58850 201426 58852
rect 273478 58850 273484 58852
rect 201420 58790 273484 58850
rect 201420 58788 201426 58790
rect 273478 58788 273484 58790
rect 273548 58788 273554 58852
rect 375966 58788 375972 58852
rect 376036 58850 376042 58852
rect 475878 58850 475884 58852
rect 376036 58790 475884 58850
rect 376036 58788 376042 58790
rect 475878 58788 475884 58790
rect 475948 58788 475954 58852
rect -960 58578 480 58668
rect 48078 58652 48084 58716
rect 48148 58714 48154 58716
rect 108246 58714 108252 58716
rect 48148 58654 108252 58714
rect 48148 58652 48154 58654
rect 108246 58652 108252 58654
rect 108316 58652 108322 58716
rect 209630 58652 209636 58716
rect 209700 58714 209706 58716
rect 276054 58714 276060 58716
rect 209700 58654 276060 58714
rect 209700 58652 209706 58654
rect 276054 58652 276060 58654
rect 276124 58652 276130 58716
rect 371734 58652 371740 58716
rect 371804 58714 371810 58716
rect 458398 58714 458404 58716
rect 371804 58654 458404 58714
rect 371804 58652 371810 58654
rect 458398 58652 458404 58654
rect 458468 58652 458474 58716
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 52310 58516 52316 58580
rect 52380 58578 52386 58580
rect 111006 58578 111012 58580
rect 52380 58518 111012 58578
rect 52380 58516 52386 58518
rect 111006 58516 111012 58518
rect 111076 58516 111082 58580
rect 202086 58516 202092 58580
rect 202156 58578 202162 58580
rect 268326 58578 268332 58580
rect 202156 58518 268332 58578
rect 202156 58516 202162 58518
rect 268326 58516 268332 58518
rect 268396 58516 268402 58580
rect 377990 58516 377996 58580
rect 378060 58578 378066 58580
rect 425278 58578 425284 58580
rect 378060 58518 425284 58578
rect 378060 58516 378066 58518
rect 425278 58516 425284 58518
rect 425348 58516 425354 58580
rect 59302 58380 59308 58444
rect 59372 58442 59378 58444
rect 101070 58442 101076 58444
rect 59372 58382 101076 58442
rect 59372 58380 59378 58382
rect 101070 58380 101076 58382
rect 101140 58380 101146 58444
rect 200614 58380 200620 58444
rect 200684 58442 200690 58444
rect 255998 58442 256004 58444
rect 200684 58382 256004 58442
rect 200684 58380 200690 58382
rect 255998 58380 256004 58382
rect 256068 58380 256074 58444
rect 377254 58380 377260 58444
rect 377324 58442 377330 58444
rect 419390 58442 419396 58444
rect 377324 58382 419396 58442
rect 377324 58380 377330 58382
rect 419390 58380 419396 58382
rect 419460 58380 419466 58444
rect 325877 58172 325943 58173
rect 85430 58108 85436 58172
rect 85500 58108 85506 58172
rect 92238 58108 92244 58172
rect 92308 58108 92314 58172
rect 128302 58108 128308 58172
rect 128372 58108 128378 58172
rect 153326 58108 153332 58172
rect 153396 58108 153402 58172
rect 235942 58108 235948 58172
rect 236012 58108 236018 58172
rect 272190 58108 272196 58172
rect 272260 58108 272266 58172
rect 275686 58108 275692 58172
rect 275756 58108 275762 58172
rect 300894 58108 300900 58172
rect 300964 58108 300970 58172
rect 325877 58168 325924 58172
rect 325988 58170 325994 58172
rect 325877 58112 325882 58168
rect 325877 58108 325924 58112
rect 325988 58110 326034 58170
rect 325988 58108 325994 58110
rect 398230 58108 398236 58172
rect 398300 58108 398306 58172
rect 401726 58108 401732 58172
rect 401796 58108 401802 58172
rect 405406 58108 405412 58172
rect 405476 58108 405482 58172
rect 416078 58108 416084 58172
rect 416148 58108 416154 58172
rect 83958 57972 83964 58036
rect 84028 58034 84034 58036
rect 84193 58034 84259 58037
rect 84028 58032 84259 58034
rect 84028 57976 84198 58032
rect 84254 57976 84259 58032
rect 84028 57974 84259 57976
rect 84028 57972 84034 57974
rect 84193 57971 84259 57974
rect 85438 57901 85498 58108
rect 76005 57900 76071 57901
rect 78213 57900 78279 57901
rect 79501 57900 79567 57901
rect 76005 57896 76052 57900
rect 76116 57898 76122 57900
rect 76005 57840 76010 57896
rect 76005 57836 76052 57840
rect 76116 57838 76162 57898
rect 78213 57896 78260 57900
rect 78324 57898 78330 57900
rect 78213 57840 78218 57896
rect 76116 57836 76122 57838
rect 78213 57836 78260 57840
rect 78324 57838 78370 57898
rect 79501 57896 79548 57900
rect 79612 57898 79618 57900
rect 80053 57898 80119 57901
rect 80462 57898 80468 57900
rect 79501 57840 79506 57896
rect 78324 57836 78330 57838
rect 79501 57836 79548 57840
rect 79612 57838 79658 57898
rect 80053 57896 80468 57898
rect 80053 57840 80058 57896
rect 80114 57840 80468 57896
rect 80053 57838 80468 57840
rect 79612 57836 79618 57838
rect 76005 57835 76071 57836
rect 78213 57835 78279 57836
rect 79501 57835 79567 57836
rect 80053 57835 80119 57838
rect 80462 57836 80468 57838
rect 80532 57836 80538 57900
rect 81801 57898 81867 57901
rect 81934 57898 81940 57900
rect 81801 57896 81940 57898
rect 81801 57840 81806 57896
rect 81862 57840 81940 57896
rect 81801 57838 81940 57840
rect 81801 57835 81867 57838
rect 81934 57836 81940 57838
rect 82004 57836 82010 57900
rect 85389 57896 85498 57901
rect 85389 57840 85394 57896
rect 85450 57840 85498 57896
rect 85389 57838 85498 57840
rect 86493 57900 86559 57901
rect 86493 57896 86540 57900
rect 86604 57898 86610 57900
rect 86953 57898 87019 57901
rect 88333 57900 88399 57901
rect 88701 57900 88767 57901
rect 87638 57898 87644 57900
rect 86493 57840 86498 57896
rect 85389 57835 85455 57838
rect 86493 57836 86540 57840
rect 86604 57838 86650 57898
rect 86953 57896 87644 57898
rect 86953 57840 86958 57896
rect 87014 57840 87644 57896
rect 86953 57838 87644 57840
rect 86604 57836 86610 57838
rect 86493 57835 86559 57836
rect 86953 57835 87019 57838
rect 87638 57836 87644 57838
rect 87708 57836 87714 57900
rect 88333 57896 88380 57900
rect 88444 57898 88450 57900
rect 88333 57840 88338 57896
rect 88333 57836 88380 57840
rect 88444 57838 88490 57898
rect 88701 57896 88748 57900
rect 88812 57898 88818 57900
rect 89713 57898 89779 57901
rect 90725 57900 90791 57901
rect 90030 57898 90036 57900
rect 88701 57840 88706 57896
rect 88444 57836 88450 57838
rect 88701 57836 88748 57840
rect 88812 57838 88858 57898
rect 89713 57896 90036 57898
rect 89713 57840 89718 57896
rect 89774 57840 90036 57896
rect 89713 57838 90036 57840
rect 88812 57836 88818 57838
rect 88333 57835 88399 57836
rect 88701 57835 88767 57836
rect 89713 57835 89779 57838
rect 90030 57836 90036 57838
rect 90100 57836 90106 57900
rect 90725 57896 90772 57900
rect 90836 57898 90842 57900
rect 91185 57898 91251 57901
rect 91318 57898 91324 57900
rect 90725 57840 90730 57896
rect 90725 57836 90772 57840
rect 90836 57838 90882 57898
rect 91185 57896 91324 57898
rect 91185 57840 91190 57896
rect 91246 57840 91324 57896
rect 91185 57838 91324 57840
rect 90836 57836 90842 57838
rect 90725 57835 90791 57836
rect 91185 57835 91251 57838
rect 91318 57836 91324 57838
rect 91388 57836 91394 57900
rect 92105 57898 92171 57901
rect 92246 57898 92306 58108
rect 128310 57901 128370 58108
rect 153334 57901 153394 58108
rect 235950 57901 236010 58108
rect 272198 57901 272258 58108
rect 92105 57896 92306 57898
rect 92105 57840 92110 57896
rect 92166 57840 92306 57896
rect 92105 57838 92306 57840
rect 92473 57898 92539 57901
rect 103789 57900 103855 57901
rect 93342 57898 93348 57900
rect 92473 57896 93348 57898
rect 92473 57840 92478 57896
rect 92534 57840 93348 57896
rect 92473 57838 93348 57840
rect 92105 57835 92171 57838
rect 92473 57835 92539 57838
rect 93342 57836 93348 57838
rect 93412 57836 93418 57900
rect 103789 57896 103836 57900
rect 103900 57898 103906 57900
rect 104985 57898 105051 57901
rect 106365 57900 106431 57901
rect 105302 57898 105308 57900
rect 103789 57840 103794 57896
rect 103789 57836 103836 57840
rect 103900 57838 103946 57898
rect 104985 57896 105308 57898
rect 104985 57840 104990 57896
rect 105046 57840 105308 57896
rect 104985 57838 105308 57840
rect 103900 57836 103906 57838
rect 103789 57835 103855 57836
rect 104985 57835 105051 57838
rect 105302 57836 105308 57838
rect 105372 57836 105378 57900
rect 106365 57896 106412 57900
rect 106476 57898 106482 57900
rect 106733 57898 106799 57901
rect 107510 57898 107516 57900
rect 106365 57840 106370 57896
rect 106365 57836 106412 57840
rect 106476 57838 106522 57898
rect 106733 57896 107516 57898
rect 106733 57840 106738 57896
rect 106794 57840 107516 57896
rect 106733 57838 107516 57840
rect 106476 57836 106482 57838
rect 106365 57835 106431 57836
rect 106733 57835 106799 57838
rect 107510 57836 107516 57838
rect 107580 57836 107586 57900
rect 108021 57898 108087 57901
rect 108614 57898 108620 57900
rect 108021 57896 108620 57898
rect 108021 57840 108026 57896
rect 108082 57840 108620 57896
rect 108021 57838 108620 57840
rect 108021 57835 108087 57838
rect 108614 57836 108620 57838
rect 108684 57836 108690 57900
rect 109217 57898 109283 57901
rect 111149 57900 111215 57901
rect 115749 57900 115815 57901
rect 123477 57900 123543 57901
rect 125869 57900 125935 57901
rect 109534 57898 109540 57900
rect 109217 57896 109540 57898
rect 109217 57840 109222 57896
rect 109278 57840 109540 57896
rect 109217 57838 109540 57840
rect 109217 57835 109283 57838
rect 109534 57836 109540 57838
rect 109604 57836 109610 57900
rect 111149 57896 111196 57900
rect 111260 57898 111266 57900
rect 111149 57840 111154 57896
rect 111149 57836 111196 57840
rect 111260 57838 111306 57898
rect 115749 57896 115796 57900
rect 115860 57898 115866 57900
rect 115749 57840 115754 57896
rect 111260 57836 111266 57838
rect 115749 57836 115796 57840
rect 115860 57838 115906 57898
rect 123477 57896 123524 57900
rect 123588 57898 123594 57900
rect 123477 57840 123482 57896
rect 115860 57836 115866 57838
rect 123477 57836 123524 57840
rect 123588 57838 123634 57898
rect 125869 57896 125916 57900
rect 125980 57898 125986 57900
rect 125869 57840 125874 57896
rect 123588 57836 123594 57838
rect 125869 57836 125916 57840
rect 125980 57838 126026 57898
rect 128310 57896 128419 57901
rect 128310 57840 128358 57896
rect 128414 57840 128419 57896
rect 128310 57838 128419 57840
rect 125980 57836 125986 57838
rect 111149 57835 111215 57836
rect 115749 57835 115815 57836
rect 123477 57835 123543 57836
rect 125869 57835 125935 57836
rect 128353 57835 128419 57838
rect 130837 57900 130903 57901
rect 133413 57900 133479 57901
rect 145557 57900 145623 57901
rect 130837 57896 130884 57900
rect 130948 57898 130954 57900
rect 130837 57840 130842 57896
rect 130837 57836 130884 57840
rect 130948 57838 130994 57898
rect 133413 57896 133460 57900
rect 133524 57898 133530 57900
rect 133413 57840 133418 57896
rect 130948 57836 130954 57838
rect 133413 57836 133460 57840
rect 133524 57838 133570 57898
rect 145557 57896 145604 57900
rect 145668 57898 145674 57900
rect 145557 57840 145562 57896
rect 133524 57836 133530 57838
rect 145557 57836 145604 57840
rect 145668 57838 145714 57898
rect 153285 57896 153394 57901
rect 153285 57840 153290 57896
rect 153346 57840 153394 57896
rect 153285 57838 153394 57840
rect 145668 57836 145674 57838
rect 130837 57835 130903 57836
rect 133413 57835 133479 57836
rect 145557 57835 145623 57836
rect 153285 57835 153351 57838
rect 183134 57836 183140 57900
rect 183204 57898 183210 57900
rect 183277 57898 183343 57901
rect 183204 57896 183343 57898
rect 183204 57840 183282 57896
rect 183338 57840 183343 57896
rect 183204 57838 183343 57840
rect 235950 57896 236059 57901
rect 235950 57840 235998 57896
rect 236054 57840 236059 57896
rect 235950 57838 236059 57840
rect 183204 57836 183210 57838
rect 183277 57835 183343 57838
rect 235993 57835 236059 57838
rect 237373 57898 237439 57901
rect 239213 57900 239279 57901
rect 242893 57900 242959 57901
rect 238150 57898 238156 57900
rect 237373 57896 238156 57898
rect 237373 57840 237378 57896
rect 237434 57840 238156 57896
rect 237373 57838 238156 57840
rect 237373 57835 237439 57838
rect 238150 57836 238156 57838
rect 238220 57836 238226 57900
rect 239213 57896 239260 57900
rect 239324 57898 239330 57900
rect 239213 57840 239218 57896
rect 239213 57836 239260 57840
rect 239324 57838 239370 57898
rect 242893 57896 242940 57900
rect 243004 57898 243010 57900
rect 244365 57898 244431 57901
rect 246389 57900 246455 57901
rect 248597 57900 248663 57901
rect 251173 57900 251239 57901
rect 253381 57900 253447 57901
rect 245326 57898 245332 57900
rect 242893 57840 242898 57896
rect 239324 57836 239330 57838
rect 242893 57836 242940 57840
rect 243004 57838 243050 57898
rect 244365 57896 245332 57898
rect 244365 57840 244370 57896
rect 244426 57840 245332 57896
rect 244365 57838 245332 57840
rect 243004 57836 243010 57838
rect 239213 57835 239279 57836
rect 242893 57835 242959 57836
rect 244365 57835 244431 57838
rect 245326 57836 245332 57838
rect 245396 57836 245402 57900
rect 246389 57896 246436 57900
rect 246500 57898 246506 57900
rect 246389 57840 246394 57896
rect 246389 57836 246436 57840
rect 246500 57838 246546 57898
rect 248597 57896 248644 57900
rect 248708 57898 248714 57900
rect 248597 57840 248602 57896
rect 246500 57836 246506 57838
rect 248597 57836 248644 57840
rect 248708 57838 248754 57898
rect 251173 57896 251220 57900
rect 251284 57898 251290 57900
rect 251173 57840 251178 57896
rect 248708 57836 248714 57838
rect 251173 57836 251220 57840
rect 251284 57838 251330 57898
rect 253381 57896 253428 57900
rect 253492 57898 253498 57900
rect 265341 57898 265407 57901
rect 266353 57900 266419 57901
rect 265934 57898 265940 57900
rect 253381 57840 253386 57896
rect 251284 57836 251290 57838
rect 253381 57836 253428 57840
rect 253492 57838 253538 57898
rect 265341 57896 265940 57898
rect 265341 57840 265346 57896
rect 265402 57840 265940 57896
rect 265341 57838 265940 57840
rect 253492 57836 253498 57838
rect 246389 57835 246455 57836
rect 248597 57835 248663 57836
rect 251173 57835 251239 57836
rect 253381 57835 253447 57836
rect 265341 57835 265407 57838
rect 265934 57836 265940 57838
rect 266004 57836 266010 57900
rect 266302 57898 266308 57900
rect 266262 57838 266308 57898
rect 266372 57896 266419 57900
rect 266414 57840 266419 57896
rect 266302 57836 266308 57838
rect 266372 57836 266419 57840
rect 266353 57835 266419 57836
rect 266997 57898 267063 57901
rect 269757 57900 269823 57901
rect 267590 57898 267596 57900
rect 266997 57896 267596 57898
rect 266997 57840 267002 57896
rect 267058 57840 267596 57896
rect 266997 57838 267596 57840
rect 266997 57835 267063 57838
rect 267590 57836 267596 57838
rect 267660 57836 267666 57900
rect 269757 57896 269804 57900
rect 269868 57898 269874 57900
rect 269757 57840 269762 57896
rect 269757 57836 269804 57840
rect 269868 57838 269914 57898
rect 272149 57896 272258 57901
rect 272149 57840 272154 57896
rect 272210 57840 272258 57896
rect 272149 57838 272258 57840
rect 273621 57898 273687 57901
rect 274398 57898 274404 57900
rect 273621 57896 274404 57898
rect 273621 57840 273626 57896
rect 273682 57840 274404 57896
rect 273621 57838 274404 57840
rect 269868 57836 269874 57838
rect 269757 57835 269823 57836
rect 272149 57835 272215 57838
rect 273621 57835 273687 57838
rect 274398 57836 274404 57838
rect 274468 57836 274474 57900
rect 274633 57898 274699 57901
rect 275694 57898 275754 58108
rect 300902 57901 300962 58108
rect 325877 58107 325943 58108
rect 279049 57900 279115 57901
rect 278998 57898 279004 57900
rect 274633 57896 275754 57898
rect 274633 57840 274638 57896
rect 274694 57840 275754 57896
rect 274633 57838 275754 57840
rect 278958 57838 279004 57898
rect 279068 57896 279115 57900
rect 279110 57840 279115 57896
rect 274633 57835 274699 57838
rect 278998 57836 279004 57838
rect 279068 57836 279115 57840
rect 279049 57835 279115 57836
rect 283649 57898 283715 57901
rect 283782 57898 283788 57900
rect 283649 57896 283788 57898
rect 283649 57840 283654 57896
rect 283710 57840 283788 57896
rect 283649 57838 283788 57840
rect 283649 57835 283715 57838
rect 283782 57836 283788 57838
rect 283852 57836 283858 57900
rect 287605 57898 287671 57901
rect 293309 57900 293375 57901
rect 288198 57898 288204 57900
rect 287605 57896 288204 57898
rect 287605 57840 287610 57896
rect 287666 57840 288204 57896
rect 287605 57838 288204 57840
rect 287605 57835 287671 57838
rect 288198 57836 288204 57838
rect 288268 57836 288274 57900
rect 293309 57896 293356 57900
rect 293420 57898 293426 57900
rect 293309 57840 293314 57896
rect 293309 57836 293356 57840
rect 293420 57838 293466 57898
rect 300853 57896 300962 57901
rect 300853 57840 300858 57896
rect 300914 57840 300962 57896
rect 300853 57838 300962 57840
rect 305821 57900 305887 57901
rect 310973 57900 311039 57901
rect 313365 57900 313431 57901
rect 318333 57900 318399 57901
rect 320909 57900 320975 57901
rect 343173 57900 343239 57901
rect 343449 57900 343515 57901
rect 305821 57896 305868 57900
rect 305932 57898 305938 57900
rect 305821 57840 305826 57896
rect 293420 57836 293426 57838
rect 293309 57835 293375 57836
rect 300853 57835 300919 57838
rect 305821 57836 305868 57840
rect 305932 57838 305978 57898
rect 310973 57896 311020 57900
rect 311084 57898 311090 57900
rect 310973 57840 310978 57896
rect 305932 57836 305938 57838
rect 310973 57836 311020 57840
rect 311084 57838 311130 57898
rect 313365 57896 313412 57900
rect 313476 57898 313482 57900
rect 313365 57840 313370 57896
rect 311084 57836 311090 57838
rect 313365 57836 313412 57840
rect 313476 57838 313522 57898
rect 318333 57896 318380 57900
rect 318444 57898 318450 57900
rect 318333 57840 318338 57896
rect 313476 57836 313482 57838
rect 318333 57836 318380 57840
rect 318444 57838 318490 57898
rect 320909 57896 320956 57900
rect 321020 57898 321026 57900
rect 343173 57898 343220 57900
rect 320909 57840 320914 57896
rect 318444 57836 318450 57838
rect 320909 57836 320956 57840
rect 321020 57838 321066 57898
rect 343128 57896 343220 57898
rect 343128 57840 343178 57896
rect 343128 57838 343220 57840
rect 321020 57836 321026 57838
rect 343173 57836 343220 57838
rect 343284 57836 343290 57900
rect 343398 57898 343404 57900
rect 343358 57838 343404 57898
rect 343468 57896 343515 57900
rect 343510 57840 343515 57896
rect 343398 57836 343404 57838
rect 343468 57836 343515 57840
rect 305821 57835 305887 57836
rect 310973 57835 311039 57836
rect 313365 57835 313431 57836
rect 318333 57835 318399 57836
rect 320909 57835 320975 57836
rect 343173 57835 343239 57836
rect 343449 57835 343515 57836
rect 397453 57898 397519 57901
rect 398238 57898 398298 58108
rect 401734 57901 401794 58108
rect 397453 57896 398298 57898
rect 397453 57840 397458 57896
rect 397514 57840 398298 57896
rect 397453 57838 398298 57840
rect 399477 57900 399543 57901
rect 399477 57896 399524 57900
rect 399588 57898 399594 57900
rect 400213 57898 400279 57901
rect 400438 57898 400444 57900
rect 399477 57840 399482 57896
rect 397453 57835 397519 57838
rect 399477 57836 399524 57840
rect 399588 57838 399634 57898
rect 400213 57896 400444 57898
rect 400213 57840 400218 57896
rect 400274 57840 400444 57896
rect 400213 57838 400444 57840
rect 399588 57836 399594 57838
rect 399477 57835 399543 57836
rect 400213 57835 400279 57838
rect 400438 57836 400444 57838
rect 400508 57836 400514 57900
rect 401685 57896 401794 57901
rect 401685 57840 401690 57896
rect 401746 57840 401794 57896
rect 401685 57838 401794 57840
rect 404353 57898 404419 57901
rect 405414 57898 405474 58108
rect 416086 57901 416146 58108
rect 404353 57896 405474 57898
rect 404353 57840 404358 57896
rect 404414 57840 405474 57896
rect 404353 57838 405474 57840
rect 405825 57898 405891 57901
rect 406510 57898 406516 57900
rect 405825 57896 406516 57898
rect 405825 57840 405830 57896
rect 405886 57840 406516 57896
rect 405825 57838 406516 57840
rect 401685 57835 401751 57838
rect 404353 57835 404419 57838
rect 405825 57835 405891 57838
rect 406510 57836 406516 57838
rect 406580 57836 406586 57900
rect 407205 57898 407271 57901
rect 408309 57900 408375 57901
rect 408677 57900 408743 57901
rect 407614 57898 407620 57900
rect 407205 57896 407620 57898
rect 407205 57840 407210 57896
rect 407266 57840 407620 57896
rect 407205 57838 407620 57840
rect 407205 57835 407271 57838
rect 407614 57836 407620 57838
rect 407684 57836 407690 57900
rect 408309 57896 408356 57900
rect 408420 57898 408426 57900
rect 408309 57840 408314 57896
rect 408309 57836 408356 57840
rect 408420 57838 408466 57898
rect 408677 57896 408724 57900
rect 408788 57898 408794 57900
rect 409873 57898 409939 57901
rect 410006 57898 410012 57900
rect 408677 57840 408682 57896
rect 408420 57836 408426 57838
rect 408677 57836 408724 57840
rect 408788 57838 408834 57898
rect 409873 57896 410012 57898
rect 409873 57840 409878 57896
rect 409934 57840 410012 57896
rect 409873 57838 410012 57840
rect 408788 57836 408794 57838
rect 408309 57835 408375 57836
rect 408677 57835 408743 57836
rect 409873 57835 409939 57838
rect 410006 57836 410012 57838
rect 410076 57836 410082 57900
rect 411345 57898 411411 57901
rect 414565 57900 414631 57901
rect 415485 57900 415551 57901
rect 412398 57898 412404 57900
rect 411345 57896 412404 57898
rect 411345 57840 411350 57896
rect 411406 57840 412404 57896
rect 411345 57838 412404 57840
rect 411345 57835 411411 57838
rect 412398 57836 412404 57838
rect 412468 57836 412474 57900
rect 414565 57896 414612 57900
rect 414676 57898 414682 57900
rect 414565 57840 414570 57896
rect 414565 57836 414612 57840
rect 414676 57838 414722 57898
rect 415485 57896 415532 57900
rect 415596 57898 415602 57900
rect 415485 57840 415490 57896
rect 414676 57836 414682 57838
rect 415485 57836 415532 57840
rect 415596 57838 415642 57898
rect 416037 57896 416146 57901
rect 426433 57900 426499 57901
rect 426382 57898 426388 57900
rect 416037 57840 416042 57896
rect 416098 57840 416146 57896
rect 416037 57838 416146 57840
rect 426342 57838 426388 57898
rect 426452 57896 426499 57900
rect 427629 57900 427695 57901
rect 427629 57898 427676 57900
rect 426494 57840 426499 57896
rect 415596 57836 415602 57838
rect 414565 57835 414631 57836
rect 415485 57835 415551 57836
rect 416037 57835 416103 57838
rect 426382 57836 426388 57838
rect 426452 57836 426499 57840
rect 427584 57896 427676 57898
rect 427584 57840 427634 57896
rect 427584 57838 427676 57840
rect 426433 57835 426499 57836
rect 427629 57836 427676 57838
rect 427740 57836 427746 57900
rect 427813 57898 427879 57901
rect 428590 57898 428596 57900
rect 427813 57896 428596 57898
rect 427813 57840 427818 57896
rect 427874 57840 428596 57896
rect 427813 57838 428596 57840
rect 427629 57835 427695 57836
rect 427813 57835 427879 57838
rect 428590 57836 428596 57838
rect 428660 57836 428666 57900
rect 429193 57898 429259 57901
rect 429694 57898 429700 57900
rect 429193 57896 429700 57898
rect 429193 57840 429198 57896
rect 429254 57840 429700 57896
rect 429193 57838 429700 57840
rect 429193 57835 429259 57838
rect 429694 57836 429700 57838
rect 429764 57836 429770 57900
rect 430573 57898 430639 57901
rect 432229 57900 432295 57901
rect 433333 57900 433399 57901
rect 433609 57900 433675 57901
rect 431166 57898 431172 57900
rect 430573 57896 431172 57898
rect 430573 57840 430578 57896
rect 430634 57840 431172 57896
rect 430573 57838 431172 57840
rect 430573 57835 430639 57838
rect 431166 57836 431172 57838
rect 431236 57836 431242 57900
rect 432229 57896 432276 57900
rect 432340 57898 432346 57900
rect 432229 57840 432234 57896
rect 432229 57836 432276 57840
rect 432340 57838 432386 57898
rect 433333 57896 433380 57900
rect 433444 57898 433450 57900
rect 433333 57840 433338 57896
rect 432340 57836 432346 57838
rect 433333 57836 433380 57840
rect 433444 57838 433490 57898
rect 433444 57836 433450 57838
rect 433558 57836 433564 57900
rect 433628 57898 433675 57900
rect 435909 57900 435975 57901
rect 435909 57898 435956 57900
rect 433628 57896 433720 57898
rect 433670 57840 433720 57896
rect 433628 57838 433720 57840
rect 435864 57896 435956 57898
rect 435864 57840 435914 57896
rect 435864 57838 435956 57840
rect 433628 57836 433675 57838
rect 432229 57835 432295 57836
rect 433333 57835 433399 57836
rect 433609 57835 433675 57836
rect 435909 57836 435956 57838
rect 436020 57836 436026 57900
rect 436093 57898 436159 57901
rect 436870 57898 436876 57900
rect 436093 57896 436876 57898
rect 436093 57840 436098 57896
rect 436154 57840 436876 57896
rect 436093 57838 436876 57840
rect 435909 57835 435975 57836
rect 436093 57835 436159 57838
rect 436870 57836 436876 57838
rect 436940 57836 436946 57900
rect 438209 57898 438275 57901
rect 438485 57900 438551 57901
rect 438342 57898 438348 57900
rect 438209 57896 438348 57898
rect 438209 57840 438214 57896
rect 438270 57840 438348 57896
rect 438209 57838 438348 57840
rect 438209 57835 438275 57838
rect 438342 57836 438348 57838
rect 438412 57836 438418 57900
rect 438485 57896 438532 57900
rect 438596 57898 438602 57900
rect 438853 57898 438919 57901
rect 440877 57900 440943 57901
rect 443453 57900 443519 57901
rect 448237 57900 448303 57901
rect 470869 57900 470935 57901
rect 478413 57900 478479 57901
rect 439078 57898 439084 57900
rect 438485 57840 438490 57896
rect 438485 57836 438532 57840
rect 438596 57838 438642 57898
rect 438853 57896 439084 57898
rect 438853 57840 438858 57896
rect 438914 57840 439084 57896
rect 438853 57838 439084 57840
rect 438596 57836 438602 57838
rect 438485 57835 438551 57836
rect 438853 57835 438919 57838
rect 439078 57836 439084 57838
rect 439148 57836 439154 57900
rect 440877 57896 440924 57900
rect 440988 57898 440994 57900
rect 440877 57840 440882 57896
rect 440877 57836 440924 57840
rect 440988 57838 441034 57898
rect 443453 57896 443500 57900
rect 443564 57898 443570 57900
rect 443453 57840 443458 57896
rect 440988 57836 440994 57838
rect 443453 57836 443500 57840
rect 443564 57838 443610 57898
rect 448237 57896 448284 57900
rect 448348 57898 448354 57900
rect 448237 57840 448242 57896
rect 443564 57836 443570 57838
rect 448237 57836 448284 57840
rect 448348 57838 448394 57898
rect 470869 57896 470916 57900
rect 470980 57898 470986 57900
rect 470869 57840 470874 57896
rect 448348 57836 448354 57838
rect 470869 57836 470916 57840
rect 470980 57838 471026 57898
rect 478413 57896 478460 57900
rect 478524 57898 478530 57900
rect 478413 57840 478418 57896
rect 470980 57836 470986 57838
rect 478413 57836 478460 57840
rect 478524 57838 478570 57898
rect 478524 57836 478530 57838
rect 503110 57836 503116 57900
rect 503180 57898 503186 57900
rect 503253 57898 503319 57901
rect 503529 57900 503595 57901
rect 503180 57896 503319 57898
rect 503180 57840 503258 57896
rect 503314 57840 503319 57896
rect 503180 57838 503319 57840
rect 503180 57836 503186 57838
rect 440877 57835 440943 57836
rect 443453 57835 443519 57836
rect 448237 57835 448303 57836
rect 470869 57835 470935 57836
rect 478413 57835 478479 57836
rect 503253 57835 503319 57838
rect 503478 57836 503484 57900
rect 503548 57898 503595 57900
rect 503548 57896 503640 57898
rect 503590 57840 503640 57896
rect 503548 57838 503640 57840
rect 503548 57836 503595 57838
rect 503529 57835 503595 57836
rect 183461 57764 183527 57765
rect 57646 57700 57652 57764
rect 57716 57762 57722 57764
rect 117998 57762 118004 57764
rect 57716 57702 98746 57762
rect 57716 57700 57722 57702
rect 44950 57564 44956 57628
rect 45020 57626 45026 57628
rect 98494 57626 98500 57628
rect 45020 57566 98500 57626
rect 45020 57564 45026 57566
rect 98494 57564 98500 57566
rect 98564 57564 98570 57628
rect 98686 57626 98746 57702
rect 103470 57702 118004 57762
rect 103470 57626 103530 57702
rect 117998 57700 118004 57702
rect 118068 57700 118074 57764
rect 183461 57760 183508 57764
rect 183572 57762 183578 57764
rect 183461 57704 183466 57760
rect 183461 57700 183508 57704
rect 183572 57702 183618 57762
rect 183572 57700 183578 57702
rect 211654 57700 211660 57764
rect 211724 57762 211730 57764
rect 270902 57762 270908 57764
rect 211724 57702 270908 57762
rect 211724 57700 211730 57702
rect 270902 57700 270908 57702
rect 270972 57700 270978 57764
rect 358118 57700 358124 57764
rect 358188 57762 358194 57764
rect 451038 57762 451044 57764
rect 358188 57702 451044 57762
rect 358188 57700 358194 57702
rect 451038 57700 451044 57702
rect 451108 57700 451114 57764
rect 183461 57699 183527 57700
rect 98686 57566 103530 57626
rect 111793 57626 111859 57629
rect 112110 57626 112116 57628
rect 111793 57624 112116 57626
rect 111793 57568 111798 57624
rect 111854 57568 112116 57624
rect 111793 57566 112116 57568
rect 111793 57563 111859 57566
rect 112110 57564 112116 57566
rect 112180 57564 112186 57628
rect 113173 57626 113239 57629
rect 115933 57628 115999 57629
rect 114318 57626 114324 57628
rect 113173 57624 114324 57626
rect 113173 57568 113178 57624
rect 113234 57568 114324 57624
rect 113173 57566 114324 57568
rect 113173 57563 113239 57566
rect 114318 57564 114324 57566
rect 114388 57564 114394 57628
rect 115933 57624 115980 57628
rect 116044 57626 116050 57628
rect 118693 57626 118759 57629
rect 155953 57628 156019 57629
rect 119102 57626 119108 57628
rect 115933 57568 115938 57624
rect 115933 57564 115980 57568
rect 116044 57566 116090 57626
rect 118693 57624 119108 57626
rect 118693 57568 118698 57624
rect 118754 57568 119108 57624
rect 118693 57566 119108 57568
rect 116044 57564 116050 57566
rect 115933 57563 115999 57564
rect 118693 57563 118759 57566
rect 119102 57564 119108 57566
rect 119172 57564 119178 57628
rect 155902 57626 155908 57628
rect 155862 57566 155908 57626
rect 155972 57624 156019 57628
rect 156014 57568 156019 57624
rect 155902 57564 155908 57566
rect 155972 57564 156019 57568
rect 155953 57563 156019 57564
rect 160093 57626 160159 57629
rect 160870 57626 160876 57628
rect 160093 57624 160876 57626
rect 160093 57568 160098 57624
rect 160154 57568 160876 57624
rect 160093 57566 160876 57568
rect 160093 57563 160159 57566
rect 160870 57564 160876 57566
rect 160940 57564 160946 57628
rect 165613 57626 165679 57629
rect 165838 57626 165844 57628
rect 165613 57624 165844 57626
rect 165613 57568 165618 57624
rect 165674 57568 165844 57624
rect 165613 57566 165844 57568
rect 165613 57563 165679 57566
rect 165838 57564 165844 57566
rect 165908 57564 165914 57628
rect 204846 57564 204852 57628
rect 204916 57626 204922 57628
rect 260966 57626 260972 57628
rect 204916 57566 260972 57626
rect 204916 57564 204922 57566
rect 260966 57564 260972 57566
rect 261036 57564 261042 57628
rect 267733 57626 267799 57629
rect 268694 57626 268700 57628
rect 267733 57624 268700 57626
rect 267733 57568 267738 57624
rect 267794 57568 268700 57624
rect 267733 57566 268700 57568
rect 267733 57563 267799 57566
rect 268694 57564 268700 57566
rect 268764 57564 268770 57628
rect 270493 57626 270559 57629
rect 273345 57628 273411 57629
rect 271086 57626 271092 57628
rect 270493 57624 271092 57626
rect 270493 57568 270498 57624
rect 270554 57568 271092 57624
rect 270493 57566 271092 57568
rect 270493 57563 270559 57566
rect 271086 57564 271092 57566
rect 271156 57564 271162 57628
rect 273294 57626 273300 57628
rect 273254 57566 273300 57626
rect 273364 57624 273411 57628
rect 273406 57568 273411 57624
rect 273294 57564 273300 57566
rect 273364 57564 273411 57568
rect 273345 57563 273411 57564
rect 277393 57626 277459 57629
rect 278078 57626 278084 57628
rect 277393 57624 278084 57626
rect 277393 57568 277398 57624
rect 277454 57568 278084 57624
rect 277393 57566 278084 57568
rect 277393 57563 277459 57566
rect 278078 57564 278084 57566
rect 278148 57564 278154 57628
rect 307753 57626 307819 57629
rect 308622 57626 308628 57628
rect 307753 57624 308628 57626
rect 307753 57568 307758 57624
rect 307814 57568 308628 57624
rect 307753 57566 308628 57568
rect 307753 57563 307819 57566
rect 308622 57564 308628 57566
rect 308692 57564 308698 57628
rect 376150 57564 376156 57628
rect 376220 57626 376226 57628
rect 460974 57626 460980 57628
rect 376220 57566 460980 57626
rect 376220 57564 376226 57566
rect 460974 57564 460980 57566
rect 461044 57564 461050 57628
rect 58750 57428 58756 57492
rect 58820 57490 58826 57492
rect 103830 57490 103836 57492
rect 58820 57430 103836 57490
rect 58820 57428 58826 57430
rect 103830 57428 103836 57430
rect 103900 57428 103906 57492
rect 214414 57428 214420 57492
rect 214484 57490 214490 57492
rect 240133 57490 240199 57493
rect 240542 57490 240548 57492
rect 214484 57430 240058 57490
rect 214484 57428 214490 57430
rect 57094 57292 57100 57356
rect 57164 57354 57170 57356
rect 97022 57354 97028 57356
rect 57164 57294 97028 57354
rect 57164 57292 57170 57294
rect 97022 57292 97028 57294
rect 97092 57292 97098 57356
rect 205030 57292 205036 57356
rect 205100 57354 205106 57356
rect 239857 57354 239923 57357
rect 205100 57352 239923 57354
rect 205100 57296 239862 57352
rect 239918 57296 239923 57352
rect 205100 57294 239923 57296
rect 239998 57354 240058 57430
rect 240133 57488 240548 57490
rect 240133 57432 240138 57488
rect 240194 57432 240548 57488
rect 240133 57430 240548 57432
rect 240133 57427 240199 57430
rect 240542 57428 240548 57430
rect 240612 57428 240618 57492
rect 241513 57490 241579 57493
rect 244273 57492 244339 57493
rect 241646 57490 241652 57492
rect 241513 57488 241652 57490
rect 241513 57432 241518 57488
rect 241574 57432 241652 57488
rect 241513 57430 241652 57432
rect 241513 57427 241579 57430
rect 241646 57428 241652 57430
rect 241716 57428 241722 57492
rect 244222 57490 244228 57492
rect 244182 57430 244228 57490
rect 244292 57488 244339 57492
rect 244334 57432 244339 57488
rect 244222 57428 244228 57430
rect 244292 57428 244339 57432
rect 244273 57427 244339 57428
rect 247033 57490 247099 57493
rect 247718 57490 247724 57492
rect 247033 57488 247724 57490
rect 247033 57432 247038 57488
rect 247094 57432 247724 57488
rect 247033 57430 247724 57432
rect 247033 57427 247099 57430
rect 247718 57428 247724 57430
rect 247788 57428 247794 57492
rect 249793 57490 249859 57493
rect 250110 57490 250116 57492
rect 249793 57488 250116 57490
rect 249793 57432 249798 57488
rect 249854 57432 250116 57488
rect 249793 57430 250116 57432
rect 249793 57427 249859 57430
rect 250110 57428 250116 57430
rect 250180 57428 250186 57492
rect 251357 57490 251423 57493
rect 252318 57490 252324 57492
rect 251357 57488 252324 57490
rect 251357 57432 251362 57488
rect 251418 57432 252324 57488
rect 251357 57430 252324 57432
rect 251357 57427 251423 57430
rect 252318 57428 252324 57430
rect 252388 57428 252394 57492
rect 253933 57490 253999 57493
rect 254526 57490 254532 57492
rect 253933 57488 254532 57490
rect 253933 57432 253938 57488
rect 253994 57432 254532 57488
rect 253933 57430 254532 57432
rect 253933 57427 253999 57430
rect 254526 57428 254532 57430
rect 254596 57428 254602 57492
rect 364926 57428 364932 57492
rect 364996 57490 365002 57492
rect 445886 57490 445892 57492
rect 364996 57430 445892 57490
rect 364996 57428 365002 57430
rect 445886 57428 445892 57430
rect 445956 57428 445962 57492
rect 258390 57354 258396 57356
rect 239998 57294 258396 57354
rect 205100 57292 205106 57294
rect 239857 57291 239923 57294
rect 258390 57292 258396 57294
rect 258460 57292 258466 57356
rect 378910 57292 378916 57356
rect 378980 57354 378986 57356
rect 456374 57354 456380 57356
rect 378980 57294 456380 57354
rect 378980 57292 378986 57294
rect 456374 57292 456380 57294
rect 456444 57292 456450 57356
rect 430941 57220 431007 57221
rect 59118 57156 59124 57220
rect 59188 57218 59194 57220
rect 96286 57218 96292 57220
rect 59188 57158 96292 57218
rect 59188 57156 59194 57158
rect 96286 57156 96292 57158
rect 96356 57156 96362 57220
rect 215886 57156 215892 57220
rect 215956 57218 215962 57220
rect 253606 57218 253612 57220
rect 215956 57158 253612 57218
rect 215956 57156 215962 57158
rect 253606 57156 253612 57158
rect 253676 57156 253682 57220
rect 379094 57156 379100 57220
rect 379164 57218 379170 57220
rect 421046 57218 421052 57220
rect 379164 57158 421052 57218
rect 379164 57156 379170 57158
rect 421046 57156 421052 57158
rect 421116 57156 421122 57220
rect 430941 57216 430988 57220
rect 431052 57218 431058 57220
rect 433425 57218 433491 57221
rect 435725 57220 435791 57221
rect 434662 57218 434668 57220
rect 430941 57160 430946 57216
rect 430941 57156 430988 57160
rect 431052 57158 431098 57218
rect 433425 57216 434668 57218
rect 433425 57160 433430 57216
rect 433486 57160 434668 57216
rect 433425 57158 434668 57160
rect 431052 57156 431058 57158
rect 430941 57155 431007 57156
rect 433425 57155 433491 57158
rect 434662 57156 434668 57158
rect 434732 57156 434738 57220
rect 435725 57216 435772 57220
rect 435836 57218 435842 57220
rect 435725 57160 435730 57216
rect 435725 57156 435772 57160
rect 435836 57158 435882 57218
rect 435836 57156 435842 57158
rect 435725 57155 435791 57156
rect 58934 57020 58940 57084
rect 59004 57082 59010 57084
rect 93710 57082 93716 57084
rect 59004 57022 93716 57082
rect 59004 57020 59010 57022
rect 93710 57020 93716 57022
rect 93780 57020 93786 57084
rect 214598 57020 214604 57084
rect 214668 57082 214674 57084
rect 250662 57082 250668 57084
rect 214668 57022 250668 57082
rect 214668 57020 214674 57022
rect 250662 57020 250668 57022
rect 250732 57020 250738 57084
rect 378726 57020 378732 57084
rect 378796 57082 378802 57084
rect 413502 57082 413508 57084
rect 378796 57022 413508 57082
rect 378796 57020 378802 57022
rect 413502 57020 413508 57022
rect 413572 57020 413578 57084
rect 239857 56946 239923 56949
rect 411253 56948 411319 56949
rect 248270 56946 248276 56948
rect 239857 56944 248276 56946
rect 239857 56888 239862 56944
rect 239918 56888 248276 56944
rect 239857 56886 248276 56888
rect 239857 56883 239923 56886
rect 248270 56884 248276 56886
rect 248340 56884 248346 56948
rect 411253 56944 411300 56948
rect 411364 56946 411370 56948
rect 412541 56946 412607 56949
rect 411253 56888 411258 56944
rect 411253 56884 411300 56888
rect 411364 56886 411410 56946
rect 412541 56944 412650 56946
rect 412541 56888 412546 56944
rect 412602 56888 412650 56944
rect 411364 56884 411370 56886
rect 411253 56883 411319 56884
rect 412541 56883 412650 56888
rect 412590 56813 412650 56883
rect 278446 56810 278452 56812
rect 258030 56750 278452 56810
rect 55070 56612 55076 56676
rect 55140 56674 55146 56676
rect 118366 56674 118372 56676
rect 55140 56614 118372 56674
rect 55140 56612 55146 56614
rect 118366 56612 118372 56614
rect 118436 56612 118442 56676
rect 163262 56612 163268 56676
rect 163332 56612 163338 56676
rect 202270 56612 202276 56676
rect 202340 56674 202346 56676
rect 258030 56674 258090 56750
rect 278446 56748 278452 56750
rect 278516 56748 278522 56812
rect 412590 56808 412699 56813
rect 412590 56752 412638 56808
rect 412694 56752 412699 56808
rect 412590 56750 412699 56752
rect 412633 56747 412699 56750
rect 202340 56614 258090 56674
rect 202340 56612 202346 56614
rect 370446 56612 370452 56676
rect 370516 56674 370522 56676
rect 465942 56674 465948 56676
rect 370516 56614 465948 56674
rect 370516 56612 370522 56614
rect 465942 56612 465948 56614
rect 466012 56612 466018 56676
rect 53598 56476 53604 56540
rect 53668 56538 53674 56540
rect 163270 56538 163330 56612
rect 53668 56478 163330 56538
rect 53668 56476 53674 56478
rect 219934 56476 219940 56540
rect 220004 56538 220010 56540
rect 410742 56538 410748 56540
rect 220004 56478 410748 56538
rect 220004 56476 220010 56478
rect 410742 56476 410748 56478
rect 410812 56476 410818 56540
rect 48630 56340 48636 56404
rect 48700 56402 48706 56404
rect 158478 56402 158484 56404
rect 48700 56342 158484 56402
rect 48700 56340 48706 56342
rect 158478 56340 158484 56342
rect 158548 56340 158554 56404
rect 217174 56340 217180 56404
rect 217244 56402 217250 56404
rect 276974 56402 276980 56404
rect 217244 56342 276980 56402
rect 217244 56340 217250 56342
rect 276974 56340 276980 56342
rect 277044 56340 277050 56404
rect 55622 56204 55628 56268
rect 55692 56266 55698 56268
rect 153285 56266 153351 56269
rect 55692 56264 153351 56266
rect 55692 56208 153290 56264
rect 153346 56208 153351 56264
rect 55692 56206 153351 56208
rect 55692 56204 55698 56206
rect 153285 56203 153351 56206
rect 50470 55116 50476 55180
rect 50540 55178 50546 55180
rect 165613 55178 165679 55181
rect 50540 55176 165679 55178
rect 50540 55120 165618 55176
rect 165674 55120 165679 55176
rect 50540 55118 165679 55120
rect 50540 55116 50546 55118
rect 165613 55115 165679 55118
rect 205214 55116 205220 55180
rect 205284 55178 205290 55180
rect 307753 55178 307819 55181
rect 205284 55176 307819 55178
rect 205284 55120 307758 55176
rect 307814 55120 307819 55176
rect 205284 55118 307819 55120
rect 205284 55116 205290 55118
rect 307753 55115 307819 55118
rect 377438 55116 377444 55180
rect 377508 55178 377514 55180
rect 438853 55178 438919 55181
rect 377508 55176 438919 55178
rect 377508 55120 438858 55176
rect 438914 55120 438919 55176
rect 377508 55118 438919 55120
rect 377508 55116 377514 55118
rect 438853 55115 438919 55118
rect 50654 54980 50660 55044
rect 50724 55042 50730 55044
rect 160093 55042 160159 55045
rect 50724 55040 160159 55042
rect 50724 54984 160098 55040
rect 160154 54984 160159 55040
rect 50724 54982 160159 54984
rect 50724 54980 50730 54982
rect 160093 54979 160159 54982
rect 217358 54980 217364 55044
rect 217428 55042 217434 55044
rect 277393 55042 277459 55045
rect 217428 55040 277459 55042
rect 217428 54984 277398 55040
rect 277454 54984 277459 55040
rect 217428 54982 277459 54984
rect 217428 54980 217434 54982
rect 277393 54979 277459 54982
rect 50838 54844 50844 54908
rect 50908 54906 50914 54908
rect 155953 54906 156019 54909
rect 50908 54904 156019 54906
rect 50908 54848 155958 54904
rect 156014 54848 156019 54904
rect 50908 54846 156019 54848
rect 50908 54844 50914 54846
rect 155953 54843 156019 54846
rect 217542 54844 217548 54908
rect 217612 54906 217618 54908
rect 249793 54906 249859 54909
rect 217612 54904 249859 54906
rect 217612 54848 249798 54904
rect 249854 54848 249859 54904
rect 217612 54846 249859 54848
rect 217612 54844 217618 54846
rect 249793 54843 249859 54846
rect 57462 54708 57468 54772
rect 57532 54770 57538 54772
rect 118693 54770 118759 54773
rect 57532 54768 118759 54770
rect 57532 54712 118698 54768
rect 118754 54712 118759 54768
rect 57532 54710 118759 54712
rect 57532 54708 57538 54710
rect 118693 54707 118759 54710
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19410 480 19500
rect 2773 19410 2839 19413
rect -960 19408 2839 19410
rect -960 19352 2778 19408
rect 2834 19352 2839 19408
rect -960 19350 2839 19352
rect -960 19260 480 19350
rect 2773 19347 2839 19350
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< via3 >>
rect 53052 630804 53116 630868
rect 54340 630668 54404 630732
rect 120028 625228 120092 625292
rect 430620 597620 430684 597684
rect 430804 592180 430868 592244
rect 120028 559540 120092 559604
rect 300164 543084 300228 543148
rect 299980 542676 300044 542740
rect 320588 541044 320652 541108
rect 300164 520100 300228 520164
rect 430620 518740 430684 518804
rect 320772 518604 320836 518668
rect 299980 517244 300044 517308
rect 430804 517244 430868 517308
rect 360700 485012 360764 485076
rect 59308 478756 59372 478820
rect 202460 478756 202524 478820
rect 357940 478756 358004 478820
rect 46796 478620 46860 478684
rect 198044 478620 198108 478684
rect 211844 478620 211908 478684
rect 360148 478620 360212 478684
rect 53236 478484 53300 478548
rect 196572 478484 196636 478548
rect 201356 478484 201420 478548
rect 206692 478484 206756 478548
rect 367692 478484 367756 478548
rect 197860 478348 197924 478412
rect 202644 478348 202708 478412
rect 371740 478348 371804 478412
rect 57652 478212 57716 478276
rect 202092 478212 202156 478276
rect 210740 478212 210804 478276
rect 219204 478212 219268 478276
rect 374500 478212 374564 478276
rect 200620 478076 200684 478140
rect 375972 478076 376036 478140
rect 54708 477940 54772 478004
rect 50660 477728 50724 477732
rect 50660 477672 50710 477728
rect 50710 477672 50724 477728
rect 50660 477668 50724 477672
rect 198228 477940 198292 478004
rect 209636 477940 209700 478004
rect 198596 477804 198660 477868
rect 199332 477668 199396 477732
rect 206508 477668 206572 477732
rect 50844 477592 50908 477596
rect 50844 477536 50894 477592
rect 50894 477536 50908 477592
rect 50844 477532 50908 477536
rect 200988 477532 201052 477596
rect 216996 477592 217060 477596
rect 216996 477536 217010 477592
rect 217010 477536 217060 477592
rect 216996 477532 217060 477536
rect 217364 477592 217428 477596
rect 217364 477536 217414 477592
rect 217414 477536 217428 477592
rect 217364 477532 217428 477536
rect 217548 477532 217612 477596
rect 219940 477532 220004 477596
rect 208348 476716 208412 476780
rect 377260 476716 377324 476780
rect 57284 475764 57348 475828
rect 211660 475628 211724 475692
rect 214420 475492 214484 475556
rect 47900 475356 47964 475420
rect 214604 475356 214668 475420
rect 378732 475356 378796 475420
rect 204852 474268 204916 474332
rect 205036 474132 205100 474196
rect 215340 473996 215404 474060
rect 378180 473996 378244 474060
rect 208900 472772 208964 472836
rect 358124 472772 358188 472836
rect 214788 472636 214852 472700
rect 370452 472636 370516 472700
rect 218836 472500 218900 472564
rect 376156 472500 376220 472564
rect 202276 471548 202340 471612
rect 214972 471412 215036 471476
rect 215892 471276 215956 471340
rect 359596 471276 359660 471340
rect 199148 471140 199212 471204
rect 378916 471140 378980 471204
rect 209820 469916 209884 469980
rect 377444 469916 377508 469980
rect 212764 469780 212828 469844
rect 379100 469780 379164 469844
rect 359412 468692 359476 468756
rect 212580 468556 212644 468620
rect 379468 468556 379532 468620
rect 196756 468420 196820 468484
rect 362908 468420 362972 468484
rect 203196 467196 203260 467260
rect 207060 467060 207124 467124
rect 217180 466244 217244 466308
rect 359964 465836 360028 465900
rect 55444 465700 55508 465764
rect 364932 465700 364996 465764
rect 376892 464340 376956 464404
rect 52316 463388 52380 463452
rect 203012 463388 203076 463452
rect 48084 463116 48148 463180
rect 204300 463116 204364 463180
rect 50476 462980 50540 463044
rect 359780 462980 359844 463044
rect 198964 462844 199028 462908
rect 377628 462844 377692 462908
rect 510844 462164 510908 462228
rect 179644 461680 179708 461684
rect 179644 461624 179658 461680
rect 179658 461624 179708 461680
rect 179644 461620 179708 461624
rect 58572 461484 58636 461548
rect 200804 461484 200868 461548
rect 178356 461408 178420 461412
rect 178356 461352 178370 461408
rect 178370 461352 178420 461408
rect 178356 461348 178420 461352
rect 190868 461000 190932 461004
rect 190868 460944 190918 461000
rect 190918 460944 190932 461000
rect 190868 460940 190932 460944
rect 338252 461000 338316 461004
rect 338252 460944 338302 461000
rect 338302 460944 338316 461000
rect 338252 460940 338316 460944
rect 339724 461000 339788 461004
rect 339724 460944 339774 461000
rect 339774 460944 339788 461000
rect 339724 460940 339788 460944
rect 350948 461000 351012 461004
rect 350948 460944 350998 461000
rect 350998 460944 351012 461000
rect 350948 460940 351012 460944
rect 498516 460940 498580 461004
rect 499804 461000 499868 461004
rect 499804 460944 499854 461000
rect 499854 460944 499868 461000
rect 499804 460940 499868 460944
rect 55076 460804 55140 460868
rect 206324 460804 206388 460868
rect 54892 460668 54956 460732
rect 210372 460668 210436 460732
rect 53420 460532 53484 460596
rect 213132 460532 213196 460596
rect 46612 460396 46676 460460
rect 205220 460396 205284 460460
rect 51948 460260 52012 460324
rect 206140 460260 206204 460324
rect 44956 460124 45020 460188
rect 215524 460124 215588 460188
rect 59124 459988 59188 460052
rect 198780 459988 198844 460052
rect 218652 459716 218716 459780
rect 48636 459640 48700 459644
rect 48636 459584 48686 459640
rect 48686 459584 48700 459640
rect 48636 459580 48700 459584
rect 51580 459640 51644 459644
rect 51580 459584 51630 459640
rect 51630 459584 51644 459640
rect 51580 459580 51644 459584
rect 52132 459580 52196 459644
rect 53604 459580 53668 459644
rect 55628 459580 55692 459644
rect 58940 459036 59004 459100
rect 207980 459036 208044 459100
rect 58756 458900 58820 458964
rect 57836 458764 57900 458828
rect 206692 408580 206756 408644
rect 360148 408580 360212 408644
rect 199148 392668 199212 392732
rect 199148 391988 199212 392052
rect 199516 391988 199580 392052
rect 51580 383556 51644 383620
rect 57468 383556 57532 383620
rect 207060 382332 207124 382396
rect 53236 375260 53300 375324
rect 198228 375260 198292 375324
rect 200988 375260 201052 375324
rect 204300 375260 204364 375324
rect 405964 375048 406028 375052
rect 405964 374992 405978 375048
rect 405978 374992 406028 375048
rect 405964 374988 406028 374992
rect 407804 375048 407868 375052
rect 407804 374992 407818 375048
rect 407818 374992 407868 375048
rect 407804 374988 407868 374992
rect 425100 375048 425164 375052
rect 425100 374992 425114 375048
rect 425114 374992 425164 375048
rect 425100 374988 425164 374992
rect 440372 375048 440436 375052
rect 440372 374992 440386 375048
rect 440386 374992 440436 375048
rect 440372 374988 440436 374992
rect 443132 375048 443196 375052
rect 443132 374992 443146 375048
rect 443146 374992 443196 375048
rect 443132 374988 443196 374992
rect 452884 375048 452948 375052
rect 452884 374992 452898 375048
rect 452898 374992 452948 375048
rect 452884 374988 452948 374992
rect 163366 374640 163430 374644
rect 163366 374584 163410 374640
rect 163410 374584 163430 374640
rect 163366 374580 163430 374584
rect 165950 374640 166014 374644
rect 165950 374584 165986 374640
rect 165986 374584 166014 374640
rect 165950 374580 166014 374584
rect 206508 374580 206572 374644
rect 208348 374580 208412 374644
rect 209820 374580 209884 374644
rect 410742 374640 410806 374644
rect 410742 374584 410762 374640
rect 410762 374584 410806 374640
rect 410742 374580 410806 374584
rect 93598 374504 93662 374508
rect 93598 374448 93638 374504
rect 93638 374448 93662 374504
rect 93598 374444 93662 374448
rect 103526 374504 103590 374508
rect 103526 374448 103574 374504
rect 103574 374448 103590 374504
rect 103526 374444 103590 374448
rect 116038 374504 116102 374508
rect 116038 374448 116086 374504
rect 116086 374448 116102 374504
rect 116038 374444 116102 374448
rect 143510 374504 143574 374508
rect 143510 374448 143538 374504
rect 143538 374448 143574 374504
rect 143510 374444 143574 374448
rect 146156 374504 146220 374508
rect 146156 374448 146206 374504
rect 146206 374448 146220 374504
rect 146156 374444 146220 374448
rect 153438 374504 153502 374508
rect 153438 374448 153474 374504
rect 153474 374448 153502 374504
rect 153438 374444 153502 374448
rect 156460 374504 156524 374508
rect 156460 374448 156510 374504
rect 156510 374448 156524 374504
rect 156460 374444 156524 374448
rect 158484 374504 158548 374508
rect 158484 374448 158534 374504
rect 158534 374448 158548 374504
rect 158484 374444 158548 374448
rect 160918 374504 160982 374508
rect 160918 374448 160926 374504
rect 160926 374448 160982 374504
rect 160918 374444 160982 374448
rect 236054 374444 236118 374508
rect 244228 374504 244292 374508
rect 244228 374448 244278 374504
rect 244278 374448 244292 374504
rect 244228 374444 244292 374448
rect 250062 374504 250126 374508
rect 250062 374448 250074 374504
rect 250074 374448 250126 374504
rect 250062 374444 250126 374448
rect 250742 374504 250806 374508
rect 250742 374448 250774 374504
rect 250774 374448 250806 374504
rect 250742 374444 250806 374448
rect 251286 374504 251350 374508
rect 251286 374448 251326 374504
rect 251326 374448 251350 374504
rect 251286 374444 251350 374448
rect 256046 374504 256110 374508
rect 256046 374448 256054 374504
rect 256054 374448 256110 374504
rect 256046 374444 256110 374448
rect 271142 374444 271206 374508
rect 320918 374504 320982 374508
rect 320918 374448 320970 374504
rect 320970 374448 320982 374504
rect 320918 374444 320982 374448
rect 433590 374504 433654 374508
rect 433590 374448 433614 374504
rect 433614 374448 433654 374504
rect 433590 374444 433654 374448
rect 436038 374504 436102 374508
rect 436038 374448 436062 374504
rect 436062 374448 436102 374504
rect 436038 374444 436102 374448
rect 438486 374504 438550 374508
rect 438486 374448 438490 374504
rect 438490 374448 438546 374504
rect 438546 374448 438550 374504
rect 438486 374444 438550 374448
rect 263732 374308 263796 374372
rect 148916 374232 148980 374236
rect 148916 374176 148966 374232
rect 148966 374176 148980 374232
rect 148916 374172 148980 374176
rect 275140 374036 275204 374100
rect 416084 374096 416148 374100
rect 416084 374040 416098 374096
rect 416098 374040 416148 374096
rect 416084 374036 416148 374040
rect 377444 373900 377508 373964
rect 485820 373900 485884 373964
rect 83780 373764 83844 373828
rect 268516 373764 268580 373828
rect 377628 373764 377692 373828
rect 460980 373764 461044 373828
rect 100892 373688 100956 373692
rect 100892 373632 100906 373688
rect 100906 373632 100956 373688
rect 100892 373628 100956 373632
rect 107884 373688 107948 373692
rect 107884 373632 107898 373688
rect 107898 373632 107948 373688
rect 107884 373628 107948 373632
rect 113588 373688 113652 373692
rect 113588 373632 113602 373688
rect 113602 373632 113652 373688
rect 113588 373628 113652 373632
rect 118372 373688 118436 373692
rect 118372 373632 118386 373688
rect 118386 373632 118436 373688
rect 118372 373628 118436 373632
rect 121316 373688 121380 373692
rect 121316 373632 121366 373688
rect 121366 373632 121380 373688
rect 121316 373628 121380 373632
rect 125732 373688 125796 373692
rect 125732 373632 125782 373688
rect 125782 373632 125796 373688
rect 125732 373628 125796 373632
rect 128860 373688 128924 373692
rect 128860 373632 128910 373688
rect 128910 373632 128924 373688
rect 128860 373628 128924 373632
rect 131068 373688 131132 373692
rect 131068 373632 131082 373688
rect 131082 373632 131132 373688
rect 131068 373628 131132 373632
rect 133644 373688 133708 373692
rect 133644 373632 133694 373688
rect 133694 373632 133708 373688
rect 133644 373628 133708 373632
rect 136404 373688 136468 373692
rect 136404 373632 136454 373688
rect 136454 373632 136468 373688
rect 136404 373628 136468 373632
rect 139164 373688 139228 373692
rect 139164 373632 139214 373688
rect 139214 373632 139228 373688
rect 139164 373628 139228 373632
rect 141556 373688 141620 373692
rect 141556 373632 141606 373688
rect 141606 373632 141620 373688
rect 141556 373628 141620 373632
rect 151676 373688 151740 373692
rect 151676 373632 151726 373688
rect 151726 373632 151740 373688
rect 151676 373628 151740 373632
rect 359596 373628 359660 373692
rect 418292 373688 418356 373692
rect 418292 373632 418306 373688
rect 418306 373632 418356 373688
rect 105492 373552 105556 373556
rect 105492 373496 105506 373552
rect 105506 373496 105556 373552
rect 105492 373492 105556 373496
rect 110460 373552 110524 373556
rect 110460 373496 110474 373552
rect 110474 373496 110524 373552
rect 110460 373492 110524 373496
rect 119844 373492 119908 373556
rect 255452 373552 255516 373556
rect 255452 373496 255466 373552
rect 255466 373496 255516 373552
rect 88380 373416 88444 373420
rect 88380 373360 88394 373416
rect 88394 373360 88444 373416
rect 88380 373356 88444 373360
rect 96108 373416 96172 373420
rect 96108 373360 96122 373416
rect 96122 373360 96172 373416
rect 96108 373356 96172 373360
rect 98316 373416 98380 373420
rect 98316 373360 98330 373416
rect 98330 373360 98380 373416
rect 98316 373356 98380 373360
rect 122972 373416 123036 373420
rect 122972 373360 122986 373416
rect 122986 373360 123036 373416
rect 122972 373356 123036 373360
rect 255452 373492 255516 373496
rect 256740 373552 256804 373556
rect 256740 373496 256754 373552
rect 256754 373496 256804 373552
rect 256740 373492 256804 373496
rect 418292 373628 418356 373632
rect 423076 373688 423140 373692
rect 423076 373632 423090 373688
rect 423090 373632 423140 373688
rect 423076 373628 423140 373632
rect 426940 373688 427004 373692
rect 426940 373632 426954 373688
rect 426954 373632 427004 373688
rect 426940 373628 427004 373632
rect 445892 373688 445956 373692
rect 445892 373632 445906 373688
rect 445906 373632 445956 373688
rect 445892 373628 445956 373632
rect 427860 373492 427924 373556
rect 450308 373552 450372 373556
rect 450308 373496 450322 373552
rect 450322 373496 450372 373552
rect 450308 373492 450372 373496
rect 455460 373552 455524 373556
rect 455460 373496 455474 373552
rect 455474 373496 455524 373552
rect 455460 373492 455524 373496
rect 236500 373416 236564 373420
rect 236500 373360 236514 373416
rect 236514 373360 236564 373416
rect 236500 373356 236564 373360
rect 242940 373416 243004 373420
rect 242940 373360 242954 373416
rect 242954 373360 243004 373416
rect 242940 373356 243004 373360
rect 260052 373416 260116 373420
rect 260052 373360 260066 373416
rect 260066 373360 260116 373416
rect 260052 373356 260116 373360
rect 269252 373416 269316 373420
rect 269252 373360 269266 373416
rect 269266 373360 269316 373416
rect 269252 373356 269316 373360
rect 447732 373416 447796 373420
rect 447732 373360 447746 373416
rect 447746 373360 447796 373416
rect 447732 373356 447796 373360
rect 462820 373416 462884 373420
rect 462820 373360 462834 373416
rect 462834 373360 462884 373416
rect 462820 373356 462884 373360
rect 278820 373220 278884 373284
rect 359964 373220 360028 373284
rect 408540 373220 408604 373284
rect 90220 373144 90284 373148
rect 90220 373088 90234 373144
rect 90234 373088 90284 373144
rect 90220 373084 90284 373088
rect 92428 373144 92492 373148
rect 92428 373088 92442 373144
rect 92442 373088 92492 373144
rect 92428 373084 92492 373088
rect 95188 373084 95252 373148
rect 247172 373144 247236 373148
rect 247172 373088 247186 373144
rect 247186 373088 247236 373144
rect 247172 373084 247236 373088
rect 253980 373144 254044 373148
rect 253980 373088 253994 373144
rect 253994 373088 254044 373144
rect 253980 373084 254044 373088
rect 257844 373084 257908 373148
rect 261340 373144 261404 373148
rect 261340 373088 261354 373144
rect 261354 373088 261404 373144
rect 261340 373084 261404 373088
rect 265020 373144 265084 373148
rect 265020 373088 265034 373144
rect 265034 373088 265084 373144
rect 265020 373084 265084 373088
rect 300900 373144 300964 373148
rect 300900 373088 300914 373144
rect 300914 373088 300964 373144
rect 300900 373084 300964 373088
rect 57284 372676 57348 372740
rect 216996 372676 217060 372740
rect 252876 372676 252940 372740
rect 362908 372676 362972 372740
rect 376892 372676 376956 372740
rect 77156 372600 77220 372604
rect 77156 372544 77206 372600
rect 77206 372544 77220 372600
rect 77156 372540 77220 372544
rect 81940 372600 82004 372604
rect 81940 372544 81990 372600
rect 81990 372544 82004 372600
rect 81940 372540 82004 372544
rect 84700 372600 84764 372604
rect 84700 372544 84750 372600
rect 84750 372544 84764 372600
rect 84700 372540 84764 372544
rect 86724 372600 86788 372604
rect 86724 372544 86774 372600
rect 86774 372544 86788 372600
rect 86724 372540 86788 372544
rect 88012 372600 88076 372604
rect 88012 372544 88062 372600
rect 88062 372544 88076 372600
rect 88012 372540 88076 372544
rect 89300 372600 89364 372604
rect 89300 372544 89350 372600
rect 89350 372544 89364 372600
rect 89300 372540 89364 372544
rect 90036 372540 90100 372604
rect 91508 372540 91572 372604
rect 93348 372540 93412 372604
rect 101996 372600 102060 372604
rect 101996 372544 102046 372600
rect 102046 372544 102060 372600
rect 101996 372540 102060 372544
rect 112852 372600 112916 372604
rect 112852 372544 112902 372600
rect 112902 372544 112916 372600
rect 112852 372540 112916 372544
rect 114508 372600 114572 372604
rect 114508 372544 114522 372600
rect 114522 372544 114572 372600
rect 114508 372540 114572 372544
rect 238156 372600 238220 372604
rect 238156 372544 238170 372600
rect 238170 372544 238220 372600
rect 238156 372540 238220 372544
rect 239260 372600 239324 372604
rect 239260 372544 239310 372600
rect 239310 372544 239324 372600
rect 239260 372540 239324 372544
rect 240364 372600 240428 372604
rect 240364 372544 240414 372600
rect 240414 372544 240428 372600
rect 240364 372540 240428 372544
rect 241652 372600 241716 372604
rect 241652 372544 241702 372600
rect 241702 372544 241716 372600
rect 241652 372540 241716 372544
rect 244780 372540 244844 372604
rect 248460 372600 248524 372604
rect 248460 372544 248474 372600
rect 248474 372544 248524 372600
rect 248460 372540 248524 372544
rect 251772 372540 251836 372604
rect 259500 372600 259564 372604
rect 259500 372544 259514 372600
rect 259514 372544 259564 372600
rect 259500 372540 259564 372544
rect 262260 372600 262324 372604
rect 262260 372544 262274 372600
rect 262274 372544 262324 372600
rect 262260 372540 262324 372544
rect 266308 372600 266372 372604
rect 266308 372544 266358 372600
rect 266358 372544 266372 372600
rect 266308 372540 266372 372544
rect 272564 372540 272628 372604
rect 310652 372540 310716 372604
rect 315068 372540 315132 372604
rect 322980 372600 323044 372604
rect 322980 372544 322994 372600
rect 322994 372544 323044 372600
rect 322980 372540 323044 372544
rect 400260 372600 400324 372604
rect 400260 372544 400274 372600
rect 400274 372544 400324 372600
rect 400260 372540 400324 372544
rect 403572 372540 403636 372604
rect 78444 372464 78508 372468
rect 78444 372408 78494 372464
rect 78494 372408 78508 372464
rect 78444 372404 78508 372408
rect 79916 372464 79980 372468
rect 79916 372408 79966 372464
rect 79966 372408 79980 372464
rect 79916 372404 79980 372408
rect 80468 372404 80532 372468
rect 84516 372404 84580 372468
rect 118188 372404 118252 372468
rect 277532 372404 277596 372468
rect 313412 372404 313476 372468
rect 376892 372404 376956 372468
rect 433564 372404 433628 372468
rect 104572 372192 104636 372196
rect 104572 372136 104622 372192
rect 104622 372136 104636 372192
rect 104572 372132 104636 372136
rect 109540 372132 109604 372196
rect 276980 372328 277044 372332
rect 276980 372272 276994 372328
rect 276994 372272 277044 372328
rect 276980 372268 277044 372272
rect 305316 372268 305380 372332
rect 438900 372268 438964 372332
rect 470732 372268 470796 372332
rect 396212 372132 396276 372196
rect 503116 372192 503180 372196
rect 503116 372136 503166 372192
rect 503166 372136 503180 372192
rect 503116 372132 503180 372136
rect 503484 372192 503548 372196
rect 503484 372136 503534 372192
rect 503534 372136 503548 372192
rect 503484 372132 503548 372136
rect 113220 371996 113284 372060
rect 273300 371996 273364 372060
rect 397500 372056 397564 372060
rect 397500 372000 397514 372056
rect 397514 372000 397564 372056
rect 397500 371996 397564 372000
rect 404860 371996 404924 372060
rect 407252 371996 407316 372060
rect 422340 372056 422404 372060
rect 422340 372000 422354 372056
rect 422354 372000 422404 372056
rect 422340 371996 422404 372000
rect 76604 371860 76668 371924
rect 108988 371860 109052 371924
rect 115796 371724 115860 371788
rect 377812 371860 377876 371924
rect 438348 371860 438412 371924
rect 483244 371860 483308 371924
rect 245884 371724 245948 371788
rect 273668 371724 273732 371788
rect 317828 371724 317892 371788
rect 402284 371724 402348 371788
rect 410012 371724 410076 371788
rect 95188 371648 95252 371652
rect 95188 371592 95238 371648
rect 95238 371592 95252 371648
rect 95188 371588 95252 371592
rect 98132 371588 98196 371652
rect 99972 371588 100036 371652
rect 105308 371588 105372 371652
rect 182956 371588 183020 371652
rect 183324 371588 183388 371652
rect 217548 371588 217612 371652
rect 398972 371588 399036 371652
rect 411300 371648 411364 371652
rect 411300 371592 411314 371648
rect 411314 371592 411364 371648
rect 411300 371588 411364 371592
rect 465396 371588 465460 371652
rect 97580 371452 97644 371516
rect 100708 371452 100772 371516
rect 111748 371452 111812 371516
rect 57100 371316 57164 371380
rect 102732 371316 102796 371380
rect 107516 371376 107580 371380
rect 107516 371320 107566 371376
rect 107566 371320 107580 371376
rect 107516 371316 107580 371320
rect 117084 371316 117148 371380
rect 278268 371452 278332 371516
rect 411852 371452 411916 371516
rect 418844 371452 418908 371516
rect 421236 371452 421300 371516
rect 423996 371452 424060 371516
rect 426388 371512 426452 371516
rect 426388 371456 426438 371512
rect 426438 371456 426452 371512
rect 426388 371452 426452 371456
rect 431172 371452 431236 371516
rect 247908 371316 247972 371380
rect 253612 371316 253676 371380
rect 258396 371316 258460 371380
rect 260972 371316 261036 371380
rect 263548 371376 263612 371380
rect 263548 371320 263598 371376
rect 263598 371320 263612 371376
rect 263548 371316 263612 371320
rect 265756 371316 265820 371380
rect 267044 371316 267108 371380
rect 267780 371376 267844 371380
rect 267780 371320 267794 371376
rect 267794 371320 267844 371376
rect 267780 371316 267844 371320
rect 270908 371316 270972 371380
rect 273852 371316 273916 371380
rect 276244 371316 276308 371380
rect 280292 371316 280356 371380
rect 283788 371316 283852 371380
rect 285812 371316 285876 371380
rect 287652 371316 287716 371380
rect 290596 371316 290660 371380
rect 292804 371316 292868 371380
rect 295380 371376 295444 371380
rect 295380 371320 295394 371376
rect 295394 371320 295444 371376
rect 295380 371316 295444 371320
rect 298140 371376 298204 371380
rect 298140 371320 298154 371376
rect 298154 371320 298204 371376
rect 298140 371316 298204 371320
rect 302924 371316 302988 371380
rect 308628 371316 308692 371380
rect 326660 371316 326724 371380
rect 343036 371316 343100 371380
rect 343404 371376 343468 371380
rect 343404 371320 343418 371376
rect 343418 371320 343468 371376
rect 343404 371316 343468 371320
rect 396580 371316 396644 371380
rect 403020 371376 403084 371380
rect 403020 371320 403034 371376
rect 403034 371320 403084 371376
rect 403020 371316 403084 371320
rect 412772 371316 412836 371380
rect 413692 371316 413756 371380
rect 414060 371376 414124 371380
rect 414060 371320 414074 371376
rect 414074 371320 414124 371376
rect 414060 371316 414124 371320
rect 415532 371316 415596 371380
rect 416820 371376 416884 371380
rect 416820 371320 416834 371376
rect 416834 371320 416884 371376
rect 416820 371316 416884 371320
rect 418108 371376 418172 371380
rect 418108 371320 418158 371376
rect 418158 371320 418172 371376
rect 418108 371316 418172 371320
rect 420316 371316 420380 371380
rect 421052 371316 421116 371380
rect 425652 371316 425716 371380
rect 428596 371316 428660 371380
rect 429332 371316 429396 371380
rect 430620 371376 430684 371380
rect 430620 371320 430634 371376
rect 430634 371320 430684 371376
rect 430620 371316 430684 371320
rect 432092 371316 432156 371380
rect 433380 371376 433444 371380
rect 433380 371320 433394 371376
rect 433394 371320 433444 371376
rect 433380 371316 433444 371320
rect 434852 371316 434916 371380
rect 436324 371316 436388 371380
rect 458220 371376 458284 371380
rect 458220 371320 458234 371376
rect 458234 371320 458284 371376
rect 458220 371316 458284 371320
rect 473308 371376 473372 371380
rect 473308 371320 473358 371376
rect 473358 371320 473372 371376
rect 473308 371316 473372 371320
rect 475332 371316 475396 371380
rect 478092 371316 478156 371380
rect 480300 371376 480364 371380
rect 480300 371320 480314 371376
rect 480314 371320 480364 371376
rect 480300 371316 480364 371320
rect 359780 371180 359844 371244
rect 467972 371180 468036 371244
rect 106412 371044 106476 371108
rect 216996 371044 217060 371108
rect 212764 369140 212828 369204
rect 215524 369140 215588 369204
rect 376892 368520 376956 368524
rect 376892 368464 376942 368520
rect 376942 368464 376956 368520
rect 376892 368460 376956 368464
rect 217364 368324 217428 368388
rect 199516 357988 199580 358052
rect 178540 355268 178604 355332
rect 190868 355268 190932 355332
rect 338436 355056 338500 355060
rect 338436 355000 338486 355056
rect 338486 355000 338500 355056
rect 338436 354996 338500 355000
rect 350948 354996 351012 355060
rect 498516 354996 498580 355060
rect 499804 354860 499868 354924
rect 179644 354784 179708 354788
rect 179644 354728 179694 354784
rect 179694 354728 179708 354784
rect 179644 354724 179708 354728
rect 339724 354784 339788 354788
rect 339724 354728 339774 354784
rect 339774 354728 339788 354784
rect 339724 354724 339788 354728
rect 510844 354784 510908 354788
rect 510844 354728 510894 354784
rect 510894 354728 510908 354784
rect 510844 354724 510908 354728
rect 217364 353364 217428 353428
rect 54340 304948 54404 305012
rect 57100 276116 57164 276180
rect 57284 275980 57348 276044
rect 216628 270540 216692 270604
rect 217364 270540 217428 270604
rect 211844 270404 211908 270468
rect 218836 270404 218900 270468
rect 378180 270404 378244 270468
rect 377996 270268 378060 270332
rect 107606 269920 107670 269924
rect 107606 269864 107622 269920
rect 107622 269864 107670 269920
rect 107606 269860 107670 269864
rect 111006 269920 111070 269924
rect 111006 269864 111026 269920
rect 111026 269864 111070 269920
rect 111006 269860 111070 269864
rect 250742 269920 250806 269924
rect 250742 269864 250774 269920
rect 250774 269864 250806 269920
rect 250742 269860 250806 269864
rect 266382 269860 266446 269924
rect 108286 269784 108350 269788
rect 108286 269728 108302 269784
rect 108302 269728 108350 269784
rect 108286 269724 108350 269728
rect 133446 269784 133510 269788
rect 133446 269728 133474 269784
rect 133474 269728 133510 269784
rect 133446 269724 133510 269728
rect 135894 269784 135958 269788
rect 135894 269728 135902 269784
rect 135902 269728 135958 269784
rect 135894 269724 135958 269728
rect 138478 269784 138542 269788
rect 138478 269728 138534 269784
rect 138534 269728 138542 269784
rect 138478 269724 138542 269728
rect 216628 269724 216692 269788
rect 274406 269724 274470 269788
rect 275766 269784 275830 269788
rect 275766 269728 275798 269784
rect 275798 269728 275830 269784
rect 275766 269724 275830 269728
rect 280934 269784 280998 269788
rect 280934 269728 280950 269784
rect 280950 269728 280998 269784
rect 280934 269724 280998 269728
rect 315886 269784 315950 269788
rect 315886 269728 315910 269784
rect 315910 269728 315950 269784
rect 315886 269724 315950 269728
rect 418494 269724 418558 269788
rect 425294 269784 425358 269788
rect 425294 269728 425298 269784
rect 425298 269728 425358 269784
rect 425294 269724 425358 269728
rect 83126 269648 83190 269652
rect 83126 269592 83150 269648
rect 83150 269592 83190 269648
rect 83126 269588 83190 269592
rect 93598 269648 93662 269652
rect 93598 269592 93638 269648
rect 93638 269592 93662 269648
rect 93598 269588 93662 269592
rect 94550 269648 94614 269652
rect 94550 269592 94558 269648
rect 94558 269592 94614 269648
rect 94550 269588 94614 269592
rect 108694 269648 108758 269652
rect 108694 269592 108726 269648
rect 108726 269592 108758 269648
rect 108694 269588 108758 269592
rect 140926 269588 140990 269652
rect 143510 269648 143574 269652
rect 143510 269592 143538 269648
rect 143538 269592 143574 269648
rect 143510 269588 143574 269592
rect 145958 269648 146022 269652
rect 145958 269592 145986 269648
rect 145986 269592 146022 269648
rect 145958 269588 146022 269592
rect 279166 269648 279230 269652
rect 279166 269592 279202 269648
rect 279202 269592 279230 269648
rect 279166 269588 279230 269592
rect 283518 269648 283582 269652
rect 283518 269592 283526 269648
rect 283526 269592 283582 269648
rect 283518 269588 283582 269592
rect 285966 269648 286030 269652
rect 285966 269592 286010 269648
rect 286010 269592 286030 269648
rect 285966 269588 286030 269592
rect 288278 269648 288342 269652
rect 288278 269592 288310 269648
rect 288310 269592 288342 269648
rect 288278 269588 288342 269592
rect 293446 269648 293510 269652
rect 293446 269592 293462 269648
rect 293462 269592 293510 269648
rect 293446 269588 293510 269592
rect 308542 269648 308606 269652
rect 308542 269592 308550 269648
rect 308550 269592 308606 269648
rect 308542 269588 308606 269592
rect 318470 269648 318534 269652
rect 318470 269592 318486 269648
rect 318486 269592 318534 269648
rect 318470 269588 318534 269592
rect 423526 269648 423590 269652
rect 423526 269592 423550 269648
rect 423550 269592 423590 269648
rect 423526 269588 423590 269592
rect 426388 269648 426452 269652
rect 426388 269592 426438 269648
rect 426438 269592 426452 269648
rect 426388 269588 426452 269592
rect 433590 269648 433654 269652
rect 433590 269592 433614 269648
rect 433614 269592 433654 269648
rect 433590 269588 433654 269592
rect 453446 269648 453510 269652
rect 453446 269592 453450 269648
rect 453450 269592 453510 269648
rect 453446 269588 453510 269592
rect 468542 269588 468606 269652
rect 480918 269648 480982 269652
rect 480918 269592 480958 269648
rect 480958 269592 480982 269648
rect 480918 269588 480982 269592
rect 376892 269316 376956 269380
rect 377628 269316 377692 269380
rect 359412 269180 359476 269244
rect 470916 269180 470980 269244
rect 57284 269044 57348 269108
rect 76052 269104 76116 269108
rect 76052 269048 76066 269104
rect 76066 269048 76116 269104
rect 76052 269044 76116 269048
rect 77156 269104 77220 269108
rect 77156 269048 77170 269104
rect 77170 269048 77220 269104
rect 77156 269044 77220 269048
rect 90772 269104 90836 269108
rect 90772 269048 90786 269104
rect 90786 269048 90836 269104
rect 90772 269044 90836 269048
rect 95924 269104 95988 269108
rect 95924 269048 95938 269104
rect 95938 269048 95988 269104
rect 95924 269044 95988 269048
rect 96108 269104 96172 269108
rect 96108 269048 96122 269104
rect 96122 269048 96172 269104
rect 96108 269044 96172 269048
rect 98500 269104 98564 269108
rect 98500 269048 98514 269104
rect 98514 269048 98564 269104
rect 98500 269044 98564 269048
rect 99420 269104 99484 269108
rect 99420 269048 99434 269104
rect 99434 269048 99484 269104
rect 99420 269044 99484 269048
rect 212580 269044 212644 269108
rect 217180 269044 217244 269108
rect 115796 268908 115860 268972
rect 199332 268908 199396 268972
rect 278452 268908 278516 268972
rect 290964 268968 291028 268972
rect 290964 268912 290978 268968
rect 290978 268912 291028 268968
rect 290964 268908 291028 268912
rect 295932 268968 295996 268972
rect 298508 269104 298572 269108
rect 298508 269048 298522 269104
rect 298522 269048 298572 269104
rect 298508 269044 298572 269048
rect 300900 269104 300964 269108
rect 300900 269048 300914 269104
rect 300914 269048 300964 269104
rect 300900 269044 300964 269048
rect 486004 269044 486068 269108
rect 295932 268912 295946 268968
rect 295946 268912 295996 268968
rect 295932 268908 295996 268912
rect 305868 268908 305932 268972
rect 377260 268908 377324 268972
rect 426020 268908 426084 268972
rect 430988 268968 431052 268972
rect 430988 268912 431002 268968
rect 431002 268912 431052 268968
rect 430988 268908 431052 268912
rect 433380 268968 433444 268972
rect 433380 268912 433394 268968
rect 433394 268912 433444 268968
rect 433380 268908 433444 268912
rect 475884 268968 475948 268972
rect 475884 268912 475898 268968
rect 475898 268912 475948 268968
rect 475884 268908 475948 268912
rect 478460 268968 478524 268972
rect 478460 268912 478474 268968
rect 478474 268912 478524 268968
rect 478460 268908 478524 268912
rect 483428 268968 483492 268972
rect 483428 268912 483442 268968
rect 483442 268912 483492 268968
rect 483428 268908 483492 268912
rect 118004 268772 118068 268836
rect 243124 268832 243188 268836
rect 243124 268776 243138 268832
rect 243138 268776 243188 268832
rect 243124 268772 243188 268776
rect 257844 268772 257908 268836
rect 261708 268832 261772 268836
rect 261708 268776 261722 268832
rect 261722 268776 261772 268832
rect 261708 268772 261772 268776
rect 377628 268772 377692 268836
rect 119108 268636 119172 268700
rect 415900 268832 415964 268836
rect 415900 268776 415914 268832
rect 415914 268776 415964 268832
rect 415900 268772 415964 268776
rect 421052 268832 421116 268836
rect 421052 268776 421066 268832
rect 421066 268776 421116 268832
rect 421052 268772 421116 268776
rect 423996 268636 424060 268700
rect 109724 268500 109788 268564
rect 111196 268364 111260 268428
rect 85436 268152 85500 268156
rect 85436 268096 85450 268152
rect 85450 268096 85500 268152
rect 85436 268092 85500 268096
rect 92428 268152 92492 268156
rect 92428 268096 92442 268152
rect 92442 268096 92492 268152
rect 92428 268092 92492 268096
rect 103284 268092 103348 268156
rect 113588 268092 113652 268156
rect 128308 268152 128372 268156
rect 128308 268096 128358 268152
rect 128358 268096 128372 268152
rect 128308 268092 128372 268096
rect 153516 268152 153580 268156
rect 153516 268096 153566 268152
rect 153566 268096 153580 268152
rect 153516 268092 153580 268096
rect 113220 268016 113284 268020
rect 113220 267960 113270 268016
rect 113270 267960 113284 268016
rect 113220 267956 113284 267960
rect 265204 268152 265268 268156
rect 265204 268096 265218 268152
rect 265218 268096 265268 268152
rect 265204 268092 265268 268096
rect 272196 268152 272260 268156
rect 272196 268096 272210 268152
rect 272210 268096 272260 268152
rect 272196 268092 272260 268096
rect 398236 268152 398300 268156
rect 398236 268096 398250 268152
rect 398250 268096 398300 268152
rect 398236 268092 398300 268096
rect 401732 268152 401796 268156
rect 401732 268096 401746 268152
rect 401746 268096 401796 268152
rect 401732 268092 401796 268096
rect 416084 268152 416148 268156
rect 416084 268096 416098 268152
rect 416098 268096 416148 268152
rect 416084 268092 416148 268096
rect 434300 268152 434364 268156
rect 434300 268096 434314 268152
rect 434314 268096 434364 268152
rect 434300 268092 434364 268096
rect 455828 268152 455892 268156
rect 455828 268096 455842 268152
rect 455842 268096 455892 268152
rect 455828 268092 455892 268096
rect 83964 267684 84028 267748
rect 87460 267684 87524 267748
rect 102732 267744 102796 267748
rect 102732 267688 102746 267744
rect 102746 267688 102796 267744
rect 102732 267684 102796 267688
rect 105308 267744 105372 267748
rect 105308 267688 105322 267744
rect 105322 267688 105372 267744
rect 105308 267684 105372 267688
rect 106412 267744 106476 267748
rect 106412 267688 106426 267744
rect 106426 267688 106476 267744
rect 106412 267684 106476 267688
rect 117084 267744 117148 267748
rect 117084 267688 117134 267744
rect 117134 267688 117148 267744
rect 117084 267684 117148 267688
rect 123524 267684 123588 267748
rect 130884 267684 130948 267748
rect 155908 267744 155972 267748
rect 155908 267688 155958 267744
rect 155958 267688 155972 267744
rect 155908 267684 155972 267688
rect 158484 267744 158548 267748
rect 158484 267688 158534 267744
rect 158534 267688 158548 267744
rect 158484 267684 158548 267688
rect 163452 267744 163516 267748
rect 163452 267688 163502 267744
rect 163502 267688 163516 267744
rect 163452 267684 163516 267688
rect 255820 267744 255884 267748
rect 255820 267688 255834 267744
rect 255834 267688 255884 267744
rect 255820 267684 255884 267688
rect 260972 267684 261036 267748
rect 263732 267684 263796 267748
rect 265940 267684 266004 267748
rect 267596 267684 267660 267748
rect 268332 267684 268396 267748
rect 270908 267744 270972 267748
rect 270908 267688 270922 267744
rect 270922 267688 270972 267744
rect 270908 267684 270972 267688
rect 273484 267684 273548 267748
rect 276244 267684 276308 267748
rect 303476 267684 303540 267748
rect 403020 267744 403084 267748
rect 403020 267688 403034 267744
rect 403034 267688 403084 267744
rect 403020 267684 403084 267688
rect 414428 267744 414492 267748
rect 414428 267688 414442 267744
rect 414442 267688 414492 267744
rect 414428 267684 414492 267688
rect 432276 267684 432340 267748
rect 435772 267744 435836 267748
rect 435772 267688 435786 267744
rect 435786 267688 435836 267744
rect 435772 267684 435836 267688
rect 435956 267744 436020 267748
rect 435956 267688 435970 267744
rect 435970 267688 436020 267744
rect 435956 267684 436020 267688
rect 445892 267684 445956 267748
rect 448284 267684 448348 267748
rect 451044 267684 451108 267748
rect 458404 267684 458468 267748
rect 473308 267744 473372 267748
rect 473308 267688 473358 267744
rect 473358 267688 473372 267744
rect 473308 267684 473372 267688
rect 79548 267548 79612 267612
rect 125916 267548 125980 267612
rect 150940 267548 151004 267612
rect 198964 267548 199028 267612
rect 323348 267548 323412 267612
rect 465948 267548 466012 267612
rect 81940 267412 82004 267476
rect 118372 267412 118436 267476
rect 120764 267412 120828 267476
rect 160876 267472 160940 267476
rect 160876 267416 160926 267472
rect 160926 267416 160940 267472
rect 160876 267412 160940 267416
rect 166028 267412 166092 267476
rect 183508 267472 183572 267476
rect 183508 267416 183522 267472
rect 183522 267416 183572 267472
rect 183508 267412 183572 267416
rect 320956 267412 321020 267476
rect 343404 267472 343468 267476
rect 343404 267416 343454 267472
rect 343454 267416 343468 267472
rect 343404 267412 343468 267416
rect 460980 267412 461044 267476
rect 503484 267472 503548 267476
rect 503484 267416 503534 267472
rect 503534 267416 503548 267472
rect 503484 267412 503548 267416
rect 115980 267336 116044 267340
rect 115980 267280 115994 267336
rect 115994 267280 116044 267336
rect 115980 267276 116044 267280
rect 183140 267276 183204 267340
rect 313412 267276 313476 267340
rect 343220 267276 343284 267340
rect 379468 267276 379532 267340
rect 428228 267276 428292 267340
rect 438532 267276 438596 267340
rect 443500 267276 443564 267340
rect 503116 267276 503180 267340
rect 88380 267200 88444 267204
rect 88380 267144 88394 267200
rect 88394 267144 88444 267200
rect 88380 267140 88444 267144
rect 101076 267140 101140 267204
rect 105860 267140 105924 267204
rect 238156 267140 238220 267204
rect 258396 267140 258460 267204
rect 269804 267200 269868 267204
rect 269804 267144 269818 267200
rect 269818 267144 269868 267200
rect 269804 267140 269868 267144
rect 271276 267200 271340 267204
rect 271276 267144 271290 267200
rect 271290 267144 271340 267200
rect 271276 267140 271340 267144
rect 276980 267140 277044 267204
rect 278084 267200 278148 267204
rect 278084 267144 278134 267200
rect 278134 267144 278148 267200
rect 278084 267140 278148 267144
rect 397132 267140 397196 267204
rect 440924 267140 440988 267204
rect 103836 267004 103900 267068
rect 236500 267004 236564 267068
rect 256188 267004 256252 267068
rect 273300 267064 273364 267068
rect 273300 267008 273314 267064
rect 273314 267008 273364 267064
rect 273300 267004 273364 267008
rect 396212 267004 396276 267068
rect 408172 267004 408236 267068
rect 410748 267004 410812 267068
rect 413692 267004 413756 267068
rect 422892 267004 422956 267068
rect 78260 266868 78324 266932
rect 80468 266868 80532 266932
rect 237052 266868 237116 266932
rect 248276 266868 248340 266932
rect 253612 266868 253676 266932
rect 263916 266868 263980 266932
rect 268700 266868 268764 266932
rect 311020 266868 311084 266932
rect 462636 266868 462700 266932
rect 326660 266732 326724 266796
rect 91324 266596 91388 266660
rect 100708 266520 100772 266524
rect 100708 266464 100758 266520
rect 100758 266464 100772 266520
rect 100708 266460 100772 266464
rect 244228 266460 244292 266524
rect 252324 266460 252388 266524
rect 260604 266460 260668 266524
rect 412404 266460 412468 266524
rect 419212 266460 419276 266524
rect 86540 266324 86604 266388
rect 88748 266324 88812 266388
rect 90036 266324 90100 266388
rect 93348 266324 93412 266388
rect 97028 266324 97092 266388
rect 98132 266324 98196 266388
rect 101812 266324 101876 266388
rect 112116 266324 112180 266388
rect 114508 266324 114572 266388
rect 148548 266324 148612 266388
rect 245332 266324 245396 266388
rect 246436 266324 246500 266388
rect 247724 266324 247788 266388
rect 248644 266324 248708 266388
rect 250116 266324 250180 266388
rect 251220 266384 251284 266388
rect 251220 266328 251234 266384
rect 251234 266328 251284 266384
rect 251220 266324 251284 266328
rect 253428 266324 253492 266388
rect 254532 266324 254596 266388
rect 256924 266324 256988 266388
rect 259500 266384 259564 266388
rect 259500 266328 259514 266384
rect 259514 266328 259564 266384
rect 259500 266324 259564 266328
rect 262812 266324 262876 266388
rect 279004 266324 279068 266388
rect 399524 266324 399588 266388
rect 400444 266324 400508 266388
rect 404124 266324 404188 266388
rect 405044 266324 405108 266388
rect 406516 266324 406580 266388
rect 407620 266324 407684 266388
rect 408724 266324 408788 266388
rect 410012 266324 410076 266388
rect 411300 266384 411364 266388
rect 411300 266328 411314 266384
rect 411314 266328 411364 266384
rect 411300 266324 411364 266328
rect 413324 266324 413388 266388
rect 417004 266324 417068 266388
rect 418108 266384 418172 266388
rect 418108 266328 418158 266384
rect 418158 266328 418172 266384
rect 418108 266324 418172 266328
rect 420684 266324 420748 266388
rect 421788 266324 421852 266388
rect 428780 266324 428844 266388
rect 429884 266324 429948 266388
rect 431172 266324 431236 266388
rect 436876 266324 436940 266388
rect 438348 266324 438412 266388
rect 439084 266324 439148 266388
rect 196756 266188 196820 266252
rect 217548 265916 217612 265980
rect 239260 266188 239324 266252
rect 240548 265644 240612 265708
rect 241652 265508 241716 265572
rect 427676 265508 427740 265572
rect 47900 264828 47964 264892
rect 377812 263468 377876 263532
rect 53052 253948 53116 254012
rect 215340 251092 215404 251156
rect 178540 249868 178604 249932
rect 179644 249868 179708 249932
rect 190868 249928 190932 249932
rect 190868 249872 190918 249928
rect 190918 249872 190932 249928
rect 190868 249868 190932 249872
rect 338436 249928 338500 249932
rect 338436 249872 338486 249928
rect 338486 249872 338500 249928
rect 338436 249868 338500 249872
rect 339724 249868 339788 249932
rect 350948 249928 351012 249932
rect 350948 249872 350998 249928
rect 350998 249872 351012 249928
rect 350948 249868 351012 249872
rect 498516 249868 498580 249932
rect 499804 249868 499868 249932
rect 510844 249928 510908 249932
rect 510844 249872 510894 249928
rect 510894 249872 510908 249928
rect 510844 249868 510908 249872
rect 58572 175204 58636 175268
rect 57468 173028 57532 173092
rect 96108 164792 96172 164796
rect 96108 164736 96122 164792
rect 96122 164736 96172 164792
rect 96108 164732 96172 164736
rect 140926 164732 140990 164796
rect 258494 164792 258558 164796
rect 258494 164736 258502 164792
rect 258502 164736 258558 164792
rect 258494 164732 258558 164736
rect 295894 164732 295958 164796
rect 425974 164792 426038 164796
rect 425974 164736 425978 164792
rect 425978 164736 426034 164792
rect 426034 164736 426038 164792
rect 425974 164732 426038 164736
rect 434406 164732 434470 164796
rect 450998 164792 451062 164796
rect 450998 164736 451002 164792
rect 451002 164736 451058 164792
rect 451058 164736 451062 164792
rect 450998 164732 451062 164736
rect 103526 164656 103590 164660
rect 103526 164600 103574 164656
rect 103574 164600 103590 164656
rect 103526 164596 103590 164600
rect 105974 164596 106038 164660
rect 116990 164656 117054 164660
rect 116990 164600 117042 164656
rect 117042 164600 117054 164656
rect 116990 164596 117054 164600
rect 153438 164596 153502 164660
rect 163366 164656 163430 164660
rect 163366 164600 163374 164656
rect 163374 164600 163430 164656
rect 163366 164596 163430 164600
rect 261078 164596 261142 164660
rect 275766 164596 275830 164660
rect 288278 164596 288342 164660
rect 305958 164656 306022 164660
rect 305958 164600 305974 164656
rect 305974 164600 306022 164656
rect 305958 164596 306022 164600
rect 318470 164656 318534 164660
rect 318470 164600 318486 164656
rect 318486 164600 318534 164656
rect 318470 164596 318534 164600
rect 423526 164656 423590 164660
rect 423526 164600 423550 164656
rect 423550 164600 423590 164656
rect 423526 164596 423590 164600
rect 436990 164596 437054 164660
rect 438078 164656 438142 164660
rect 438078 164600 438086 164656
rect 438086 164600 438142 164656
rect 438078 164596 438142 164600
rect 480918 164656 480982 164660
rect 480918 164600 480958 164656
rect 480958 164600 480982 164656
rect 480918 164596 480982 164600
rect 55444 164324 55508 164388
rect 138428 164324 138492 164388
rect 213132 164324 213196 164388
rect 98500 164248 98564 164252
rect 98500 164192 98514 164248
rect 98514 164192 98564 164248
rect 98500 164188 98564 164192
rect 101076 164248 101140 164252
rect 101076 164192 101090 164248
rect 101090 164192 101140 164248
rect 101076 164188 101140 164192
rect 108252 164248 108316 164252
rect 108252 164192 108266 164248
rect 108266 164192 108316 164248
rect 108252 164188 108316 164192
rect 145972 164248 146036 164252
rect 145972 164192 145986 164248
rect 145986 164192 146036 164248
rect 145972 164188 146036 164192
rect 148548 164248 148612 164252
rect 148548 164192 148562 164248
rect 148562 164192 148612 164248
rect 148548 164188 148612 164192
rect 150940 164248 151004 164252
rect 150940 164192 150954 164248
rect 150954 164192 151004 164248
rect 150940 164188 151004 164192
rect 210372 164188 210436 164252
rect 298508 164248 298572 164252
rect 298508 164192 298522 164248
rect 298522 164192 298572 164248
rect 298508 164188 298572 164192
rect 300900 164248 300964 164252
rect 300900 164192 300914 164248
rect 300914 164192 300964 164248
rect 300900 164188 300964 164192
rect 377812 164188 377876 164252
rect 416084 164248 416148 164252
rect 416084 164192 416098 164248
rect 416098 164192 416148 164248
rect 416084 164188 416148 164192
rect 421052 164248 421116 164252
rect 421052 164192 421066 164248
rect 421066 164192 421116 164248
rect 421052 164188 421116 164192
rect 428228 164248 428292 164252
rect 428228 164192 428242 164248
rect 428242 164192 428292 164248
rect 428228 164188 428292 164192
rect 430988 164248 431052 164252
rect 430988 164192 431002 164248
rect 431002 164192 431052 164248
rect 430988 164188 431052 164192
rect 473492 164248 473556 164252
rect 473492 164192 473506 164248
rect 473506 164192 473556 164248
rect 473492 164188 473556 164192
rect 475884 164248 475948 164252
rect 475884 164192 475898 164248
rect 475898 164192 475948 164248
rect 475884 164188 475948 164192
rect 478460 164248 478524 164252
rect 478460 164192 478474 164248
rect 478474 164192 478524 164248
rect 478460 164188 478524 164192
rect 57652 164052 57716 164116
rect 143580 164052 143644 164116
rect 202460 164052 202524 164116
rect 323348 164052 323412 164116
rect 486004 164052 486068 164116
rect 203012 163916 203076 163980
rect 311020 163916 311084 163980
rect 483428 163916 483492 163980
rect 206324 163780 206388 163844
rect 313412 163780 313476 163844
rect 470364 163780 470428 163844
rect 207980 163644 208044 163708
rect 315804 163644 315868 163708
rect 198044 163508 198108 163572
rect 290964 163508 291028 163572
rect 196572 163372 196636 163436
rect 270908 163372 270972 163436
rect 85436 163100 85500 163164
rect 95924 163100 95988 163164
rect 99420 163160 99484 163164
rect 99420 163104 99434 163160
rect 99434 163104 99484 163160
rect 99420 163100 99484 163104
rect 113588 163160 113652 163164
rect 113588 163104 113602 163160
rect 113602 163104 113652 163160
rect 113588 163100 113652 163104
rect 128308 163160 128372 163164
rect 128308 163104 128358 163160
rect 128358 163104 128372 163160
rect 128308 163100 128372 163104
rect 235948 163160 236012 163164
rect 235948 163104 235998 163160
rect 235998 163104 236012 163160
rect 235948 163100 236012 163104
rect 261708 163100 261772 163164
rect 54708 162692 54772 162756
rect 76052 162692 76116 162756
rect 78260 162692 78324 162756
rect 79548 162692 79612 162756
rect 80468 162692 80532 162756
rect 81940 162692 82004 162756
rect 83044 162692 83108 162756
rect 86540 162692 86604 162756
rect 87644 162692 87708 162756
rect 88748 162692 88812 162756
rect 90036 162692 90100 162756
rect 90772 162752 90836 162756
rect 90772 162696 90786 162752
rect 90786 162696 90836 162752
rect 90772 162692 90836 162696
rect 91324 162692 91388 162756
rect 93348 162692 93412 162756
rect 93716 162752 93780 162756
rect 93716 162696 93730 162752
rect 93730 162696 93780 162752
rect 93716 162692 93780 162696
rect 94452 162692 94516 162756
rect 97028 162692 97092 162756
rect 98132 162692 98196 162756
rect 100708 162752 100772 162756
rect 100708 162696 100758 162752
rect 100758 162696 100772 162752
rect 100708 162692 100772 162696
rect 102732 162692 102796 162756
rect 103836 162692 103900 162756
rect 105308 162692 105372 162756
rect 106412 162692 106476 162756
rect 108620 162692 108684 162756
rect 109540 162692 109604 162756
rect 111196 162692 111260 162756
rect 112116 162692 112180 162756
rect 113220 162692 113284 162756
rect 115796 162692 115860 162756
rect 115980 162752 116044 162756
rect 115980 162696 115994 162752
rect 115994 162696 116044 162752
rect 115980 162692 116044 162696
rect 118004 162692 118068 162756
rect 118372 162752 118436 162756
rect 118372 162696 118386 162752
rect 118386 162696 118436 162752
rect 118372 162692 118436 162696
rect 119108 162692 119172 162756
rect 120764 162752 120828 162756
rect 120764 162696 120778 162752
rect 120778 162696 120828 162752
rect 120764 162692 120828 162696
rect 122604 162692 122668 162756
rect 125916 162752 125980 162756
rect 125916 162696 125930 162752
rect 125930 162696 125980 162752
rect 125916 162692 125980 162696
rect 130884 162752 130948 162756
rect 130884 162696 130898 162752
rect 130898 162696 130948 162752
rect 130884 162692 130948 162696
rect 133460 162752 133524 162756
rect 133460 162696 133474 162752
rect 133474 162696 133524 162752
rect 133460 162692 133524 162696
rect 183508 162752 183572 162756
rect 183508 162696 183522 162752
rect 183522 162696 183572 162752
rect 183508 162692 183572 162696
rect 237052 162692 237116 162756
rect 238156 162692 238220 162756
rect 240548 162692 240612 162756
rect 241652 162692 241716 162756
rect 242940 162752 243004 162756
rect 242940 162696 242954 162752
rect 242954 162696 243004 162752
rect 242940 162692 243004 162696
rect 244228 162752 244292 162756
rect 244228 162696 244278 162752
rect 244278 162696 244292 162752
rect 244228 162692 244292 162696
rect 246436 162692 246500 162756
rect 247724 162692 247788 162756
rect 248276 162692 248340 162756
rect 248644 162692 248708 162756
rect 250116 162692 250180 162756
rect 251220 162752 251284 162756
rect 251220 162696 251270 162752
rect 251270 162696 251284 162752
rect 251220 162692 251284 162696
rect 253428 162692 253492 162756
rect 254532 162692 254596 162756
rect 255820 162692 255884 162756
rect 256004 162752 256068 162756
rect 256004 162696 256018 162752
rect 256018 162696 256068 162752
rect 256004 162692 256068 162696
rect 256924 162692 256988 162756
rect 259500 162752 259564 162756
rect 259500 162696 259550 162752
rect 259550 162696 259564 162752
rect 259500 162692 259564 162696
rect 265204 163100 265268 163164
rect 272196 163100 272260 163164
rect 325924 163100 325988 163164
rect 398236 163100 398300 163164
rect 262812 162692 262876 162756
rect 263916 162692 263980 162756
rect 265940 162692 266004 162756
rect 266308 162752 266372 162756
rect 266308 162696 266358 162752
rect 266358 162696 266372 162752
rect 266308 162692 266372 162696
rect 267596 162752 267660 162756
rect 267596 162696 267610 162752
rect 267610 162696 267660 162752
rect 267596 162692 267660 162696
rect 268700 162692 268764 162756
rect 269804 162692 269868 162756
rect 271092 162692 271156 162756
rect 274404 162692 274468 162756
rect 276980 162692 277044 162756
rect 278452 162752 278516 162756
rect 278452 162696 278466 162752
rect 278466 162696 278516 162752
rect 278452 162692 278516 162696
rect 279004 162692 279068 162756
rect 280844 162752 280908 162756
rect 280844 162696 280858 162752
rect 280858 162696 280908 162752
rect 280844 162692 280908 162696
rect 283788 162752 283852 162756
rect 283788 162696 283802 162752
rect 283802 162696 283852 162752
rect 283788 162692 283852 162696
rect 285996 162752 286060 162756
rect 285996 162696 286010 162752
rect 286010 162696 286060 162752
rect 285996 162692 286060 162696
rect 293356 162752 293420 162756
rect 293356 162696 293370 162752
rect 293370 162696 293420 162752
rect 293356 162692 293420 162696
rect 303476 162752 303540 162756
rect 303476 162696 303490 162752
rect 303490 162696 303540 162752
rect 303476 162692 303540 162696
rect 308628 162752 308692 162756
rect 308628 162696 308642 162752
rect 308642 162696 308692 162752
rect 308628 162692 308692 162696
rect 343404 162752 343468 162756
rect 343404 162696 343454 162752
rect 343454 162696 343468 162752
rect 158484 162556 158548 162620
rect 166028 162556 166092 162620
rect 198780 162556 198844 162620
rect 214788 162556 214852 162620
rect 155908 162420 155972 162484
rect 183140 162480 183204 162484
rect 183140 162424 183190 162480
rect 183190 162424 183204 162480
rect 183140 162420 183204 162424
rect 203196 162420 203260 162484
rect 136036 162284 136100 162348
rect 214972 162284 215036 162348
rect 250668 162284 250732 162348
rect 252324 162420 252388 162484
rect 260604 162556 260668 162620
rect 263548 162556 263612 162620
rect 268332 162616 268396 162620
rect 268332 162560 268346 162616
rect 268346 162560 268396 162616
rect 268332 162556 268396 162560
rect 273300 162556 273364 162620
rect 276244 162420 276308 162484
rect 253612 162284 253676 162348
rect 273484 162344 273548 162348
rect 273484 162288 273498 162344
rect 273498 162288 273548 162344
rect 273484 162284 273548 162288
rect 77156 162148 77220 162212
rect 88380 162208 88444 162212
rect 88380 162152 88394 162208
rect 88394 162152 88444 162208
rect 88380 162148 88444 162152
rect 91508 162148 91572 162212
rect 101812 162148 101876 162212
rect 107516 162148 107580 162212
rect 111012 162208 111076 162212
rect 111012 162152 111026 162208
rect 111026 162152 111076 162208
rect 111012 162148 111076 162152
rect 245332 162148 245396 162212
rect 258396 162148 258460 162212
rect 114508 162012 114572 162076
rect 196756 162012 196820 162076
rect 160876 161876 160940 161940
rect 200804 161876 200868 161940
rect 343404 162692 343468 162696
rect 396028 162752 396092 162756
rect 396028 162696 396078 162752
rect 396078 162696 396092 162752
rect 396028 162692 396092 162696
rect 401732 163100 401796 163164
rect 455828 163160 455892 163164
rect 455828 163104 455842 163160
rect 455842 163104 455892 163160
rect 455828 163100 455892 163104
rect 418108 162888 418172 162892
rect 418108 162832 418158 162888
rect 418158 162832 418172 162888
rect 418108 162828 418172 162832
rect 399524 162692 399588 162756
rect 400444 162692 400508 162756
rect 403020 162752 403084 162756
rect 403020 162696 403070 162752
rect 403070 162696 403084 162752
rect 403020 162692 403084 162696
rect 405044 162692 405108 162756
rect 406516 162692 406580 162756
rect 407620 162692 407684 162756
rect 408356 162752 408420 162756
rect 408356 162696 408370 162752
rect 408370 162696 408420 162752
rect 408356 162692 408420 162696
rect 408724 162692 408788 162756
rect 410012 162752 410076 162756
rect 410012 162696 410026 162752
rect 410026 162696 410076 162752
rect 410012 162692 410076 162696
rect 410748 162692 410812 162756
rect 411300 162752 411364 162756
rect 411300 162696 411350 162752
rect 411350 162696 411364 162752
rect 411300 162692 411364 162696
rect 413508 162692 413572 162756
rect 413692 162752 413756 162756
rect 413692 162696 413706 162752
rect 413706 162696 413756 162752
rect 413692 162692 413756 162696
rect 414612 162692 414676 162756
rect 415532 162692 415596 162756
rect 417004 162692 417068 162756
rect 419212 162692 419276 162756
rect 420684 162692 420748 162756
rect 421788 162692 421852 162756
rect 422892 162692 422956 162756
rect 423996 162692 424060 162756
rect 425284 162692 425348 162756
rect 426388 162752 426452 162756
rect 426388 162696 426438 162752
rect 426438 162696 426452 162752
rect 426388 162692 426452 162696
rect 428780 162692 428844 162756
rect 429700 162692 429764 162756
rect 431172 162692 431236 162756
rect 431724 162692 431788 162756
rect 433380 162692 433444 162756
rect 435772 162692 435836 162756
rect 435956 162752 436020 162756
rect 435956 162696 435970 162752
rect 435970 162696 436020 162752
rect 435956 162692 436020 162696
rect 438532 162752 438596 162756
rect 438532 162696 438546 162752
rect 438546 162696 438596 162752
rect 438532 162692 438596 162696
rect 439084 162752 439148 162756
rect 439084 162696 439098 162752
rect 439098 162696 439148 162752
rect 439084 162692 439148 162696
rect 440924 162752 440988 162756
rect 440924 162696 440938 162752
rect 440938 162696 440988 162752
rect 440924 162692 440988 162696
rect 443500 162752 443564 162756
rect 443500 162696 443514 162752
rect 443514 162696 443564 162752
rect 443500 162692 443564 162696
rect 445892 162752 445956 162756
rect 445892 162696 445906 162752
rect 445906 162696 445956 162752
rect 445892 162692 445956 162696
rect 448284 162752 448348 162756
rect 448284 162696 448298 162752
rect 448298 162696 448348 162752
rect 448284 162692 448348 162696
rect 453436 162692 453500 162756
rect 458404 162752 458468 162756
rect 458404 162696 458418 162752
rect 458418 162696 458468 162752
rect 458404 162692 458468 162696
rect 503116 162692 503180 162756
rect 320956 162616 321020 162620
rect 320956 162560 320970 162616
rect 320970 162560 321020 162616
rect 320956 162556 321020 162560
rect 343220 162556 343284 162620
rect 465948 162556 466012 162620
rect 503484 162556 503548 162620
rect 462636 162420 462700 162484
rect 460980 162284 461044 162348
rect 397132 162148 397196 162212
rect 404124 162148 404188 162212
rect 412404 162148 412468 162212
rect 418476 162208 418540 162212
rect 418476 162152 418490 162208
rect 418490 162152 418540 162208
rect 418476 162148 418540 162152
rect 427676 162148 427740 162212
rect 433564 162208 433628 162212
rect 433564 162152 433578 162208
rect 433578 162152 433628 162208
rect 433564 162148 433628 162152
rect 468524 161876 468588 161940
rect 84148 161468 84212 161532
rect 238708 161528 238772 161532
rect 238708 161472 238758 161528
rect 238758 161472 238772 161528
rect 238708 161468 238772 161472
rect 277348 161468 277412 161532
rect 57652 160108 57716 160172
rect 377260 158748 377324 158812
rect 360700 149092 360764 149156
rect 217364 148276 217428 148340
rect 217180 146372 217244 146436
rect 377996 146236 378060 146300
rect 510844 146100 510908 146164
rect 57468 145964 57532 146028
rect 217548 145964 217612 146028
rect 190868 145420 190932 145484
rect 178540 144876 178604 144940
rect 179644 144936 179708 144940
rect 179644 144880 179694 144936
rect 179694 144880 179708 144936
rect 179644 144876 179708 144880
rect 338436 144936 338500 144940
rect 338436 144880 338486 144936
rect 338486 144880 338500 144936
rect 338436 144876 338500 144880
rect 339724 144876 339788 144940
rect 350948 144876 351012 144940
rect 498516 144876 498580 144940
rect 499804 144936 499868 144940
rect 499804 144880 499854 144936
rect 499854 144880 499868 144936
rect 499804 144876 499868 144880
rect 57100 144740 57164 144804
rect 57468 144740 57532 144804
rect 377444 143652 377508 143716
rect 57468 140796 57532 140860
rect 57836 70348 57900 70412
rect 208900 69940 208964 70004
rect 46796 67764 46860 67828
rect 206140 68036 206204 68100
rect 218652 60556 218716 60620
rect 219204 60616 219268 60620
rect 219204 60560 219254 60616
rect 219254 60560 219268 60616
rect 219204 60556 219268 60560
rect 77142 59800 77206 59804
rect 77142 59744 77170 59800
rect 77170 59744 77206 59800
rect 77142 59740 77206 59744
rect 83126 59800 83190 59804
rect 83126 59744 83150 59800
rect 83150 59744 83190 59800
rect 83126 59740 83190 59744
rect 99446 59800 99510 59804
rect 99446 59744 99470 59800
rect 99470 59744 99510 59800
rect 99446 59740 99510 59744
rect 113590 59800 113654 59804
rect 113590 59744 113602 59800
rect 113602 59744 113654 59800
rect 113590 59740 113654 59744
rect 120934 59800 120998 59804
rect 120934 59744 120962 59800
rect 120962 59744 120998 59800
rect 120934 59740 120998 59744
rect 237142 59800 237206 59804
rect 237142 59744 237158 59800
rect 237158 59744 237206 59800
rect 237142 59740 237206 59744
rect 255910 59800 255974 59804
rect 255910 59744 255926 59800
rect 255926 59744 255974 59800
rect 255910 59740 255974 59744
rect 259446 59800 259510 59804
rect 259446 59744 259458 59800
rect 259458 59744 259510 59800
rect 259446 59740 259510 59744
rect 260670 59800 260734 59804
rect 260670 59744 260710 59800
rect 260710 59744 260734 59800
rect 260670 59740 260734 59744
rect 261758 59800 261822 59804
rect 261758 59744 261814 59800
rect 261814 59744 261822 59800
rect 261758 59740 261822 59744
rect 263934 59740 263998 59804
rect 396054 59800 396118 59804
rect 396054 59744 396078 59800
rect 396078 59744 396118 59800
rect 396054 59740 396118 59744
rect 397142 59800 397206 59804
rect 397142 59744 397146 59800
rect 397146 59744 397206 59800
rect 397142 59740 397206 59744
rect 416998 59800 417062 59804
rect 416998 59744 417018 59800
rect 417018 59744 417062 59800
rect 416998 59740 417062 59744
rect 418494 59740 418558 59804
rect 422846 59800 422910 59804
rect 422846 59744 422850 59800
rect 422850 59744 422906 59800
rect 422906 59744 422910 59800
rect 422846 59740 422910 59744
rect 423934 59800 423998 59804
rect 423934 59744 423954 59800
rect 423954 59744 423998 59800
rect 423934 59740 423998 59744
rect 94550 59664 94614 59668
rect 94550 59608 94558 59664
rect 94558 59608 94614 59664
rect 94550 59604 94614 59608
rect 102846 59604 102910 59668
rect 105974 59604 106038 59668
rect 113318 59664 113382 59668
rect 113318 59608 113326 59664
rect 113326 59608 113382 59664
rect 113318 59604 113382 59608
rect 116990 59664 117054 59668
rect 116990 59608 117006 59664
rect 117006 59608 117054 59664
rect 116990 59604 117054 59608
rect 256998 59664 257062 59668
rect 256998 59608 257030 59664
rect 257030 59608 257062 59664
rect 256998 59604 257062 59608
rect 258086 59664 258150 59668
rect 258086 59608 258134 59664
rect 258134 59608 258150 59664
rect 258086 59604 258150 59608
rect 265294 59664 265358 59668
rect 265294 59608 265310 59664
rect 265310 59608 265358 59664
rect 265294 59604 265358 59608
rect 315886 59664 315950 59668
rect 315886 59608 315910 59664
rect 315910 59608 315950 59664
rect 315886 59604 315950 59608
rect 403126 59604 403190 59668
rect 404214 59664 404278 59668
rect 404214 59608 404230 59664
rect 404230 59608 404278 59664
rect 404214 59604 404278 59608
rect 46612 59468 46676 59532
rect 413462 59604 413526 59668
rect 423526 59664 423590 59668
rect 423526 59608 423550 59664
rect 423550 59608 423590 59664
rect 423526 59604 423590 59608
rect 480918 59664 480982 59668
rect 480918 59608 480958 59664
rect 480958 59608 480982 59664
rect 480918 59604 480982 59608
rect 262812 59528 262876 59532
rect 262812 59472 262826 59528
rect 262826 59472 262876 59528
rect 262812 59468 262876 59472
rect 418108 59528 418172 59532
rect 418108 59472 418158 59528
rect 418158 59472 418172 59528
rect 418108 59468 418172 59472
rect 95924 59392 95988 59396
rect 95924 59336 95938 59392
rect 95938 59336 95988 59392
rect 95924 59332 95988 59336
rect 98132 59392 98196 59396
rect 98132 59336 98146 59392
rect 98146 59336 98196 59392
rect 98132 59332 98196 59336
rect 100708 59392 100772 59396
rect 100708 59336 100758 59392
rect 100758 59336 100772 59392
rect 100708 59332 100772 59336
rect 101812 59392 101876 59396
rect 101812 59336 101826 59392
rect 101826 59336 101876 59392
rect 101812 59332 101876 59336
rect 197860 59332 197924 59396
rect 263548 59332 263612 59396
rect 420684 59392 420748 59396
rect 420684 59336 420698 59392
rect 420698 59336 420748 59392
rect 420684 59332 420748 59336
rect 421788 59392 421852 59396
rect 421788 59336 421802 59392
rect 421802 59336 421852 59392
rect 421788 59332 421852 59336
rect 426020 59392 426084 59396
rect 426020 59336 426034 59392
rect 426034 59336 426084 59392
rect 426020 59332 426084 59336
rect 428228 59392 428292 59396
rect 428228 59336 428242 59392
rect 428242 59336 428292 59392
rect 428228 59332 428292 59336
rect 453436 59392 453500 59396
rect 453436 59336 453450 59392
rect 453450 59336 453500 59392
rect 453436 59332 453500 59336
rect 463556 59392 463620 59396
rect 463556 59336 463570 59392
rect 463570 59336 463620 59392
rect 463556 59332 463620 59336
rect 52132 59196 52196 59260
rect 143580 59196 143644 59260
rect 148548 59256 148612 59260
rect 148548 59200 148562 59256
rect 148562 59200 148612 59256
rect 148548 59196 148612 59200
rect 150940 59256 151004 59260
rect 150940 59200 150954 59256
rect 150954 59200 151004 59256
rect 150940 59196 151004 59200
rect 202644 59196 202708 59260
rect 285996 59196 286060 59260
rect 295932 59256 295996 59260
rect 295932 59200 295946 59256
rect 295946 59200 295996 59256
rect 295932 59196 295996 59200
rect 298508 59256 298572 59260
rect 298508 59200 298522 59256
rect 298522 59200 298572 59256
rect 298508 59196 298572 59200
rect 303476 59256 303540 59260
rect 303476 59200 303490 59256
rect 303490 59200 303540 59256
rect 303476 59196 303540 59200
rect 323348 59256 323412 59260
rect 323348 59200 323362 59256
rect 323362 59200 323412 59256
rect 323348 59196 323412 59200
rect 357940 59196 358004 59260
rect 483428 59196 483492 59260
rect 486004 59256 486068 59260
rect 486004 59200 486018 59256
rect 486018 59200 486068 59256
rect 486004 59196 486068 59200
rect 54892 59060 54956 59124
rect 140820 59060 140884 59124
rect 198596 59060 198660 59124
rect 280844 59060 280908 59124
rect 367692 59060 367756 59124
rect 468524 59060 468588 59124
rect 53420 58924 53484 58988
rect 138428 58924 138492 58988
rect 210740 58924 210804 58988
rect 290964 58924 291028 58988
rect 374500 58924 374564 58988
rect 473492 58924 473556 58988
rect 51948 58788 52012 58852
rect 135852 58788 135916 58852
rect 201356 58788 201420 58852
rect 273484 58788 273548 58852
rect 375972 58788 376036 58852
rect 475884 58788 475948 58852
rect 48084 58652 48148 58716
rect 108252 58652 108316 58716
rect 209636 58652 209700 58716
rect 276060 58652 276124 58716
rect 371740 58652 371804 58716
rect 458404 58652 458468 58716
rect 52316 58516 52380 58580
rect 111012 58516 111076 58580
rect 202092 58516 202156 58580
rect 268332 58516 268396 58580
rect 377996 58516 378060 58580
rect 425284 58516 425348 58580
rect 59308 58380 59372 58444
rect 101076 58380 101140 58444
rect 200620 58380 200684 58444
rect 256004 58380 256068 58444
rect 377260 58380 377324 58444
rect 419396 58380 419460 58444
rect 85436 58108 85500 58172
rect 92244 58108 92308 58172
rect 128308 58108 128372 58172
rect 153332 58108 153396 58172
rect 235948 58108 236012 58172
rect 272196 58108 272260 58172
rect 275692 58108 275756 58172
rect 300900 58108 300964 58172
rect 325924 58168 325988 58172
rect 325924 58112 325938 58168
rect 325938 58112 325988 58168
rect 325924 58108 325988 58112
rect 398236 58108 398300 58172
rect 401732 58108 401796 58172
rect 405412 58108 405476 58172
rect 416084 58108 416148 58172
rect 83964 57972 84028 58036
rect 76052 57896 76116 57900
rect 76052 57840 76066 57896
rect 76066 57840 76116 57896
rect 76052 57836 76116 57840
rect 78260 57896 78324 57900
rect 78260 57840 78274 57896
rect 78274 57840 78324 57896
rect 78260 57836 78324 57840
rect 79548 57896 79612 57900
rect 79548 57840 79562 57896
rect 79562 57840 79612 57896
rect 79548 57836 79612 57840
rect 80468 57836 80532 57900
rect 81940 57836 82004 57900
rect 86540 57896 86604 57900
rect 86540 57840 86554 57896
rect 86554 57840 86604 57896
rect 86540 57836 86604 57840
rect 87644 57836 87708 57900
rect 88380 57896 88444 57900
rect 88380 57840 88394 57896
rect 88394 57840 88444 57896
rect 88380 57836 88444 57840
rect 88748 57896 88812 57900
rect 88748 57840 88762 57896
rect 88762 57840 88812 57896
rect 88748 57836 88812 57840
rect 90036 57836 90100 57900
rect 90772 57896 90836 57900
rect 90772 57840 90786 57896
rect 90786 57840 90836 57896
rect 90772 57836 90836 57840
rect 91324 57836 91388 57900
rect 93348 57836 93412 57900
rect 103836 57896 103900 57900
rect 103836 57840 103850 57896
rect 103850 57840 103900 57896
rect 103836 57836 103900 57840
rect 105308 57836 105372 57900
rect 106412 57896 106476 57900
rect 106412 57840 106426 57896
rect 106426 57840 106476 57896
rect 106412 57836 106476 57840
rect 107516 57836 107580 57900
rect 108620 57836 108684 57900
rect 109540 57836 109604 57900
rect 111196 57896 111260 57900
rect 111196 57840 111210 57896
rect 111210 57840 111260 57896
rect 111196 57836 111260 57840
rect 115796 57896 115860 57900
rect 115796 57840 115810 57896
rect 115810 57840 115860 57896
rect 115796 57836 115860 57840
rect 123524 57896 123588 57900
rect 123524 57840 123538 57896
rect 123538 57840 123588 57896
rect 123524 57836 123588 57840
rect 125916 57896 125980 57900
rect 125916 57840 125930 57896
rect 125930 57840 125980 57896
rect 125916 57836 125980 57840
rect 130884 57896 130948 57900
rect 130884 57840 130898 57896
rect 130898 57840 130948 57896
rect 130884 57836 130948 57840
rect 133460 57896 133524 57900
rect 133460 57840 133474 57896
rect 133474 57840 133524 57896
rect 133460 57836 133524 57840
rect 145604 57896 145668 57900
rect 145604 57840 145618 57896
rect 145618 57840 145668 57896
rect 145604 57836 145668 57840
rect 183140 57836 183204 57900
rect 238156 57836 238220 57900
rect 239260 57896 239324 57900
rect 239260 57840 239274 57896
rect 239274 57840 239324 57896
rect 239260 57836 239324 57840
rect 242940 57896 243004 57900
rect 242940 57840 242954 57896
rect 242954 57840 243004 57896
rect 242940 57836 243004 57840
rect 245332 57836 245396 57900
rect 246436 57896 246500 57900
rect 246436 57840 246450 57896
rect 246450 57840 246500 57896
rect 246436 57836 246500 57840
rect 248644 57896 248708 57900
rect 248644 57840 248658 57896
rect 248658 57840 248708 57896
rect 248644 57836 248708 57840
rect 251220 57896 251284 57900
rect 251220 57840 251234 57896
rect 251234 57840 251284 57896
rect 251220 57836 251284 57840
rect 253428 57896 253492 57900
rect 253428 57840 253442 57896
rect 253442 57840 253492 57896
rect 253428 57836 253492 57840
rect 265940 57836 266004 57900
rect 266308 57896 266372 57900
rect 266308 57840 266358 57896
rect 266358 57840 266372 57896
rect 266308 57836 266372 57840
rect 267596 57836 267660 57900
rect 269804 57896 269868 57900
rect 269804 57840 269818 57896
rect 269818 57840 269868 57896
rect 269804 57836 269868 57840
rect 274404 57836 274468 57900
rect 279004 57896 279068 57900
rect 279004 57840 279054 57896
rect 279054 57840 279068 57896
rect 279004 57836 279068 57840
rect 283788 57836 283852 57900
rect 288204 57836 288268 57900
rect 293356 57896 293420 57900
rect 293356 57840 293370 57896
rect 293370 57840 293420 57896
rect 293356 57836 293420 57840
rect 305868 57896 305932 57900
rect 305868 57840 305882 57896
rect 305882 57840 305932 57896
rect 305868 57836 305932 57840
rect 311020 57896 311084 57900
rect 311020 57840 311034 57896
rect 311034 57840 311084 57896
rect 311020 57836 311084 57840
rect 313412 57896 313476 57900
rect 313412 57840 313426 57896
rect 313426 57840 313476 57896
rect 313412 57836 313476 57840
rect 318380 57896 318444 57900
rect 318380 57840 318394 57896
rect 318394 57840 318444 57896
rect 318380 57836 318444 57840
rect 320956 57896 321020 57900
rect 320956 57840 320970 57896
rect 320970 57840 321020 57896
rect 320956 57836 321020 57840
rect 343220 57896 343284 57900
rect 343220 57840 343234 57896
rect 343234 57840 343284 57896
rect 343220 57836 343284 57840
rect 343404 57896 343468 57900
rect 343404 57840 343454 57896
rect 343454 57840 343468 57896
rect 343404 57836 343468 57840
rect 399524 57896 399588 57900
rect 399524 57840 399538 57896
rect 399538 57840 399588 57896
rect 399524 57836 399588 57840
rect 400444 57836 400508 57900
rect 406516 57836 406580 57900
rect 407620 57836 407684 57900
rect 408356 57896 408420 57900
rect 408356 57840 408370 57896
rect 408370 57840 408420 57896
rect 408356 57836 408420 57840
rect 408724 57896 408788 57900
rect 408724 57840 408738 57896
rect 408738 57840 408788 57896
rect 408724 57836 408788 57840
rect 410012 57836 410076 57900
rect 412404 57836 412468 57900
rect 414612 57896 414676 57900
rect 414612 57840 414626 57896
rect 414626 57840 414676 57896
rect 414612 57836 414676 57840
rect 415532 57896 415596 57900
rect 415532 57840 415546 57896
rect 415546 57840 415596 57896
rect 415532 57836 415596 57840
rect 426388 57896 426452 57900
rect 426388 57840 426438 57896
rect 426438 57840 426452 57896
rect 426388 57836 426452 57840
rect 427676 57896 427740 57900
rect 427676 57840 427690 57896
rect 427690 57840 427740 57896
rect 427676 57836 427740 57840
rect 428596 57836 428660 57900
rect 429700 57836 429764 57900
rect 431172 57836 431236 57900
rect 432276 57896 432340 57900
rect 432276 57840 432290 57896
rect 432290 57840 432340 57896
rect 432276 57836 432340 57840
rect 433380 57896 433444 57900
rect 433380 57840 433394 57896
rect 433394 57840 433444 57896
rect 433380 57836 433444 57840
rect 433564 57896 433628 57900
rect 433564 57840 433614 57896
rect 433614 57840 433628 57896
rect 433564 57836 433628 57840
rect 435956 57896 436020 57900
rect 435956 57840 435970 57896
rect 435970 57840 436020 57896
rect 435956 57836 436020 57840
rect 436876 57836 436940 57900
rect 438348 57836 438412 57900
rect 438532 57896 438596 57900
rect 438532 57840 438546 57896
rect 438546 57840 438596 57896
rect 438532 57836 438596 57840
rect 439084 57836 439148 57900
rect 440924 57896 440988 57900
rect 440924 57840 440938 57896
rect 440938 57840 440988 57896
rect 440924 57836 440988 57840
rect 443500 57896 443564 57900
rect 443500 57840 443514 57896
rect 443514 57840 443564 57896
rect 443500 57836 443564 57840
rect 448284 57896 448348 57900
rect 448284 57840 448298 57896
rect 448298 57840 448348 57896
rect 448284 57836 448348 57840
rect 470916 57896 470980 57900
rect 470916 57840 470930 57896
rect 470930 57840 470980 57896
rect 470916 57836 470980 57840
rect 478460 57896 478524 57900
rect 478460 57840 478474 57896
rect 478474 57840 478524 57896
rect 478460 57836 478524 57840
rect 503116 57836 503180 57900
rect 503484 57896 503548 57900
rect 503484 57840 503534 57896
rect 503534 57840 503548 57896
rect 503484 57836 503548 57840
rect 57652 57700 57716 57764
rect 44956 57564 45020 57628
rect 98500 57564 98564 57628
rect 118004 57700 118068 57764
rect 183508 57760 183572 57764
rect 183508 57704 183522 57760
rect 183522 57704 183572 57760
rect 183508 57700 183572 57704
rect 211660 57700 211724 57764
rect 270908 57700 270972 57764
rect 358124 57700 358188 57764
rect 451044 57700 451108 57764
rect 112116 57564 112180 57628
rect 114324 57564 114388 57628
rect 115980 57624 116044 57628
rect 115980 57568 115994 57624
rect 115994 57568 116044 57624
rect 115980 57564 116044 57568
rect 119108 57564 119172 57628
rect 155908 57624 155972 57628
rect 155908 57568 155958 57624
rect 155958 57568 155972 57624
rect 155908 57564 155972 57568
rect 160876 57564 160940 57628
rect 165844 57564 165908 57628
rect 204852 57564 204916 57628
rect 260972 57564 261036 57628
rect 268700 57564 268764 57628
rect 271092 57564 271156 57628
rect 273300 57624 273364 57628
rect 273300 57568 273350 57624
rect 273350 57568 273364 57624
rect 273300 57564 273364 57568
rect 278084 57564 278148 57628
rect 308628 57564 308692 57628
rect 376156 57564 376220 57628
rect 460980 57564 461044 57628
rect 58756 57428 58820 57492
rect 103836 57428 103900 57492
rect 214420 57428 214484 57492
rect 57100 57292 57164 57356
rect 97028 57292 97092 57356
rect 205036 57292 205100 57356
rect 240548 57428 240612 57492
rect 241652 57428 241716 57492
rect 244228 57488 244292 57492
rect 244228 57432 244278 57488
rect 244278 57432 244292 57488
rect 244228 57428 244292 57432
rect 247724 57428 247788 57492
rect 250116 57428 250180 57492
rect 252324 57428 252388 57492
rect 254532 57428 254596 57492
rect 364932 57428 364996 57492
rect 445892 57428 445956 57492
rect 258396 57292 258460 57356
rect 378916 57292 378980 57356
rect 456380 57292 456444 57356
rect 59124 57156 59188 57220
rect 96292 57156 96356 57220
rect 215892 57156 215956 57220
rect 253612 57156 253676 57220
rect 379100 57156 379164 57220
rect 421052 57156 421116 57220
rect 430988 57216 431052 57220
rect 430988 57160 431002 57216
rect 431002 57160 431052 57216
rect 430988 57156 431052 57160
rect 434668 57156 434732 57220
rect 435772 57216 435836 57220
rect 435772 57160 435786 57216
rect 435786 57160 435836 57216
rect 435772 57156 435836 57160
rect 58940 57020 59004 57084
rect 93716 57020 93780 57084
rect 214604 57020 214668 57084
rect 250668 57020 250732 57084
rect 378732 57020 378796 57084
rect 413508 57020 413572 57084
rect 248276 56884 248340 56948
rect 411300 56944 411364 56948
rect 411300 56888 411314 56944
rect 411314 56888 411364 56944
rect 411300 56884 411364 56888
rect 55076 56612 55140 56676
rect 118372 56612 118436 56676
rect 163268 56612 163332 56676
rect 202276 56612 202340 56676
rect 278452 56748 278516 56812
rect 370452 56612 370516 56676
rect 465948 56612 466012 56676
rect 53604 56476 53668 56540
rect 219940 56476 220004 56540
rect 410748 56476 410812 56540
rect 48636 56340 48700 56404
rect 158484 56340 158548 56404
rect 217180 56340 217244 56404
rect 276980 56340 277044 56404
rect 55628 56204 55692 56268
rect 50476 55116 50540 55180
rect 205220 55116 205284 55180
rect 377444 55116 377508 55180
rect 50660 54980 50724 55044
rect 217364 54980 217428 55044
rect 50844 54844 50908 54908
rect 217548 54844 217612 54908
rect 57468 54708 57532 54772
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 53051 630868 53117 630869
rect 53051 630804 53052 630868
rect 53116 630804 53117 630868
rect 53051 630803 53117 630804
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 45234 478574 45854 478658
rect 46795 478684 46861 478685
rect 46795 478620 46796 478684
rect 46860 478620 46861 478684
rect 46795 478619 46861 478620
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 44955 460188 45021 460189
rect 44955 460124 44956 460188
rect 45020 460124 45021 460188
rect 44955 460123 45021 460124
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 44958 57629 45018 460123
rect 45234 442894 45854 478338
rect 46611 460460 46677 460461
rect 46611 460396 46612 460460
rect 46676 460396 46677 460460
rect 46611 460395 46677 460396
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 44955 57628 45021 57629
rect 44955 57564 44956 57628
rect 45020 57564 45021 57628
rect 44955 57563 45021 57564
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 46894 45854 82338
rect 46614 59533 46674 460395
rect 46798 67829 46858 478619
rect 47899 475420 47965 475421
rect 47899 475356 47900 475420
rect 47964 475356 47965 475420
rect 47899 475355 47965 475356
rect 47902 264893 47962 475355
rect 48083 463180 48149 463181
rect 48083 463116 48084 463180
rect 48148 463116 48149 463180
rect 48083 463115 48149 463116
rect 47899 264892 47965 264893
rect 47899 264828 47900 264892
rect 47964 264828 47965 264892
rect 47899 264827 47965 264828
rect 46795 67828 46861 67829
rect 46795 67764 46796 67828
rect 46860 67764 46861 67828
rect 46795 67763 46861 67764
rect 46611 59532 46677 59533
rect 46611 59468 46612 59532
rect 46676 59468 46677 59532
rect 46611 59467 46677 59468
rect 48086 58717 48146 463115
rect 48635 459644 48701 459645
rect 48635 459580 48636 459644
rect 48700 459580 48701 459644
rect 48635 459579 48701 459580
rect 48083 58716 48149 58717
rect 48083 58652 48084 58716
rect 48148 58652 48149 58716
rect 48083 58651 48149 58652
rect 48638 56405 48698 459579
rect 48954 446614 49574 482058
rect 50659 477732 50725 477733
rect 50659 477668 50660 477732
rect 50724 477668 50725 477732
rect 50659 477667 50725 477668
rect 50475 463044 50541 463045
rect 50475 462980 50476 463044
rect 50540 462980 50541 463044
rect 50475 462979 50541 462980
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48635 56404 48701 56405
rect 48635 56340 48636 56404
rect 48700 56340 48701 56404
rect 48635 56339 48701 56340
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 50614 49574 86058
rect 50478 55181 50538 462979
rect 50475 55180 50541 55181
rect 50475 55116 50476 55180
rect 50540 55116 50541 55180
rect 50475 55115 50541 55116
rect 50662 55045 50722 477667
rect 50843 477596 50909 477597
rect 50843 477532 50844 477596
rect 50908 477532 50909 477596
rect 50843 477531 50909 477532
rect 50659 55044 50725 55045
rect 50659 54980 50660 55044
rect 50724 54980 50725 55044
rect 50659 54979 50725 54980
rect 50846 54909 50906 477531
rect 52315 463452 52381 463453
rect 52315 463388 52316 463452
rect 52380 463388 52381 463452
rect 52315 463387 52381 463388
rect 51947 460324 52013 460325
rect 51947 460260 51948 460324
rect 52012 460260 52013 460324
rect 51947 460259 52013 460260
rect 51579 459644 51645 459645
rect 51579 459580 51580 459644
rect 51644 459580 51645 459644
rect 51579 459579 51645 459580
rect 51582 383621 51642 459579
rect 51579 383620 51645 383621
rect 51579 383556 51580 383620
rect 51644 383556 51645 383620
rect 51579 383555 51645 383556
rect 51950 58853 52010 460259
rect 52131 459644 52197 459645
rect 52131 459580 52132 459644
rect 52196 459580 52197 459644
rect 52131 459579 52197 459580
rect 52134 59261 52194 459579
rect 52131 59260 52197 59261
rect 52131 59196 52132 59260
rect 52196 59196 52197 59260
rect 52131 59195 52197 59196
rect 51947 58852 52013 58853
rect 51947 58788 51948 58852
rect 52012 58788 52013 58852
rect 51947 58787 52013 58788
rect 52318 58581 52378 463387
rect 53054 254013 53114 630803
rect 54339 630732 54405 630733
rect 54339 630668 54340 630732
rect 54404 630668 54405 630732
rect 54339 630667 54405 630668
rect 53235 478548 53301 478549
rect 53235 478484 53236 478548
rect 53300 478484 53301 478548
rect 53235 478483 53301 478484
rect 53238 375325 53298 478483
rect 53419 460596 53485 460597
rect 53419 460532 53420 460596
rect 53484 460532 53485 460596
rect 53419 460531 53485 460532
rect 53235 375324 53301 375325
rect 53235 375260 53236 375324
rect 53300 375260 53301 375324
rect 53235 375259 53301 375260
rect 53051 254012 53117 254013
rect 53051 253948 53052 254012
rect 53116 253948 53117 254012
rect 53051 253947 53117 253948
rect 53422 58989 53482 460531
rect 53603 459644 53669 459645
rect 53603 459580 53604 459644
rect 53668 459580 53669 459644
rect 53603 459579 53669 459580
rect 53419 58988 53485 58989
rect 53419 58924 53420 58988
rect 53484 58924 53485 58988
rect 53419 58923 53485 58924
rect 52315 58580 52381 58581
rect 52315 58516 52316 58580
rect 52380 58516 52381 58580
rect 52315 58515 52381 58516
rect 53606 56541 53666 459579
rect 54342 305013 54402 630667
rect 55794 597454 56414 632898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 625099 60134 636618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 625099 63854 640338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 625099 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 625099 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 625099 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 625099 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 625099 85574 626058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 625099 92414 632898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 625099 96134 636618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 625099 99854 640338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 625099 103574 644058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 625099 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 625099 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 625099 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120027 625292 120093 625293
rect 120027 625228 120028 625292
rect 120092 625228 120093 625292
rect 120027 625227 120093 625228
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 79568 597454 79888 597486
rect 79568 597218 79610 597454
rect 79846 597218 79888 597454
rect 79568 597134 79888 597218
rect 79568 596898 79610 597134
rect 79846 596898 79888 597134
rect 79568 596866 79888 596898
rect 110288 597454 110608 597486
rect 110288 597218 110330 597454
rect 110566 597218 110608 597454
rect 110288 597134 110608 597218
rect 110288 596898 110330 597134
rect 110566 596898 110608 597134
rect 110288 596866 110608 596898
rect 64208 579454 64528 579486
rect 64208 579218 64250 579454
rect 64486 579218 64528 579454
rect 64208 579134 64528 579218
rect 64208 578898 64250 579134
rect 64486 578898 64528 579134
rect 64208 578866 64528 578898
rect 94928 579454 95248 579486
rect 94928 579218 94970 579454
rect 95206 579218 95248 579454
rect 94928 579134 95248 579218
rect 94928 578898 94970 579134
rect 95206 578898 95248 579134
rect 94928 578866 95248 578898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 120030 559605 120090 625227
rect 120954 625099 121574 626058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 120027 559604 120093 559605
rect 120027 559540 120028 559604
rect 120092 559540 120093 559604
rect 120027 559539 120093 559540
rect 59514 548114 60134 558000
rect 59514 547878 59546 548114
rect 59782 547878 59866 548114
rect 60102 547878 60134 548114
rect 59514 547794 60134 547878
rect 59514 547558 59546 547794
rect 59782 547558 59866 547794
rect 60102 547558 60134 547794
rect 59514 542000 60134 547558
rect 63234 549954 63854 558000
rect 63234 549718 63266 549954
rect 63502 549718 63586 549954
rect 63822 549718 63854 549954
rect 63234 549634 63854 549718
rect 63234 549398 63266 549634
rect 63502 549398 63586 549634
rect 63822 549398 63854 549634
rect 63234 542000 63854 549398
rect 66954 553674 67574 558000
rect 66954 553438 66986 553674
rect 67222 553438 67306 553674
rect 67542 553438 67574 553674
rect 66954 553354 67574 553438
rect 66954 553118 66986 553354
rect 67222 553118 67306 553354
rect 67542 553118 67574 553354
rect 66954 542000 67574 553118
rect 73794 543454 74414 558000
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 542000 74414 542898
rect 77514 547174 78134 558000
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 542000 78134 546618
rect 81234 550894 81854 558000
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 542000 81854 550338
rect 84954 554614 85574 558000
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 542000 85574 554058
rect 91794 544394 92414 558000
rect 91794 544158 91826 544394
rect 92062 544158 92146 544394
rect 92382 544158 92414 544394
rect 91794 544074 92414 544158
rect 91794 543838 91826 544074
rect 92062 543838 92146 544074
rect 92382 543838 92414 544074
rect 91794 542000 92414 543838
rect 95514 548114 96134 558000
rect 95514 547878 95546 548114
rect 95782 547878 95866 548114
rect 96102 547878 96134 548114
rect 95514 547794 96134 547878
rect 95514 547558 95546 547794
rect 95782 547558 95866 547794
rect 96102 547558 96134 547794
rect 95514 542000 96134 547558
rect 99234 549954 99854 558000
rect 99234 549718 99266 549954
rect 99502 549718 99586 549954
rect 99822 549718 99854 549954
rect 99234 549634 99854 549718
rect 99234 549398 99266 549634
rect 99502 549398 99586 549634
rect 99822 549398 99854 549634
rect 99234 542000 99854 549398
rect 102954 553674 103574 558000
rect 102954 553438 102986 553674
rect 103222 553438 103306 553674
rect 103542 553438 103574 553674
rect 102954 553354 103574 553438
rect 102954 553118 102986 553354
rect 103222 553118 103306 553354
rect 103542 553118 103574 553354
rect 102954 542000 103574 553118
rect 109794 543454 110414 558000
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 542000 110414 542898
rect 113514 547174 114134 558000
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 542000 114134 546618
rect 117234 550894 117854 558000
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 542000 117854 550338
rect 120954 554614 121574 558000
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 542000 121574 554058
rect 127794 544394 128414 560898
rect 127794 544158 127826 544394
rect 128062 544158 128146 544394
rect 128382 544158 128414 544394
rect 127794 544074 128414 544158
rect 127794 543838 127826 544074
rect 128062 543838 128146 544074
rect 128382 543838 128414 544074
rect 127794 542000 128414 543838
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 548114 132134 564618
rect 131514 547878 131546 548114
rect 131782 547878 131866 548114
rect 132102 547878 132134 548114
rect 131514 547794 132134 547878
rect 131514 547558 131546 547794
rect 131782 547558 131866 547794
rect 132102 547558 132134 547794
rect 131514 542000 132134 547558
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 625099 139574 644058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 625099 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 625099 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 625099 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 625099 157574 626058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 625099 164414 632898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 625099 168134 636618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 625099 171854 640338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 625099 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 625099 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 625099 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 625099 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 625099 193574 626058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 625099 200414 632898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 144208 615454 144528 615486
rect 144208 615218 144250 615454
rect 144486 615218 144528 615454
rect 144208 615134 144528 615218
rect 144208 614898 144250 615134
rect 144486 614898 144528 615134
rect 144208 614866 144528 614898
rect 174928 615454 175248 615486
rect 174928 615218 174970 615454
rect 175206 615218 175248 615454
rect 174928 615134 175248 615218
rect 174928 614898 174970 615134
rect 175206 614898 175248 615134
rect 174928 614866 175248 614898
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 159568 597454 159888 597486
rect 159568 597218 159610 597454
rect 159846 597218 159888 597454
rect 159568 597134 159888 597218
rect 159568 596898 159610 597134
rect 159846 596898 159888 597134
rect 159568 596866 159888 596898
rect 190288 597454 190608 597486
rect 190288 597218 190330 597454
rect 190566 597218 190608 597454
rect 190288 597134 190608 597218
rect 190288 596898 190330 597134
rect 190566 596898 190608 597134
rect 190288 596866 190608 596898
rect 144208 579454 144528 579486
rect 144208 579218 144250 579454
rect 144486 579218 144528 579454
rect 144208 579134 144528 579218
rect 144208 578898 144250 579134
rect 144486 578898 144528 579134
rect 144208 578866 144528 578898
rect 174928 579454 175248 579486
rect 174928 579218 174970 579454
rect 175206 579218 175248 579454
rect 174928 579134 175248 579218
rect 174928 578898 174970 579134
rect 175206 578898 175248 579134
rect 174928 578866 175248 578898
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 549954 135854 568338
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 135234 549718 135266 549954
rect 135502 549718 135586 549954
rect 135822 549718 135854 549954
rect 135234 549634 135854 549718
rect 135234 549398 135266 549634
rect 135502 549398 135586 549634
rect 135822 549398 135854 549634
rect 135234 542000 135854 549398
rect 138954 553674 139574 558000
rect 138954 553438 138986 553674
rect 139222 553438 139306 553674
rect 139542 553438 139574 553674
rect 138954 553354 139574 553438
rect 138954 553118 138986 553354
rect 139222 553118 139306 553354
rect 139542 553118 139574 553354
rect 138954 542000 139574 553118
rect 145794 543454 146414 558000
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 542000 146414 542898
rect 149514 547174 150134 558000
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 542000 150134 546618
rect 153234 550894 153854 558000
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 542000 153854 550338
rect 156954 554614 157574 558000
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 542000 157574 554058
rect 163794 544394 164414 558000
rect 163794 544158 163826 544394
rect 164062 544158 164146 544394
rect 164382 544158 164414 544394
rect 163794 544074 164414 544158
rect 163794 543838 163826 544074
rect 164062 543838 164146 544074
rect 164382 543838 164414 544074
rect 163794 542000 164414 543838
rect 167514 548114 168134 558000
rect 167514 547878 167546 548114
rect 167782 547878 167866 548114
rect 168102 547878 168134 548114
rect 167514 547794 168134 547878
rect 167514 547558 167546 547794
rect 167782 547558 167866 547794
rect 168102 547558 168134 547794
rect 167514 542000 168134 547558
rect 171234 549954 171854 558000
rect 171234 549718 171266 549954
rect 171502 549718 171586 549954
rect 171822 549718 171854 549954
rect 171234 549634 171854 549718
rect 171234 549398 171266 549634
rect 171502 549398 171586 549634
rect 171822 549398 171854 549634
rect 171234 542000 171854 549398
rect 174954 553674 175574 558000
rect 174954 553438 174986 553674
rect 175222 553438 175306 553674
rect 175542 553438 175574 553674
rect 174954 553354 175574 553438
rect 174954 553118 174986 553354
rect 175222 553118 175306 553354
rect 175542 553118 175574 553354
rect 174954 542000 175574 553118
rect 181794 543454 182414 558000
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 542000 182414 542898
rect 185514 547174 186134 558000
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 542000 186134 546618
rect 189234 550894 189854 558000
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 542000 189854 550338
rect 192954 554614 193574 558000
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 542000 193574 554058
rect 199794 544394 200414 558000
rect 199794 544158 199826 544394
rect 200062 544158 200146 544394
rect 200382 544158 200414 544394
rect 199794 544074 200414 544158
rect 199794 543838 199826 544074
rect 200062 543838 200146 544074
rect 200382 543838 200414 544074
rect 199794 542000 200414 543838
rect 203514 548114 204134 564618
rect 203514 547878 203546 548114
rect 203782 547878 203866 548114
rect 204102 547878 204134 548114
rect 203514 547794 204134 547878
rect 203514 547558 203546 547794
rect 203782 547558 203866 547794
rect 204102 547558 204134 547794
rect 203514 542000 204134 547558
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 549954 207854 568338
rect 207234 549718 207266 549954
rect 207502 549718 207586 549954
rect 207822 549718 207854 549954
rect 207234 549634 207854 549718
rect 207234 549398 207266 549634
rect 207502 549398 207586 549634
rect 207822 549398 207854 549634
rect 207234 542000 207854 549398
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 625099 218414 650898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 625099 222134 654618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 625099 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 625099 229574 626058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 625099 236414 632898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 625099 240134 636618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 625099 243854 640338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 625099 247574 644058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 625099 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 625099 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 625099 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 625099 265574 626058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 625099 272414 632898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 625099 276134 636618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 625099 279854 640338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 625099 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 224208 615454 224528 615486
rect 224208 615218 224250 615454
rect 224486 615218 224528 615454
rect 224208 615134 224528 615218
rect 224208 614898 224250 615134
rect 224486 614898 224528 615134
rect 224208 614866 224528 614898
rect 254928 615454 255248 615486
rect 254928 615218 254970 615454
rect 255206 615218 255248 615454
rect 254928 615134 255248 615218
rect 254928 614898 254970 615134
rect 255206 614898 255248 615134
rect 254928 614866 255248 614898
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 239568 597454 239888 597486
rect 239568 597218 239610 597454
rect 239846 597218 239888 597454
rect 239568 597134 239888 597218
rect 239568 596898 239610 597134
rect 239846 596898 239888 597134
rect 239568 596866 239888 596898
rect 270288 597454 270608 597486
rect 270288 597218 270330 597454
rect 270566 597218 270608 597454
rect 270288 597134 270608 597218
rect 270288 596898 270330 597134
rect 270566 596898 270608 597134
rect 270288 596866 270608 596898
rect 224208 579454 224528 579486
rect 224208 579218 224250 579454
rect 224486 579218 224528 579454
rect 224208 579134 224528 579218
rect 224208 578898 224250 579134
rect 224486 578898 224528 579134
rect 224208 578866 224528 578898
rect 254928 579454 255248 579486
rect 254928 579218 254970 579454
rect 255206 579218 255248 579454
rect 254928 579134 255248 579218
rect 254928 578898 254970 579134
rect 255206 578898 255248 579134
rect 254928 578866 255248 578898
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 553674 211574 572058
rect 210954 553438 210986 553674
rect 211222 553438 211306 553674
rect 211542 553438 211574 553674
rect 210954 553354 211574 553438
rect 210954 553118 210986 553354
rect 211222 553118 211306 553354
rect 211542 553118 211574 553354
rect 210954 542000 211574 553118
rect 217794 543454 218414 558000
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 542000 218414 542898
rect 221514 547174 222134 558000
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 542000 222134 546618
rect 225234 550894 225854 558000
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 542000 225854 550338
rect 228954 554614 229574 558000
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 542000 229574 554058
rect 235794 544394 236414 558000
rect 235794 544158 235826 544394
rect 236062 544158 236146 544394
rect 236382 544158 236414 544394
rect 235794 544074 236414 544158
rect 235794 543838 235826 544074
rect 236062 543838 236146 544074
rect 236382 543838 236414 544074
rect 235794 542000 236414 543838
rect 239514 548114 240134 558000
rect 239514 547878 239546 548114
rect 239782 547878 239866 548114
rect 240102 547878 240134 548114
rect 239514 547794 240134 547878
rect 239514 547558 239546 547794
rect 239782 547558 239866 547794
rect 240102 547558 240134 547794
rect 239514 542000 240134 547558
rect 243234 549954 243854 558000
rect 243234 549718 243266 549954
rect 243502 549718 243586 549954
rect 243822 549718 243854 549954
rect 243234 549634 243854 549718
rect 243234 549398 243266 549634
rect 243502 549398 243586 549634
rect 243822 549398 243854 549634
rect 243234 542000 243854 549398
rect 246954 553674 247574 558000
rect 246954 553438 246986 553674
rect 247222 553438 247306 553674
rect 247542 553438 247574 553674
rect 246954 553354 247574 553438
rect 246954 553118 246986 553354
rect 247222 553118 247306 553354
rect 247542 553118 247574 553354
rect 246954 542000 247574 553118
rect 253794 543454 254414 558000
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 542000 254414 542898
rect 257514 547174 258134 558000
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 542000 258134 546618
rect 261234 550894 261854 558000
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 542000 261854 550338
rect 264954 554614 265574 558000
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 542000 265574 554058
rect 271794 544394 272414 558000
rect 271794 544158 271826 544394
rect 272062 544158 272146 544394
rect 272382 544158 272414 544394
rect 271794 544074 272414 544158
rect 271794 543838 271826 544074
rect 272062 543838 272146 544074
rect 272382 543838 272414 544074
rect 271794 542000 272414 543838
rect 275514 548114 276134 558000
rect 275514 547878 275546 548114
rect 275782 547878 275866 548114
rect 276102 547878 276134 548114
rect 275514 547794 276134 547878
rect 275514 547558 275546 547794
rect 275782 547558 275866 547794
rect 276102 547558 276134 547794
rect 275514 542000 276134 547558
rect 279234 549954 279854 558000
rect 279234 549718 279266 549954
rect 279502 549718 279586 549954
rect 279822 549718 279854 549954
rect 279234 549634 279854 549718
rect 279234 549398 279266 549634
rect 279502 549398 279586 549634
rect 279822 549398 279854 549634
rect 279234 542000 279854 549398
rect 282954 553674 283574 558000
rect 282954 553438 282986 553674
rect 283222 553438 283306 553674
rect 283542 553438 283574 553674
rect 282954 553354 283574 553438
rect 282954 553118 282986 553354
rect 283222 553118 283306 553354
rect 283542 553118 283574 553354
rect 282954 542000 283574 553118
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 542000 290414 542898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 542000 294134 546618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 542000 297854 550338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300163 543148 300229 543149
rect 300163 543084 300164 543148
rect 300228 543084 300229 543148
rect 300163 543083 300229 543084
rect 299979 542740 300045 542741
rect 299979 542676 299980 542740
rect 300044 542676 300045 542740
rect 299979 542675 300045 542676
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 79568 525454 79888 525486
rect 79568 525218 79610 525454
rect 79846 525218 79888 525454
rect 79568 525134 79888 525218
rect 79568 524898 79610 525134
rect 79846 524898 79888 525134
rect 79568 524866 79888 524898
rect 110288 525454 110608 525486
rect 110288 525218 110330 525454
rect 110566 525218 110608 525454
rect 110288 525134 110608 525218
rect 110288 524898 110330 525134
rect 110566 524898 110608 525134
rect 110288 524866 110608 524898
rect 141008 525454 141328 525486
rect 141008 525218 141050 525454
rect 141286 525218 141328 525454
rect 141008 525134 141328 525218
rect 141008 524898 141050 525134
rect 141286 524898 141328 525134
rect 141008 524866 141328 524898
rect 171728 525454 172048 525486
rect 171728 525218 171770 525454
rect 172006 525218 172048 525454
rect 171728 525134 172048 525218
rect 171728 524898 171770 525134
rect 172006 524898 172048 525134
rect 171728 524866 172048 524898
rect 202448 525454 202768 525486
rect 202448 525218 202490 525454
rect 202726 525218 202768 525454
rect 202448 525134 202768 525218
rect 202448 524898 202490 525134
rect 202726 524898 202768 525134
rect 202448 524866 202768 524898
rect 233168 525454 233488 525486
rect 233168 525218 233210 525454
rect 233446 525218 233488 525454
rect 233168 525134 233488 525218
rect 233168 524898 233210 525134
rect 233446 524898 233488 525134
rect 233168 524866 233488 524898
rect 263888 525454 264208 525486
rect 263888 525218 263930 525454
rect 264166 525218 264208 525454
rect 263888 525134 264208 525218
rect 263888 524898 263930 525134
rect 264166 524898 264208 525134
rect 263888 524866 264208 524898
rect 294608 525454 294928 525486
rect 294608 525218 294650 525454
rect 294886 525218 294928 525454
rect 294608 525134 294928 525218
rect 294608 524898 294650 525134
rect 294886 524898 294928 525134
rect 294608 524866 294928 524898
rect 299982 517309 300042 542675
rect 300166 520165 300226 543083
rect 300954 542000 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 300163 520164 300229 520165
rect 300163 520100 300164 520164
rect 300228 520100 300229 520164
rect 300163 520099 300229 520100
rect 299979 517308 300045 517309
rect 299979 517244 299980 517308
rect 300044 517244 300045 517308
rect 299979 517243 300045 517244
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 54707 478004 54773 478005
rect 54707 477940 54708 478004
rect 54772 477940 54773 478004
rect 54707 477939 54773 477940
rect 54339 305012 54405 305013
rect 54339 304948 54340 305012
rect 54404 304948 54405 305012
rect 54339 304947 54405 304948
rect 54710 162757 54770 477939
rect 55443 465764 55509 465765
rect 55443 465700 55444 465764
rect 55508 465700 55509 465764
rect 55443 465699 55509 465700
rect 55075 460868 55141 460869
rect 55075 460804 55076 460868
rect 55140 460804 55141 460868
rect 55075 460803 55141 460804
rect 54891 460732 54957 460733
rect 54891 460668 54892 460732
rect 54956 460668 54957 460732
rect 54891 460667 54957 460668
rect 54707 162756 54773 162757
rect 54707 162692 54708 162756
rect 54772 162692 54773 162756
rect 54707 162691 54773 162692
rect 54894 59125 54954 460667
rect 54891 59124 54957 59125
rect 54891 59060 54892 59124
rect 54956 59060 54957 59124
rect 54891 59059 54957 59060
rect 55078 56677 55138 460803
rect 55446 164389 55506 465699
rect 55627 459644 55693 459645
rect 55627 459580 55628 459644
rect 55692 459580 55693 459644
rect 55627 459579 55693 459580
rect 55443 164388 55509 164389
rect 55443 164324 55444 164388
rect 55508 164324 55509 164388
rect 55443 164323 55509 164324
rect 55075 56676 55141 56677
rect 55075 56612 55076 56676
rect 55140 56612 55141 56676
rect 55075 56611 55141 56612
rect 53603 56540 53669 56541
rect 53603 56476 53604 56540
rect 53668 56476 53669 56540
rect 53603 56475 53669 56476
rect 55630 56269 55690 459579
rect 55794 453454 56414 488898
rect 79568 489454 79888 489486
rect 79568 489218 79610 489454
rect 79846 489218 79888 489454
rect 79568 489134 79888 489218
rect 79568 488898 79610 489134
rect 79846 488898 79888 489134
rect 79568 488866 79888 488898
rect 110288 489454 110608 489486
rect 110288 489218 110330 489454
rect 110566 489218 110608 489454
rect 110288 489134 110608 489218
rect 110288 488898 110330 489134
rect 110566 488898 110608 489134
rect 110288 488866 110608 488898
rect 141008 489454 141328 489486
rect 141008 489218 141050 489454
rect 141286 489218 141328 489454
rect 141008 489134 141328 489218
rect 141008 488898 141050 489134
rect 141286 488898 141328 489134
rect 141008 488866 141328 488898
rect 171728 489454 172048 489486
rect 171728 489218 171770 489454
rect 172006 489218 172048 489454
rect 171728 489134 172048 489218
rect 171728 488898 171770 489134
rect 172006 488898 172048 489134
rect 171728 488866 172048 488898
rect 202448 489454 202768 489486
rect 202448 489218 202490 489454
rect 202726 489218 202768 489454
rect 202448 489134 202768 489218
rect 202448 488898 202490 489134
rect 202726 488898 202768 489134
rect 202448 488866 202768 488898
rect 233168 489454 233488 489486
rect 233168 489218 233210 489454
rect 233446 489218 233488 489454
rect 233168 489134 233488 489218
rect 233168 488898 233210 489134
rect 233446 488898 233488 489134
rect 233168 488866 233488 488898
rect 263888 489454 264208 489486
rect 263888 489218 263930 489454
rect 264166 489218 264208 489454
rect 263888 489134 264208 489218
rect 263888 488898 263930 489134
rect 264166 488898 264208 489134
rect 263888 488866 264208 488898
rect 294608 489454 294928 489486
rect 294608 489218 294650 489454
rect 294886 489218 294928 489454
rect 294608 489134 294928 489218
rect 294608 488898 294650 489134
rect 294886 488898 294928 489134
rect 294608 488866 294928 488898
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 59307 478820 59373 478821
rect 59307 478756 59308 478820
rect 59372 478756 59373 478820
rect 59307 478755 59373 478756
rect 202459 478820 202525 478821
rect 202459 478756 202460 478820
rect 202524 478756 202525 478820
rect 202459 478755 202525 478756
rect 57651 478276 57717 478277
rect 57651 478212 57652 478276
rect 57716 478212 57717 478276
rect 57651 478211 57717 478212
rect 57283 475828 57349 475829
rect 57283 475764 57284 475828
rect 57348 475764 57349 475828
rect 57283 475763 57349 475764
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 57286 372741 57346 475763
rect 57467 383620 57533 383621
rect 57467 383556 57468 383620
rect 57532 383556 57533 383620
rect 57467 383555 57533 383556
rect 57283 372740 57349 372741
rect 57283 372676 57284 372740
rect 57348 372676 57349 372740
rect 57283 372675 57349 372676
rect 57099 371380 57165 371381
rect 57099 371316 57100 371380
rect 57164 371316 57165 371380
rect 57099 371315 57165 371316
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 57102 276181 57162 371315
rect 57099 276180 57165 276181
rect 57099 276116 57100 276180
rect 57164 276116 57165 276180
rect 57099 276115 57165 276116
rect 57283 276044 57349 276045
rect 57283 275980 57284 276044
rect 57348 275980 57349 276044
rect 57283 275979 57349 275980
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57286 269109 57346 275979
rect 57283 269108 57349 269109
rect 57283 269044 57284 269108
rect 57348 269044 57349 269108
rect 57283 269043 57349 269044
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 57470 173093 57530 383555
rect 57467 173092 57533 173093
rect 57467 173028 57468 173092
rect 57532 173028 57533 173092
rect 57467 173027 57533 173028
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57654 164117 57714 478211
rect 58571 461548 58637 461549
rect 58571 461484 58572 461548
rect 58636 461484 58637 461548
rect 58571 461483 58637 461484
rect 57835 458828 57901 458829
rect 57835 458764 57836 458828
rect 57900 458764 57901 458828
rect 57835 458763 57901 458764
rect 57651 164116 57717 164117
rect 57651 164052 57652 164116
rect 57716 164052 57717 164116
rect 57651 164051 57717 164052
rect 57651 160172 57717 160173
rect 57651 160108 57652 160172
rect 57716 160108 57717 160172
rect 57651 160107 57717 160108
rect 57467 146028 57533 146029
rect 57467 145964 57468 146028
rect 57532 145964 57533 146028
rect 57467 145963 57533 145964
rect 57470 144805 57530 145963
rect 57099 144804 57165 144805
rect 57099 144740 57100 144804
rect 57164 144740 57165 144804
rect 57099 144739 57165 144740
rect 57467 144804 57533 144805
rect 57467 144740 57468 144804
rect 57532 144740 57533 144804
rect 57467 144739 57533 144740
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 57102 57357 57162 144739
rect 57467 140860 57533 140861
rect 57467 140796 57468 140860
rect 57532 140796 57533 140860
rect 57467 140795 57533 140796
rect 57099 57356 57165 57357
rect 57099 57292 57100 57356
rect 57164 57292 57165 57356
rect 57099 57291 57165 57292
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55627 56268 55693 56269
rect 55627 56204 55628 56268
rect 55692 56204 55693 56268
rect 55627 56203 55693 56204
rect 50843 54908 50909 54909
rect 50843 54844 50844 54908
rect 50908 54844 50909 54908
rect 50843 54843 50909 54844
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 56898
rect 57470 54773 57530 140795
rect 57654 57765 57714 160107
rect 57838 70413 57898 458763
rect 58574 175269 58634 461483
rect 59123 460052 59189 460053
rect 59123 459988 59124 460052
rect 59188 459988 59189 460052
rect 59123 459987 59189 459988
rect 58939 459100 59005 459101
rect 58939 459036 58940 459100
rect 59004 459036 59005 459100
rect 58939 459035 59005 459036
rect 58755 458964 58821 458965
rect 58755 458900 58756 458964
rect 58820 458900 58821 458964
rect 58755 458899 58821 458900
rect 58571 175268 58637 175269
rect 58571 175204 58572 175268
rect 58636 175204 58637 175268
rect 58571 175203 58637 175204
rect 57835 70412 57901 70413
rect 57835 70348 57836 70412
rect 57900 70348 57901 70412
rect 57835 70347 57901 70348
rect 57651 57764 57717 57765
rect 57651 57700 57652 57764
rect 57716 57700 57717 57764
rect 57651 57699 57717 57700
rect 58758 57493 58818 458899
rect 58755 57492 58821 57493
rect 58755 57428 58756 57492
rect 58820 57428 58821 57492
rect 58755 57427 58821 57428
rect 58942 57085 59002 459035
rect 59126 57221 59186 459987
rect 59310 58445 59370 478755
rect 198043 478684 198109 478685
rect 198043 478620 198044 478684
rect 198108 478620 198109 478684
rect 198043 478619 198109 478620
rect 196571 478548 196637 478549
rect 196571 478484 196572 478548
rect 196636 478484 196637 478548
rect 196571 478483 196637 478484
rect 59514 474234 60134 478000
rect 59514 473998 59546 474234
rect 59782 473998 59866 474234
rect 60102 473998 60134 474234
rect 59514 473914 60134 473998
rect 59514 473678 59546 473914
rect 59782 473678 59866 473914
rect 60102 473678 60134 473914
rect 59514 460308 60134 473678
rect 63234 470078 63854 478000
rect 63234 469842 63266 470078
rect 63502 469842 63586 470078
rect 63822 469842 63854 470078
rect 63234 469758 63854 469842
rect 63234 469522 63266 469758
rect 63502 469522 63586 469758
rect 63822 469522 63854 469758
rect 63234 460308 63854 469522
rect 66954 464614 67574 478000
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 460308 67574 464058
rect 73794 471454 74414 478000
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 460308 74414 470898
rect 77514 475174 78134 478000
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 460308 78134 474618
rect 81234 469138 81854 478000
rect 81234 468902 81266 469138
rect 81502 468902 81586 469138
rect 81822 468902 81854 469138
rect 81234 468818 81854 468902
rect 81234 468582 81266 468818
rect 81502 468582 81586 468818
rect 81822 468582 81854 468818
rect 81234 460308 81854 468582
rect 84954 465554 85574 478000
rect 84954 465318 84986 465554
rect 85222 465318 85306 465554
rect 85542 465318 85574 465554
rect 84954 465234 85574 465318
rect 84954 464998 84986 465234
rect 85222 464998 85306 465234
rect 85542 464998 85574 465234
rect 84954 460308 85574 464998
rect 91794 470514 92414 478000
rect 91794 470278 91826 470514
rect 92062 470278 92146 470514
rect 92382 470278 92414 470514
rect 91794 470194 92414 470278
rect 91794 469958 91826 470194
rect 92062 469958 92146 470194
rect 92382 469958 92414 470194
rect 91794 460308 92414 469958
rect 95514 474234 96134 478000
rect 95514 473998 95546 474234
rect 95782 473998 95866 474234
rect 96102 473998 96134 474234
rect 95514 473914 96134 473998
rect 95514 473678 95546 473914
rect 95782 473678 95866 473914
rect 96102 473678 96134 473914
rect 95514 460308 96134 473678
rect 99234 470078 99854 478000
rect 99234 469842 99266 470078
rect 99502 469842 99586 470078
rect 99822 469842 99854 470078
rect 99234 469758 99854 469842
rect 99234 469522 99266 469758
rect 99502 469522 99586 469758
rect 99822 469522 99854 469758
rect 99234 460308 99854 469522
rect 102954 464614 103574 478000
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 460308 103574 464058
rect 109794 471454 110414 478000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 460308 110414 470898
rect 113514 475174 114134 478000
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 460308 114134 474618
rect 117234 469138 117854 478000
rect 117234 468902 117266 469138
rect 117502 468902 117586 469138
rect 117822 468902 117854 469138
rect 117234 468818 117854 468902
rect 117234 468582 117266 468818
rect 117502 468582 117586 468818
rect 117822 468582 117854 468818
rect 117234 460308 117854 468582
rect 120954 465554 121574 478000
rect 120954 465318 120986 465554
rect 121222 465318 121306 465554
rect 121542 465318 121574 465554
rect 120954 465234 121574 465318
rect 120954 464998 120986 465234
rect 121222 464998 121306 465234
rect 121542 464998 121574 465234
rect 120954 460308 121574 464998
rect 127794 470514 128414 478000
rect 127794 470278 127826 470514
rect 128062 470278 128146 470514
rect 128382 470278 128414 470514
rect 127794 470194 128414 470278
rect 127794 469958 127826 470194
rect 128062 469958 128146 470194
rect 128382 469958 128414 470194
rect 127794 460308 128414 469958
rect 131514 474234 132134 478000
rect 131514 473998 131546 474234
rect 131782 473998 131866 474234
rect 132102 473998 132134 474234
rect 131514 473914 132134 473998
rect 131514 473678 131546 473914
rect 131782 473678 131866 473914
rect 132102 473678 132134 473914
rect 131514 460308 132134 473678
rect 135234 470078 135854 478000
rect 135234 469842 135266 470078
rect 135502 469842 135586 470078
rect 135822 469842 135854 470078
rect 135234 469758 135854 469842
rect 135234 469522 135266 469758
rect 135502 469522 135586 469758
rect 135822 469522 135854 469758
rect 135234 460308 135854 469522
rect 138954 464614 139574 478000
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 460308 139574 464058
rect 145794 471454 146414 478000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 460308 146414 470898
rect 149514 475174 150134 478000
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 460308 150134 474618
rect 153234 469138 153854 478000
rect 153234 468902 153266 469138
rect 153502 468902 153586 469138
rect 153822 468902 153854 469138
rect 153234 468818 153854 468902
rect 153234 468582 153266 468818
rect 153502 468582 153586 468818
rect 153822 468582 153854 468818
rect 153234 460308 153854 468582
rect 156954 465554 157574 478000
rect 156954 465318 156986 465554
rect 157222 465318 157306 465554
rect 157542 465318 157574 465554
rect 156954 465234 157574 465318
rect 156954 464998 156986 465234
rect 157222 464998 157306 465234
rect 157542 464998 157574 465234
rect 156954 460308 157574 464998
rect 163794 470514 164414 478000
rect 163794 470278 163826 470514
rect 164062 470278 164146 470514
rect 164382 470278 164414 470514
rect 163794 470194 164414 470278
rect 163794 469958 163826 470194
rect 164062 469958 164146 470194
rect 164382 469958 164414 470194
rect 163794 460308 164414 469958
rect 167514 474234 168134 478000
rect 167514 473998 167546 474234
rect 167782 473998 167866 474234
rect 168102 473998 168134 474234
rect 167514 473914 168134 473998
rect 167514 473678 167546 473914
rect 167782 473678 167866 473914
rect 168102 473678 168134 473914
rect 167514 460308 168134 473678
rect 171234 470078 171854 478000
rect 171234 469842 171266 470078
rect 171502 469842 171586 470078
rect 171822 469842 171854 470078
rect 171234 469758 171854 469842
rect 171234 469522 171266 469758
rect 171502 469522 171586 469758
rect 171822 469522 171854 469758
rect 171234 460308 171854 469522
rect 174954 464614 175574 478000
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 460308 175574 464058
rect 181794 471454 182414 478000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 179643 461684 179709 461685
rect 179643 461620 179644 461684
rect 179708 461620 179709 461684
rect 179643 461619 179709 461620
rect 178355 461412 178421 461413
rect 178355 461348 178356 461412
rect 178420 461348 178421 461412
rect 178355 461347 178421 461348
rect 178358 458690 178418 461347
rect 179646 458690 179706 461619
rect 181794 460308 182414 470898
rect 185514 475174 186134 478000
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 460308 186134 474618
rect 189234 469138 189854 478000
rect 189234 468902 189266 469138
rect 189502 468902 189586 469138
rect 189822 468902 189854 469138
rect 189234 468818 189854 468902
rect 189234 468582 189266 468818
rect 189502 468582 189586 468818
rect 189822 468582 189854 468818
rect 189234 460308 189854 468582
rect 192954 465554 193574 478000
rect 192954 465318 192986 465554
rect 193222 465318 193306 465554
rect 193542 465318 193574 465554
rect 192954 465234 193574 465318
rect 192954 464998 192986 465234
rect 193222 464998 193306 465234
rect 193542 464998 193574 465234
rect 190867 461004 190933 461005
rect 190867 460940 190868 461004
rect 190932 460940 190933 461004
rect 190867 460939 190933 460940
rect 190870 458690 190930 460939
rect 192954 460308 193574 464998
rect 178358 458630 178524 458690
rect 179646 458630 179748 458690
rect 178464 458202 178524 458630
rect 179688 458202 179748 458630
rect 190840 458630 190930 458690
rect 190840 458202 190900 458630
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 60952 399454 61300 399486
rect 60952 399218 61008 399454
rect 61244 399218 61300 399454
rect 60952 399134 61300 399218
rect 60952 398898 61008 399134
rect 61244 398898 61300 399134
rect 60952 398866 61300 398898
rect 195320 399454 195668 399486
rect 195320 399218 195376 399454
rect 195612 399218 195668 399454
rect 195320 399134 195668 399218
rect 195320 398898 195376 399134
rect 195612 398898 195668 399134
rect 195320 398866 195668 398898
rect 60272 381454 60620 381486
rect 60272 381218 60328 381454
rect 60564 381218 60620 381454
rect 60272 381134 60620 381218
rect 60272 380898 60328 381134
rect 60564 380898 60620 381134
rect 60272 380866 60620 380898
rect 196000 381454 196348 381486
rect 196000 381218 196056 381454
rect 196292 381218 196348 381454
rect 196000 381134 196348 381218
rect 196000 380898 196056 381134
rect 196292 380898 196348 381134
rect 196000 380866 196348 380898
rect 76086 374990 76666 375050
rect 59514 366234 60134 373000
rect 59514 365998 59546 366234
rect 59782 365998 59866 366234
rect 60102 365998 60134 366234
rect 59514 365914 60134 365998
rect 59514 365678 59546 365914
rect 59782 365678 59866 365914
rect 60102 365678 60134 365914
rect 59514 355308 60134 365678
rect 63234 369954 63854 373000
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 63854 369954
rect 63234 369634 63854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 63854 369634
rect 63234 355308 63854 369398
rect 66954 356614 67574 373000
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 355308 67574 356058
rect 73794 363454 74414 373000
rect 76606 371925 76666 374990
rect 77158 372605 77218 375050
rect 78262 374990 78506 375050
rect 79622 374990 79978 375050
rect 77155 372604 77221 372605
rect 77155 372540 77156 372604
rect 77220 372540 77221 372604
rect 77155 372539 77221 372540
rect 76603 371924 76669 371925
rect 76603 371860 76604 371924
rect 76668 371860 76669 371924
rect 76603 371859 76669 371860
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 355308 74414 362898
rect 77514 367174 78134 373000
rect 78446 372469 78506 374990
rect 79918 372469 79978 374990
rect 80470 374990 80574 375050
rect 81798 374990 82002 375050
rect 83158 374990 83842 375050
rect 84246 374990 84578 375050
rect 80470 372469 80530 374990
rect 78443 372468 78509 372469
rect 78443 372404 78444 372468
rect 78508 372404 78509 372468
rect 78443 372403 78509 372404
rect 79915 372468 79981 372469
rect 79915 372404 79916 372468
rect 79980 372404 79981 372468
rect 79915 372403 79981 372404
rect 80467 372468 80533 372469
rect 80467 372404 80468 372468
rect 80532 372404 80533 372468
rect 80467 372403 80533 372404
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 355308 78134 366618
rect 81234 370894 81854 373000
rect 81942 372605 82002 374990
rect 83782 373829 83842 374990
rect 83779 373828 83845 373829
rect 83779 373764 83780 373828
rect 83844 373764 83845 373828
rect 83779 373763 83845 373764
rect 81939 372604 82005 372605
rect 81939 372540 81940 372604
rect 82004 372540 82005 372604
rect 81939 372539 82005 372540
rect 84518 372469 84578 374990
rect 84702 374990 85470 375050
rect 86558 374990 86786 375050
rect 87646 374990 88074 375050
rect 88326 374990 88442 375050
rect 88734 374990 89362 375050
rect 84702 372605 84762 374990
rect 84699 372604 84765 372605
rect 84699 372540 84700 372604
rect 84764 372540 84765 372604
rect 84699 372539 84765 372540
rect 84515 372468 84581 372469
rect 84515 372404 84516 372468
rect 84580 372404 84581 372468
rect 84515 372403 84581 372404
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 355308 81854 370338
rect 84954 357554 85574 373000
rect 86726 372605 86786 374990
rect 88014 372605 88074 374990
rect 88382 373421 88442 374990
rect 88379 373420 88445 373421
rect 88379 373356 88380 373420
rect 88444 373356 88445 373420
rect 88379 373355 88445 373356
rect 89302 372605 89362 374990
rect 90038 372605 90098 375050
rect 90222 374990 90774 375050
rect 91318 374990 91570 375050
rect 92406 374990 92490 375050
rect 90222 373149 90282 374990
rect 90219 373148 90285 373149
rect 90219 373084 90220 373148
rect 90284 373084 90285 373148
rect 90219 373083 90285 373084
rect 91510 372605 91570 374990
rect 92430 373149 92490 374990
rect 93350 374990 93494 375050
rect 92427 373148 92493 373149
rect 92427 373084 92428 373148
rect 92492 373084 92493 373148
rect 92427 373083 92493 373084
rect 86723 372604 86789 372605
rect 86723 372540 86724 372604
rect 86788 372540 86789 372604
rect 86723 372539 86789 372540
rect 88011 372604 88077 372605
rect 88011 372540 88012 372604
rect 88076 372540 88077 372604
rect 88011 372539 88077 372540
rect 89299 372604 89365 372605
rect 89299 372540 89300 372604
rect 89364 372540 89365 372604
rect 89299 372539 89365 372540
rect 90035 372604 90101 372605
rect 90035 372540 90036 372604
rect 90100 372540 90101 372604
rect 90035 372539 90101 372540
rect 91507 372604 91573 372605
rect 91507 372540 91508 372604
rect 91572 372540 91573 372604
rect 91507 372539 91573 372540
rect 84954 357318 84986 357554
rect 85222 357318 85306 357554
rect 85542 357318 85574 357554
rect 84954 357234 85574 357318
rect 84954 356998 84986 357234
rect 85222 356998 85306 357234
rect 85542 356998 85574 357234
rect 84954 355308 85574 356998
rect 91794 364394 92414 373000
rect 93350 372605 93410 374990
rect 93600 374509 93660 375020
rect 94582 374990 95250 375050
rect 93597 374508 93663 374509
rect 93597 374444 93598 374508
rect 93662 374444 93663 374508
rect 93597 374443 93663 374444
rect 95190 373149 95250 374990
rect 95374 374990 95942 375050
rect 96078 374990 96170 375050
rect 97030 374990 97642 375050
rect 98118 374990 98194 375050
rect 95187 373148 95253 373149
rect 95187 373084 95188 373148
rect 95252 373084 95253 373148
rect 95187 373083 95253 373084
rect 93347 372604 93413 372605
rect 93347 372540 93348 372604
rect 93412 372540 93413 372604
rect 93347 372539 93413 372540
rect 95187 371652 95253 371653
rect 95187 371588 95188 371652
rect 95252 371650 95253 371652
rect 95374 371650 95434 374990
rect 96110 373421 96170 374990
rect 96107 373420 96173 373421
rect 96107 373356 96108 373420
rect 96172 373356 96173 373420
rect 96107 373355 96173 373356
rect 95252 371590 95434 371650
rect 95252 371588 95253 371590
rect 95187 371587 95253 371588
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 92414 364394
rect 91794 364074 92414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 92414 364074
rect 91794 355308 92414 363838
rect 95514 366234 96134 373000
rect 97582 371517 97642 374990
rect 98134 371653 98194 374990
rect 98318 374990 98526 375050
rect 99478 374990 100034 375050
rect 100702 374990 100770 375050
rect 98318 373421 98378 374990
rect 98315 373420 98381 373421
rect 98315 373356 98316 373420
rect 98380 373356 98381 373420
rect 98315 373355 98381 373356
rect 98131 371652 98197 371653
rect 98131 371588 98132 371652
rect 98196 371588 98197 371652
rect 98131 371587 98197 371588
rect 97579 371516 97645 371517
rect 97579 371452 97580 371516
rect 97644 371452 97645 371516
rect 97579 371451 97645 371452
rect 95514 365998 95546 366234
rect 95782 365998 95866 366234
rect 96102 365998 96134 366234
rect 95514 365914 96134 365998
rect 95514 365678 95546 365914
rect 95782 365678 95866 365914
rect 96102 365678 96134 365914
rect 95514 355308 96134 365678
rect 99234 369954 99854 373000
rect 99974 371653 100034 374990
rect 99971 371652 100037 371653
rect 99971 371588 99972 371652
rect 100036 371588 100037 371652
rect 99971 371587 100037 371588
rect 100710 371517 100770 374990
rect 100894 374990 101110 375050
rect 101790 374990 102058 375050
rect 100894 373693 100954 374990
rect 100891 373692 100957 373693
rect 100891 373628 100892 373692
rect 100956 373628 100957 373692
rect 100891 373627 100957 373628
rect 101998 372605 102058 374990
rect 102734 374990 102878 375050
rect 101995 372604 102061 372605
rect 101995 372540 101996 372604
rect 102060 372540 102061 372604
rect 101995 372539 102061 372540
rect 100707 371516 100773 371517
rect 100707 371452 100708 371516
rect 100772 371452 100773 371516
rect 100707 371451 100773 371452
rect 102734 371381 102794 374990
rect 103528 374509 103588 375020
rect 103966 374990 104634 375050
rect 103525 374508 103591 374509
rect 103525 374444 103526 374508
rect 103590 374444 103591 374508
rect 103525 374443 103591 374444
rect 102731 371380 102797 371381
rect 102731 371316 102732 371380
rect 102796 371316 102797 371380
rect 102731 371315 102797 371316
rect 99234 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 99854 369954
rect 99234 369634 99854 369718
rect 99234 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 99854 369634
rect 99234 355308 99854 369398
rect 102954 356614 103574 373000
rect 104574 372197 104634 374990
rect 104571 372196 104637 372197
rect 104571 372132 104572 372196
rect 104636 372132 104637 372196
rect 104571 372131 104637 372132
rect 105310 371653 105370 375050
rect 105494 374990 106006 375050
rect 105494 373557 105554 374990
rect 105491 373556 105557 373557
rect 105491 373492 105492 373556
rect 105556 373492 105557 373556
rect 105491 373491 105557 373492
rect 105307 371652 105373 371653
rect 105307 371588 105308 371652
rect 105372 371588 105373 371652
rect 105307 371587 105373 371588
rect 106414 371109 106474 375050
rect 107518 374990 107638 375050
rect 107886 374990 108318 375050
rect 108726 374990 109050 375050
rect 107518 371381 107578 374990
rect 107886 373693 107946 374990
rect 107883 373692 107949 373693
rect 107883 373628 107884 373692
rect 107948 373628 107949 373692
rect 107883 373627 107949 373628
rect 108990 371925 109050 374990
rect 109542 374990 109814 375050
rect 110462 374990 111038 375050
rect 111174 374990 111810 375050
rect 112262 374990 112914 375050
rect 109542 372197 109602 374990
rect 110462 373557 110522 374990
rect 110459 373556 110525 373557
rect 110459 373492 110460 373556
rect 110524 373492 110525 373556
rect 110459 373491 110525 373492
rect 109539 372196 109605 372197
rect 109539 372132 109540 372196
rect 109604 372132 109605 372196
rect 109539 372131 109605 372132
rect 108987 371924 109053 371925
rect 108987 371860 108988 371924
rect 109052 371860 109053 371924
rect 108987 371859 109053 371860
rect 107515 371380 107581 371381
rect 107515 371316 107516 371380
rect 107580 371316 107581 371380
rect 107515 371315 107581 371316
rect 106411 371108 106477 371109
rect 106411 371044 106412 371108
rect 106476 371044 106477 371108
rect 106411 371043 106477 371044
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 355308 103574 356058
rect 109794 363454 110414 373000
rect 111750 371517 111810 374990
rect 112854 372605 112914 374990
rect 113222 374990 113350 375050
rect 112851 372604 112917 372605
rect 112851 372540 112852 372604
rect 112916 372540 112917 372604
rect 112851 372539 112917 372540
rect 113222 372061 113282 374990
rect 113592 374370 113652 375020
rect 114438 374990 114570 375050
rect 113590 374310 113652 374370
rect 113590 373693 113650 374310
rect 113587 373692 113653 373693
rect 113587 373628 113588 373692
rect 113652 373628 113653 373692
rect 113587 373627 113653 373628
rect 113219 372060 113285 372061
rect 113219 371996 113220 372060
rect 113284 371996 113285 372060
rect 113219 371995 113285 371996
rect 111747 371516 111813 371517
rect 111747 371452 111748 371516
rect 111812 371452 111813 371516
rect 111747 371451 111813 371452
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 355308 110414 362898
rect 113514 367174 114134 373000
rect 114510 372605 114570 374990
rect 115768 374370 115828 375020
rect 116040 374509 116100 375020
rect 117022 374990 117146 375050
rect 118110 374990 118250 375050
rect 116037 374508 116103 374509
rect 116037 374444 116038 374508
rect 116102 374444 116103 374508
rect 116037 374443 116103 374444
rect 115768 374310 115858 374370
rect 114507 372604 114573 372605
rect 114507 372540 114508 372604
rect 114572 372540 114573 372604
rect 114507 372539 114573 372540
rect 115798 371789 115858 374310
rect 115795 371788 115861 371789
rect 115795 371724 115796 371788
rect 115860 371724 115861 371788
rect 115795 371723 115861 371724
rect 117086 371381 117146 374990
rect 117083 371380 117149 371381
rect 117083 371316 117084 371380
rect 117148 371316 117149 371380
rect 117083 371315 117149 371316
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 355308 114134 366618
rect 117234 370894 117854 373000
rect 118190 372469 118250 374990
rect 118374 374990 118518 375050
rect 119198 374990 119906 375050
rect 120966 374990 121378 375050
rect 118374 373693 118434 374990
rect 118371 373692 118437 373693
rect 118371 373628 118372 373692
rect 118436 373628 118437 373692
rect 118371 373627 118437 373628
rect 119846 373557 119906 374990
rect 121318 373693 121378 374990
rect 122974 374990 123550 375050
rect 125734 374990 125998 375050
rect 128310 374990 128922 375050
rect 131030 374990 131130 375050
rect 133478 374990 133706 375050
rect 135926 374990 136466 375050
rect 138510 374990 139226 375050
rect 140958 374990 141618 375050
rect 121315 373692 121381 373693
rect 121315 373628 121316 373692
rect 121380 373628 121381 373692
rect 121315 373627 121381 373628
rect 119843 373556 119909 373557
rect 119843 373492 119844 373556
rect 119908 373492 119909 373556
rect 119843 373491 119909 373492
rect 122974 373421 123034 374990
rect 125734 373693 125794 374990
rect 128862 373693 128922 374990
rect 131070 373693 131130 374990
rect 133646 373693 133706 374990
rect 136406 373693 136466 374990
rect 139166 373693 139226 374990
rect 141558 373693 141618 374990
rect 143512 374509 143572 375020
rect 145990 374990 146218 375050
rect 148574 374990 148978 375050
rect 151022 374990 151738 375050
rect 146158 374509 146218 374990
rect 143509 374508 143575 374509
rect 143509 374444 143510 374508
rect 143574 374444 143575 374508
rect 143509 374443 143575 374444
rect 146155 374508 146221 374509
rect 146155 374444 146156 374508
rect 146220 374444 146221 374508
rect 146155 374443 146221 374444
rect 148918 374237 148978 374990
rect 148915 374236 148981 374237
rect 148915 374172 148916 374236
rect 148980 374172 148981 374236
rect 148915 374171 148981 374172
rect 151678 373693 151738 374990
rect 153440 374509 153500 375020
rect 155918 374990 156522 375050
rect 156462 374509 156522 374990
rect 158486 374509 158546 375050
rect 160920 374509 160980 375020
rect 163368 374645 163428 375020
rect 165952 374645 166012 375020
rect 182958 374990 183254 375050
rect 163365 374644 163431 374645
rect 163365 374580 163366 374644
rect 163430 374580 163431 374644
rect 163365 374579 163431 374580
rect 165949 374644 166015 374645
rect 165949 374580 165950 374644
rect 166014 374580 166015 374644
rect 165949 374579 166015 374580
rect 153437 374508 153503 374509
rect 153437 374444 153438 374508
rect 153502 374444 153503 374508
rect 153437 374443 153503 374444
rect 156459 374508 156525 374509
rect 156459 374444 156460 374508
rect 156524 374444 156525 374508
rect 156459 374443 156525 374444
rect 158483 374508 158549 374509
rect 158483 374444 158484 374508
rect 158548 374444 158549 374508
rect 158483 374443 158549 374444
rect 160917 374508 160983 374509
rect 160917 374444 160918 374508
rect 160982 374444 160983 374508
rect 160917 374443 160983 374444
rect 125731 373692 125797 373693
rect 125731 373628 125732 373692
rect 125796 373628 125797 373692
rect 125731 373627 125797 373628
rect 128859 373692 128925 373693
rect 128859 373628 128860 373692
rect 128924 373628 128925 373692
rect 128859 373627 128925 373628
rect 131067 373692 131133 373693
rect 131067 373628 131068 373692
rect 131132 373628 131133 373692
rect 131067 373627 131133 373628
rect 133643 373692 133709 373693
rect 133643 373628 133644 373692
rect 133708 373628 133709 373692
rect 133643 373627 133709 373628
rect 136403 373692 136469 373693
rect 136403 373628 136404 373692
rect 136468 373628 136469 373692
rect 136403 373627 136469 373628
rect 139163 373692 139229 373693
rect 139163 373628 139164 373692
rect 139228 373628 139229 373692
rect 139163 373627 139229 373628
rect 141555 373692 141621 373693
rect 141555 373628 141556 373692
rect 141620 373628 141621 373692
rect 141555 373627 141621 373628
rect 151675 373692 151741 373693
rect 151675 373628 151676 373692
rect 151740 373628 151741 373692
rect 151675 373627 151741 373628
rect 122971 373420 123037 373421
rect 122971 373356 122972 373420
rect 123036 373356 123037 373420
rect 122971 373355 123037 373356
rect 118187 372468 118253 372469
rect 118187 372404 118188 372468
rect 118252 372404 118253 372468
rect 118187 372403 118253 372404
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 355308 117854 370338
rect 120954 357554 121574 373000
rect 120954 357318 120986 357554
rect 121222 357318 121306 357554
rect 121542 357318 121574 357554
rect 120954 357234 121574 357318
rect 120954 356998 120986 357234
rect 121222 356998 121306 357234
rect 121542 356998 121574 357234
rect 120954 355308 121574 356998
rect 127794 364394 128414 373000
rect 127794 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 128414 364394
rect 127794 364074 128414 364158
rect 127794 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 128414 364074
rect 127794 355308 128414 363838
rect 131514 366234 132134 373000
rect 131514 365998 131546 366234
rect 131782 365998 131866 366234
rect 132102 365998 132134 366234
rect 131514 365914 132134 365998
rect 131514 365678 131546 365914
rect 131782 365678 131866 365914
rect 132102 365678 132134 365914
rect 131514 355308 132134 365678
rect 135234 369954 135854 373000
rect 135234 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 135854 369954
rect 135234 369634 135854 369718
rect 135234 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 135854 369634
rect 135234 355308 135854 369398
rect 138954 356614 139574 373000
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 355308 139574 356058
rect 145794 363454 146414 373000
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 355308 146414 362898
rect 149514 367174 150134 373000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 355308 150134 366618
rect 153234 370894 153854 373000
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 355308 153854 370338
rect 156954 357554 157574 373000
rect 156954 357318 156986 357554
rect 157222 357318 157306 357554
rect 157542 357318 157574 357554
rect 156954 357234 157574 357318
rect 156954 356998 156986 357234
rect 157222 356998 157306 357234
rect 157542 356998 157574 357234
rect 156954 355308 157574 356998
rect 163794 364394 164414 373000
rect 163794 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 164414 364394
rect 163794 364074 164414 364158
rect 163794 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 164414 364074
rect 163794 355308 164414 363838
rect 167514 366234 168134 373000
rect 167514 365998 167546 366234
rect 167782 365998 167866 366234
rect 168102 365998 168134 366234
rect 167514 365914 168134 365998
rect 167514 365678 167546 365914
rect 167782 365678 167866 365914
rect 168102 365678 168134 365914
rect 167514 355308 168134 365678
rect 171234 369954 171854 373000
rect 171234 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 171854 369954
rect 171234 369634 171854 369718
rect 171234 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 171854 369634
rect 171234 355308 171854 369398
rect 174954 356614 175574 373000
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 355308 175574 356058
rect 181794 363454 182414 373000
rect 182958 371653 183018 374990
rect 183360 374370 183420 375020
rect 183326 374310 183420 374370
rect 183326 371653 183386 374310
rect 182955 371652 183021 371653
rect 182955 371588 182956 371652
rect 183020 371588 183021 371652
rect 182955 371587 183021 371588
rect 183323 371652 183389 371653
rect 183323 371588 183324 371652
rect 183388 371588 183389 371652
rect 183323 371587 183389 371588
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 178539 355332 178605 355333
rect 178539 355268 178540 355332
rect 178604 355268 178605 355332
rect 181794 355308 182414 362898
rect 185514 367174 186134 373000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 355308 186134 366618
rect 189234 370894 189854 373000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 355308 189854 370338
rect 192954 357554 193574 373000
rect 192954 357318 192986 357554
rect 193222 357318 193306 357554
rect 193542 357318 193574 357554
rect 192954 357234 193574 357318
rect 192954 356998 192986 357234
rect 193222 356998 193306 357234
rect 193542 356998 193574 357234
rect 190867 355332 190933 355333
rect 178539 355267 178605 355268
rect 190867 355268 190868 355332
rect 190932 355268 190933 355332
rect 192954 355308 193574 356998
rect 190867 355267 190933 355268
rect 178542 353970 178602 355267
rect 179643 354788 179709 354789
rect 179643 354724 179644 354788
rect 179708 354724 179709 354788
rect 179643 354723 179709 354724
rect 178464 353910 178602 353970
rect 179646 353970 179706 354723
rect 190870 353970 190930 355267
rect 179646 353910 179748 353970
rect 178464 353260 178524 353910
rect 179688 353260 179748 353910
rect 190840 353910 190930 353970
rect 190840 353260 190900 353910
rect 60272 345454 60620 345486
rect 60272 345218 60328 345454
rect 60564 345218 60620 345454
rect 60272 345134 60620 345218
rect 60272 344898 60328 345134
rect 60564 344898 60620 345134
rect 60272 344866 60620 344898
rect 196000 345454 196348 345486
rect 196000 345218 196056 345454
rect 196292 345218 196348 345454
rect 196000 345134 196348 345218
rect 196000 344898 196056 345134
rect 196292 344898 196348 345134
rect 196000 344866 196348 344898
rect 60952 327454 61300 327486
rect 60952 327218 61008 327454
rect 61244 327218 61300 327454
rect 60952 327134 61300 327218
rect 60952 326898 61008 327134
rect 61244 326898 61300 327134
rect 60952 326866 61300 326898
rect 195320 327454 195668 327486
rect 195320 327218 195376 327454
rect 195612 327218 195668 327454
rect 195320 327134 195668 327218
rect 195320 326898 195376 327134
rect 195612 326898 195668 327134
rect 195320 326866 195668 326898
rect 60272 309454 60620 309486
rect 60272 309218 60328 309454
rect 60564 309218 60620 309454
rect 60272 309134 60620 309218
rect 60272 308898 60328 309134
rect 60564 308898 60620 309134
rect 60272 308866 60620 308898
rect 196000 309454 196348 309486
rect 196000 309218 196056 309454
rect 196292 309218 196348 309454
rect 196000 309134 196348 309218
rect 196000 308898 196056 309134
rect 196292 308898 196348 309134
rect 196000 308866 196348 308898
rect 60952 291454 61300 291486
rect 60952 291218 61008 291454
rect 61244 291218 61300 291454
rect 60952 291134 61300 291218
rect 60952 290898 61008 291134
rect 61244 290898 61300 291134
rect 60952 290866 61300 290898
rect 195320 291454 195668 291486
rect 195320 291218 195376 291454
rect 195612 291218 195668 291454
rect 195320 291134 195668 291218
rect 195320 290898 195376 291134
rect 195612 290898 195668 291134
rect 195320 290866 195668 290898
rect 60272 273454 60620 273486
rect 60272 273218 60328 273454
rect 60564 273218 60620 273454
rect 60272 273134 60620 273218
rect 60272 272898 60328 273134
rect 60564 272898 60620 273134
rect 60272 272866 60620 272898
rect 196000 273454 196348 273486
rect 196000 273218 196056 273454
rect 196292 273218 196348 273454
rect 196000 273134 196348 273218
rect 196000 272898 196056 273134
rect 196292 272898 196348 273134
rect 196000 272866 196348 272898
rect 76056 269650 76116 270106
rect 76054 269590 76116 269650
rect 77144 269650 77204 270106
rect 78232 269650 78292 270106
rect 79592 269650 79652 270106
rect 80544 269650 80604 270106
rect 77144 269590 77218 269650
rect 78232 269590 78322 269650
rect 76054 269109 76114 269590
rect 77158 269109 77218 269590
rect 76051 269108 76117 269109
rect 76051 269044 76052 269108
rect 76116 269044 76117 269108
rect 76051 269043 76117 269044
rect 77155 269108 77221 269109
rect 77155 269044 77156 269108
rect 77220 269044 77221 269108
rect 77155 269043 77221 269044
rect 59514 260114 60134 268000
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 60134 260114
rect 59514 259794 60134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 60134 259794
rect 59514 250308 60134 259558
rect 63234 261954 63854 268000
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 63854 261954
rect 63234 261634 63854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 63854 261634
rect 63234 250308 63854 261398
rect 66954 265674 67574 268000
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 67574 265674
rect 66954 265354 67574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 67574 265354
rect 66954 250308 67574 265118
rect 73794 255454 74414 268000
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 250308 74414 254898
rect 77514 259174 78134 268000
rect 78262 266933 78322 269590
rect 79550 269590 79652 269650
rect 80470 269590 80604 269650
rect 81768 269650 81828 270106
rect 83128 269653 83188 270106
rect 83125 269652 83191 269653
rect 81768 269590 82002 269650
rect 79550 267613 79610 269590
rect 79547 267612 79613 267613
rect 79547 267548 79548 267612
rect 79612 267548 79613 267612
rect 79547 267547 79613 267548
rect 80470 266933 80530 269590
rect 78259 266932 78325 266933
rect 78259 266868 78260 266932
rect 78324 266868 78325 266932
rect 78259 266867 78325 266868
rect 80467 266932 80533 266933
rect 80467 266868 80468 266932
rect 80532 266868 80533 266932
rect 80467 266867 80533 266868
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 250308 78134 258618
rect 81234 262894 81854 268000
rect 81942 267477 82002 269590
rect 83125 269588 83126 269652
rect 83190 269588 83191 269652
rect 84216 269650 84276 270106
rect 85440 269650 85500 270106
rect 83125 269587 83191 269588
rect 83966 269590 84276 269650
rect 85438 269590 85500 269650
rect 86528 269650 86588 270106
rect 87616 269650 87676 270106
rect 86528 269590 86602 269650
rect 83966 267749 84026 269590
rect 85438 268157 85498 269590
rect 85435 268156 85501 268157
rect 85435 268092 85436 268156
rect 85500 268092 85501 268156
rect 85435 268091 85501 268092
rect 83963 267748 84029 267749
rect 83963 267684 83964 267748
rect 84028 267684 84029 267748
rect 83963 267683 84029 267684
rect 81939 267476 82005 267477
rect 81939 267412 81940 267476
rect 82004 267412 82005 267476
rect 81939 267411 82005 267412
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 250308 81854 262338
rect 84954 266614 85574 268000
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 86542 266389 86602 269590
rect 87462 269590 87676 269650
rect 88296 269650 88356 270106
rect 88704 269650 88764 270106
rect 90064 269650 90124 270106
rect 88296 269590 88442 269650
rect 88704 269590 88810 269650
rect 87462 267749 87522 269590
rect 87459 267748 87525 267749
rect 87459 267684 87460 267748
rect 87524 267684 87525 267748
rect 87459 267683 87525 267684
rect 88382 267205 88442 269590
rect 88379 267204 88445 267205
rect 88379 267140 88380 267204
rect 88444 267140 88445 267204
rect 88379 267139 88445 267140
rect 88750 266389 88810 269590
rect 90038 269590 90124 269650
rect 90744 269650 90804 270106
rect 91288 269650 91348 270106
rect 92376 269650 92436 270106
rect 93464 269650 93524 270106
rect 93600 269653 93660 270106
rect 94552 269653 94612 270106
rect 90744 269590 90834 269650
rect 91288 269590 91386 269650
rect 92376 269590 92490 269650
rect 90038 266389 90098 269590
rect 90774 269109 90834 269590
rect 90771 269108 90837 269109
rect 90771 269044 90772 269108
rect 90836 269044 90837 269108
rect 90771 269043 90837 269044
rect 91326 266661 91386 269590
rect 92430 268157 92490 269590
rect 93350 269590 93524 269650
rect 93597 269652 93663 269653
rect 92427 268156 92493 268157
rect 92427 268092 92428 268156
rect 92492 268092 92493 268156
rect 92427 268091 92493 268092
rect 91323 266660 91389 266661
rect 91323 266596 91324 266660
rect 91388 266596 91389 266660
rect 91323 266595 91389 266596
rect 84954 266294 85574 266378
rect 86539 266388 86605 266389
rect 86539 266324 86540 266388
rect 86604 266324 86605 266388
rect 86539 266323 86605 266324
rect 88747 266388 88813 266389
rect 88747 266324 88748 266388
rect 88812 266324 88813 266388
rect 88747 266323 88813 266324
rect 90035 266388 90101 266389
rect 90035 266324 90036 266388
rect 90100 266324 90101 266388
rect 90035 266323 90101 266324
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 250308 85574 266058
rect 91794 256394 92414 268000
rect 93350 266389 93410 269590
rect 93597 269588 93598 269652
rect 93662 269588 93663 269652
rect 93597 269587 93663 269588
rect 94549 269652 94615 269653
rect 94549 269588 94550 269652
rect 94614 269588 94615 269652
rect 95912 269650 95972 270106
rect 96048 269650 96108 270106
rect 97000 269650 97060 270106
rect 98088 269650 98148 270106
rect 98496 269650 98556 270106
rect 99448 269650 99508 270106
rect 95912 269590 95986 269650
rect 96048 269590 96170 269650
rect 97000 269590 97090 269650
rect 98088 269590 98194 269650
rect 98496 269590 98562 269650
rect 94549 269587 94615 269588
rect 95926 269109 95986 269590
rect 96110 269109 96170 269590
rect 95923 269108 95989 269109
rect 95923 269044 95924 269108
rect 95988 269044 95989 269108
rect 95923 269043 95989 269044
rect 96107 269108 96173 269109
rect 96107 269044 96108 269108
rect 96172 269044 96173 269108
rect 96107 269043 96173 269044
rect 93347 266388 93413 266389
rect 93347 266324 93348 266388
rect 93412 266324 93413 266388
rect 93347 266323 93413 266324
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 92414 256394
rect 91794 256074 92414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 92414 256074
rect 91794 250308 92414 255838
rect 95514 260114 96134 268000
rect 97030 266389 97090 269590
rect 98134 266389 98194 269590
rect 98502 269109 98562 269590
rect 99422 269590 99508 269650
rect 100672 269650 100732 270106
rect 101080 269650 101140 270106
rect 100672 269590 100770 269650
rect 99422 269109 99482 269590
rect 98499 269108 98565 269109
rect 98499 269044 98500 269108
rect 98564 269044 98565 269108
rect 98499 269043 98565 269044
rect 99419 269108 99485 269109
rect 99419 269044 99420 269108
rect 99484 269044 99485 269108
rect 99419 269043 99485 269044
rect 97027 266388 97093 266389
rect 97027 266324 97028 266388
rect 97092 266324 97093 266388
rect 97027 266323 97093 266324
rect 98131 266388 98197 266389
rect 98131 266324 98132 266388
rect 98196 266324 98197 266388
rect 98131 266323 98197 266324
rect 95514 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 96134 260114
rect 95514 259794 96134 259878
rect 95514 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 96134 259794
rect 95514 250308 96134 259558
rect 99234 261954 99854 268000
rect 100710 266525 100770 269590
rect 101078 269590 101140 269650
rect 101760 269650 101820 270106
rect 102848 269650 102908 270106
rect 103528 269650 103588 270106
rect 103936 269650 103996 270106
rect 101760 269590 101874 269650
rect 101078 267205 101138 269590
rect 101075 267204 101141 267205
rect 101075 267140 101076 267204
rect 101140 267140 101141 267204
rect 101075 267139 101141 267140
rect 100707 266524 100773 266525
rect 100707 266460 100708 266524
rect 100772 266460 100773 266524
rect 100707 266459 100773 266460
rect 101814 266389 101874 269590
rect 102734 269590 102908 269650
rect 103286 269590 103588 269650
rect 103838 269590 103996 269650
rect 105296 269650 105356 270106
rect 105976 269650 106036 270106
rect 105296 269590 105370 269650
rect 102734 267749 102794 269590
rect 103286 268157 103346 269590
rect 103283 268156 103349 268157
rect 103283 268092 103284 268156
rect 103348 268092 103349 268156
rect 103283 268091 103349 268092
rect 102731 267748 102797 267749
rect 102731 267684 102732 267748
rect 102796 267684 102797 267748
rect 102731 267683 102797 267684
rect 101811 266388 101877 266389
rect 101811 266324 101812 266388
rect 101876 266324 101877 266388
rect 101811 266323 101877 266324
rect 99234 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 99854 261954
rect 99234 261634 99854 261718
rect 99234 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 99854 261634
rect 99234 250308 99854 261398
rect 102954 265674 103574 268000
rect 103838 267069 103898 269590
rect 105310 267749 105370 269590
rect 105862 269590 106036 269650
rect 106384 269650 106444 270106
rect 107608 269925 107668 270106
rect 107605 269924 107671 269925
rect 107605 269860 107606 269924
rect 107670 269860 107671 269924
rect 107605 269859 107671 269860
rect 108288 269789 108348 270106
rect 108285 269788 108351 269789
rect 108285 269724 108286 269788
rect 108350 269724 108351 269788
rect 108285 269723 108351 269724
rect 108696 269653 108756 270106
rect 108693 269652 108759 269653
rect 106384 269590 106474 269650
rect 105307 267748 105373 267749
rect 105307 267684 105308 267748
rect 105372 267684 105373 267748
rect 105307 267683 105373 267684
rect 105862 267205 105922 269590
rect 106414 267749 106474 269590
rect 108693 269588 108694 269652
rect 108758 269588 108759 269652
rect 109784 269650 109844 270106
rect 111008 269925 111068 270106
rect 111005 269924 111071 269925
rect 111005 269860 111006 269924
rect 111070 269860 111071 269924
rect 111005 269859 111071 269860
rect 108693 269587 108759 269588
rect 109726 269590 109844 269650
rect 111144 269650 111204 270106
rect 112232 269650 112292 270106
rect 113320 269650 113380 270106
rect 113592 269650 113652 270106
rect 111144 269590 111258 269650
rect 109726 268565 109786 269590
rect 109723 268564 109789 268565
rect 109723 268500 109724 268564
rect 109788 268500 109789 268564
rect 109723 268499 109789 268500
rect 111198 268429 111258 269590
rect 112118 269590 112292 269650
rect 113222 269590 113380 269650
rect 113590 269590 113652 269650
rect 114408 269650 114468 270106
rect 115768 269650 115828 270106
rect 116040 269650 116100 270106
rect 114408 269590 114570 269650
rect 115768 269590 115858 269650
rect 111195 268428 111261 268429
rect 111195 268364 111196 268428
rect 111260 268364 111261 268428
rect 111195 268363 111261 268364
rect 106411 267748 106477 267749
rect 106411 267684 106412 267748
rect 106476 267684 106477 267748
rect 106411 267683 106477 267684
rect 105859 267204 105925 267205
rect 105859 267140 105860 267204
rect 105924 267140 105925 267204
rect 105859 267139 105925 267140
rect 103835 267068 103901 267069
rect 103835 267004 103836 267068
rect 103900 267004 103901 267068
rect 103835 267003 103901 267004
rect 102954 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 103574 265674
rect 102954 265354 103574 265438
rect 102954 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 103574 265354
rect 102954 250308 103574 265118
rect 109794 255454 110414 268000
rect 112118 266389 112178 269590
rect 113222 268021 113282 269590
rect 113590 268157 113650 269590
rect 113587 268156 113653 268157
rect 113587 268092 113588 268156
rect 113652 268092 113653 268156
rect 113587 268091 113653 268092
rect 113219 268020 113285 268021
rect 113219 267956 113220 268020
rect 113284 267956 113285 268020
rect 113219 267955 113285 267956
rect 112115 266388 112181 266389
rect 112115 266324 112116 266388
rect 112180 266324 112181 266388
rect 112115 266323 112181 266324
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 250308 110414 254898
rect 113514 259174 114134 268000
rect 114510 266389 114570 269590
rect 115798 268973 115858 269590
rect 115982 269590 116100 269650
rect 116992 269650 117052 270106
rect 118080 269650 118140 270106
rect 118488 269650 118548 270106
rect 119168 269650 119228 270106
rect 120936 269650 120996 270106
rect 116992 269590 117146 269650
rect 115795 268972 115861 268973
rect 115795 268908 115796 268972
rect 115860 268908 115861 268972
rect 115795 268907 115861 268908
rect 115982 267341 116042 269590
rect 117086 267749 117146 269590
rect 118006 269590 118140 269650
rect 118374 269590 118548 269650
rect 119110 269590 119228 269650
rect 120766 269590 120996 269650
rect 123520 269650 123580 270106
rect 125968 269650 126028 270106
rect 123520 269590 123586 269650
rect 118006 268837 118066 269590
rect 118003 268836 118069 268837
rect 118003 268772 118004 268836
rect 118068 268772 118069 268836
rect 118003 268771 118069 268772
rect 117083 267748 117149 267749
rect 117083 267684 117084 267748
rect 117148 267684 117149 267748
rect 117083 267683 117149 267684
rect 115979 267340 116045 267341
rect 115979 267276 115980 267340
rect 116044 267276 116045 267340
rect 115979 267275 116045 267276
rect 114507 266388 114573 266389
rect 114507 266324 114508 266388
rect 114572 266324 114573 266388
rect 114507 266323 114573 266324
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 250308 114134 258618
rect 117234 262894 117854 268000
rect 118374 267477 118434 269590
rect 119110 268701 119170 269590
rect 119107 268700 119173 268701
rect 119107 268636 119108 268700
rect 119172 268636 119173 268700
rect 119107 268635 119173 268636
rect 120766 267477 120826 269590
rect 118371 267476 118437 267477
rect 118371 267412 118372 267476
rect 118436 267412 118437 267476
rect 118371 267411 118437 267412
rect 120763 267476 120829 267477
rect 120763 267412 120764 267476
rect 120828 267412 120829 267476
rect 120763 267411 120829 267412
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 250308 117854 262338
rect 120954 266614 121574 268000
rect 123526 267749 123586 269590
rect 125918 269590 126028 269650
rect 128280 269650 128340 270106
rect 131000 269650 131060 270106
rect 133448 269789 133508 270106
rect 135896 269789 135956 270106
rect 138480 269789 138540 270106
rect 133445 269788 133511 269789
rect 133445 269724 133446 269788
rect 133510 269724 133511 269788
rect 133445 269723 133511 269724
rect 135893 269788 135959 269789
rect 135893 269724 135894 269788
rect 135958 269724 135959 269788
rect 135893 269723 135959 269724
rect 138477 269788 138543 269789
rect 138477 269724 138478 269788
rect 138542 269724 138543 269788
rect 138477 269723 138543 269724
rect 140928 269653 140988 270106
rect 143512 269653 143572 270106
rect 145960 269653 146020 270106
rect 128280 269590 128370 269650
rect 123523 267748 123589 267749
rect 123523 267684 123524 267748
rect 123588 267684 123589 267748
rect 123523 267683 123589 267684
rect 125918 267613 125978 269590
rect 128310 268157 128370 269590
rect 130886 269590 131060 269650
rect 140925 269652 140991 269653
rect 128307 268156 128373 268157
rect 128307 268092 128308 268156
rect 128372 268092 128373 268156
rect 128307 268091 128373 268092
rect 125915 267612 125981 267613
rect 125915 267548 125916 267612
rect 125980 267548 125981 267612
rect 125915 267547 125981 267548
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 250308 121574 266058
rect 127794 256394 128414 268000
rect 130886 267749 130946 269590
rect 140925 269588 140926 269652
rect 140990 269588 140991 269652
rect 140925 269587 140991 269588
rect 143509 269652 143575 269653
rect 143509 269588 143510 269652
rect 143574 269588 143575 269652
rect 143509 269587 143575 269588
rect 145957 269652 146023 269653
rect 145957 269588 145958 269652
rect 146022 269588 146023 269652
rect 148544 269650 148604 270106
rect 150992 269650 151052 270106
rect 148544 269590 148610 269650
rect 145957 269587 146023 269588
rect 130883 267748 130949 267749
rect 130883 267684 130884 267748
rect 130948 267684 130949 267748
rect 130883 267683 130949 267684
rect 127794 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 128414 256394
rect 127794 256074 128414 256158
rect 127794 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 128414 256074
rect 127794 250308 128414 255838
rect 131514 260114 132134 268000
rect 131514 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 132134 260114
rect 131514 259794 132134 259878
rect 131514 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 132134 259794
rect 131514 250308 132134 259558
rect 135234 261954 135854 268000
rect 135234 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 135854 261954
rect 135234 261634 135854 261718
rect 135234 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 135854 261634
rect 135234 250308 135854 261398
rect 138954 265674 139574 268000
rect 138954 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 139574 265674
rect 138954 265354 139574 265438
rect 138954 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 139574 265354
rect 138954 250308 139574 265118
rect 145794 255454 146414 268000
rect 148550 266389 148610 269590
rect 150942 269590 151052 269650
rect 153440 269650 153500 270106
rect 155888 269650 155948 270106
rect 158472 269650 158532 270106
rect 160920 269650 160980 270106
rect 153440 269590 153578 269650
rect 155888 269590 155970 269650
rect 158472 269590 158546 269650
rect 148547 266388 148613 266389
rect 148547 266324 148548 266388
rect 148612 266324 148613 266388
rect 148547 266323 148613 266324
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 250308 146414 254898
rect 149514 259174 150134 268000
rect 150942 267613 151002 269590
rect 153518 268157 153578 269590
rect 153515 268156 153581 268157
rect 153515 268092 153516 268156
rect 153580 268092 153581 268156
rect 153515 268091 153581 268092
rect 150939 267612 151005 267613
rect 150939 267548 150940 267612
rect 151004 267548 151005 267612
rect 150939 267547 151005 267548
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 250308 150134 258618
rect 153234 262894 153854 268000
rect 155910 267749 155970 269590
rect 155907 267748 155973 267749
rect 155907 267684 155908 267748
rect 155972 267684 155973 267748
rect 155907 267683 155973 267684
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 250308 153854 262338
rect 156954 266614 157574 268000
rect 158486 267749 158546 269590
rect 160878 269590 160980 269650
rect 163368 269650 163428 270106
rect 165952 269650 166012 270106
rect 183224 269650 183284 270106
rect 163368 269590 163514 269650
rect 165952 269590 166090 269650
rect 158483 267748 158549 267749
rect 158483 267684 158484 267748
rect 158548 267684 158549 267748
rect 158483 267683 158549 267684
rect 160878 267477 160938 269590
rect 163454 267749 163514 269590
rect 163451 267748 163517 267749
rect 163451 267684 163452 267748
rect 163516 267684 163517 267748
rect 163451 267683 163517 267684
rect 160875 267476 160941 267477
rect 160875 267412 160876 267476
rect 160940 267412 160941 267476
rect 160875 267411 160941 267412
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 250308 157574 266058
rect 163794 256394 164414 268000
rect 166030 267477 166090 269590
rect 183142 269590 183284 269650
rect 183360 269650 183420 270106
rect 183360 269590 183570 269650
rect 166027 267476 166093 267477
rect 166027 267412 166028 267476
rect 166092 267412 166093 267476
rect 166027 267411 166093 267412
rect 163794 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 164414 256394
rect 163794 256074 164414 256158
rect 163794 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 164414 256074
rect 163794 250308 164414 255838
rect 167514 260114 168134 268000
rect 167514 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 168134 260114
rect 167514 259794 168134 259878
rect 167514 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 168134 259794
rect 167514 250308 168134 259558
rect 171234 261954 171854 268000
rect 171234 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 171854 261954
rect 171234 261634 171854 261718
rect 171234 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 171854 261634
rect 171234 250308 171854 261398
rect 174954 265674 175574 268000
rect 174954 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 175574 265674
rect 174954 265354 175574 265438
rect 174954 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 175574 265354
rect 174954 250308 175574 265118
rect 181794 255454 182414 268000
rect 183142 267341 183202 269590
rect 183510 267477 183570 269590
rect 183507 267476 183573 267477
rect 183507 267412 183508 267476
rect 183572 267412 183573 267476
rect 183507 267411 183573 267412
rect 183139 267340 183205 267341
rect 183139 267276 183140 267340
rect 183204 267276 183205 267340
rect 183139 267275 183205 267276
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 250308 182414 254898
rect 185514 259174 186134 268000
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 250308 186134 258618
rect 189234 262894 189854 268000
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 250308 189854 262338
rect 192954 266614 193574 268000
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 250308 193574 266058
rect 178539 249932 178605 249933
rect 178539 249868 178540 249932
rect 178604 249868 178605 249932
rect 178539 249867 178605 249868
rect 179643 249932 179709 249933
rect 179643 249868 179644 249932
rect 179708 249868 179709 249932
rect 179643 249867 179709 249868
rect 190867 249932 190933 249933
rect 190867 249868 190868 249932
rect 190932 249868 190933 249932
rect 190867 249867 190933 249868
rect 178542 248430 178602 249867
rect 178464 248370 178602 248430
rect 179646 248430 179706 249867
rect 190870 248430 190930 249867
rect 179646 248370 179748 248430
rect 178464 248202 178524 248370
rect 179688 248202 179748 248370
rect 190840 248370 190930 248430
rect 190840 248202 190900 248370
rect 60272 237454 60620 237486
rect 60272 237218 60328 237454
rect 60564 237218 60620 237454
rect 60272 237134 60620 237218
rect 60272 236898 60328 237134
rect 60564 236898 60620 237134
rect 60272 236866 60620 236898
rect 196000 237454 196348 237486
rect 196000 237218 196056 237454
rect 196292 237218 196348 237454
rect 196000 237134 196348 237218
rect 196000 236898 196056 237134
rect 196292 236898 196348 237134
rect 196000 236866 196348 236898
rect 60952 219454 61300 219486
rect 60952 219218 61008 219454
rect 61244 219218 61300 219454
rect 60952 219134 61300 219218
rect 60952 218898 61008 219134
rect 61244 218898 61300 219134
rect 60952 218866 61300 218898
rect 195320 219454 195668 219486
rect 195320 219218 195376 219454
rect 195612 219218 195668 219454
rect 195320 219134 195668 219218
rect 195320 218898 195376 219134
rect 195612 218898 195668 219134
rect 195320 218866 195668 218898
rect 60272 201454 60620 201486
rect 60272 201218 60328 201454
rect 60564 201218 60620 201454
rect 60272 201134 60620 201218
rect 60272 200898 60328 201134
rect 60564 200898 60620 201134
rect 60272 200866 60620 200898
rect 196000 201454 196348 201486
rect 196000 201218 196056 201454
rect 196292 201218 196348 201454
rect 196000 201134 196348 201218
rect 196000 200898 196056 201134
rect 196292 200898 196348 201134
rect 196000 200866 196348 200898
rect 60952 183454 61300 183486
rect 60952 183218 61008 183454
rect 61244 183218 61300 183454
rect 60952 183134 61300 183218
rect 60952 182898 61008 183134
rect 61244 182898 61300 183134
rect 60952 182866 61300 182898
rect 195320 183454 195668 183486
rect 195320 183218 195376 183454
rect 195612 183218 195668 183454
rect 195320 183134 195668 183218
rect 195320 182898 195376 183134
rect 195612 182898 195668 183134
rect 195320 182866 195668 182898
rect 76056 164930 76116 165106
rect 76054 164870 76116 164930
rect 77144 164930 77204 165106
rect 78232 164930 78292 165106
rect 79592 164930 79652 165106
rect 80544 164930 80604 165106
rect 77144 164870 77218 164930
rect 78232 164870 78322 164930
rect 59514 152114 60134 163000
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 60134 152114
rect 59514 151794 60134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 60134 151794
rect 59514 145308 60134 151558
rect 63234 153954 63854 163000
rect 63234 153718 63266 153954
rect 63502 153718 63586 153954
rect 63822 153718 63854 153954
rect 63234 153634 63854 153718
rect 63234 153398 63266 153634
rect 63502 153398 63586 153634
rect 63822 153398 63854 153634
rect 63234 145308 63854 153398
rect 66954 157674 67574 163000
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 67574 157674
rect 66954 157354 67574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 67574 157354
rect 66954 145308 67574 157118
rect 73794 147454 74414 163000
rect 76054 162757 76114 164870
rect 76051 162756 76117 162757
rect 76051 162692 76052 162756
rect 76116 162692 76117 162756
rect 76051 162691 76117 162692
rect 77158 162213 77218 164870
rect 77155 162212 77221 162213
rect 77155 162148 77156 162212
rect 77220 162148 77221 162212
rect 77155 162147 77221 162148
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 145308 74414 146898
rect 77514 151174 78134 163000
rect 78262 162757 78322 164870
rect 79550 164870 79652 164930
rect 80470 164870 80604 164930
rect 81768 164930 81828 165106
rect 83128 164930 83188 165106
rect 84216 164930 84276 165106
rect 85440 164930 85500 165106
rect 81768 164870 82002 164930
rect 79550 162757 79610 164870
rect 80470 162757 80530 164870
rect 78259 162756 78325 162757
rect 78259 162692 78260 162756
rect 78324 162692 78325 162756
rect 78259 162691 78325 162692
rect 79547 162756 79613 162757
rect 79547 162692 79548 162756
rect 79612 162692 79613 162756
rect 79547 162691 79613 162692
rect 80467 162756 80533 162757
rect 80467 162692 80468 162756
rect 80532 162692 80533 162756
rect 80467 162691 80533 162692
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 145308 78134 150618
rect 81234 154894 81854 163000
rect 81942 162757 82002 164870
rect 83046 164870 83188 164930
rect 83966 164870 84276 164930
rect 85438 164870 85500 164930
rect 86528 164930 86588 165106
rect 87616 164930 87676 165106
rect 88296 164930 88356 165106
rect 88704 164930 88764 165106
rect 90064 164930 90124 165106
rect 86528 164870 86602 164930
rect 87616 164870 87706 164930
rect 88296 164870 88442 164930
rect 88704 164870 88810 164930
rect 83046 162757 83106 164870
rect 81939 162756 82005 162757
rect 81939 162692 81940 162756
rect 82004 162692 82005 162756
rect 81939 162691 82005 162692
rect 83043 162756 83109 162757
rect 83043 162692 83044 162756
rect 83108 162692 83109 162756
rect 83043 162691 83109 162692
rect 83966 161530 84026 164870
rect 85438 163165 85498 164870
rect 85435 163164 85501 163165
rect 85435 163100 85436 163164
rect 85500 163100 85501 163164
rect 85435 163099 85501 163100
rect 84147 161532 84213 161533
rect 84147 161530 84148 161532
rect 83966 161470 84148 161530
rect 84147 161468 84148 161470
rect 84212 161468 84213 161532
rect 84147 161467 84213 161468
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 145308 81854 154338
rect 84954 158614 85574 163000
rect 86542 162757 86602 164870
rect 87646 162757 87706 164870
rect 86539 162756 86605 162757
rect 86539 162692 86540 162756
rect 86604 162692 86605 162756
rect 86539 162691 86605 162692
rect 87643 162756 87709 162757
rect 87643 162692 87644 162756
rect 87708 162692 87709 162756
rect 87643 162691 87709 162692
rect 88382 162213 88442 164870
rect 88750 162757 88810 164870
rect 90038 164870 90124 164930
rect 90744 164930 90804 165106
rect 91288 164930 91348 165106
rect 92376 164930 92436 165106
rect 93464 164930 93524 165106
rect 90744 164870 90834 164930
rect 91288 164870 91386 164930
rect 90038 162757 90098 164870
rect 90774 162757 90834 164870
rect 91326 162757 91386 164870
rect 91510 164870 92436 164930
rect 93350 164870 93524 164930
rect 93600 164930 93660 165106
rect 94552 164930 94612 165106
rect 93600 164870 93778 164930
rect 88747 162756 88813 162757
rect 88747 162692 88748 162756
rect 88812 162692 88813 162756
rect 88747 162691 88813 162692
rect 90035 162756 90101 162757
rect 90035 162692 90036 162756
rect 90100 162692 90101 162756
rect 90035 162691 90101 162692
rect 90771 162756 90837 162757
rect 90771 162692 90772 162756
rect 90836 162692 90837 162756
rect 90771 162691 90837 162692
rect 91323 162756 91389 162757
rect 91323 162692 91324 162756
rect 91388 162692 91389 162756
rect 91323 162691 91389 162692
rect 91510 162213 91570 164870
rect 88379 162212 88445 162213
rect 88379 162148 88380 162212
rect 88444 162148 88445 162212
rect 88379 162147 88445 162148
rect 91507 162212 91573 162213
rect 91507 162148 91508 162212
rect 91572 162148 91573 162212
rect 91507 162147 91573 162148
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 145308 85574 158058
rect 91794 148394 92414 163000
rect 93350 162757 93410 164870
rect 93718 162757 93778 164870
rect 94454 164870 94612 164930
rect 95912 164930 95972 165106
rect 96048 164930 96108 165106
rect 97000 164930 97060 165106
rect 98088 164930 98148 165106
rect 98496 164930 98556 165106
rect 99448 164930 99508 165106
rect 95912 164870 95986 164930
rect 96048 164870 96170 164930
rect 97000 164870 97090 164930
rect 98088 164870 98194 164930
rect 98496 164870 98562 164930
rect 94454 162757 94514 164870
rect 95926 163165 95986 164870
rect 96110 164797 96170 164870
rect 96107 164796 96173 164797
rect 96107 164732 96108 164796
rect 96172 164732 96173 164796
rect 96107 164731 96173 164732
rect 95923 163164 95989 163165
rect 95923 163100 95924 163164
rect 95988 163100 95989 163164
rect 95923 163099 95989 163100
rect 93347 162756 93413 162757
rect 93347 162692 93348 162756
rect 93412 162692 93413 162756
rect 93347 162691 93413 162692
rect 93715 162756 93781 162757
rect 93715 162692 93716 162756
rect 93780 162692 93781 162756
rect 93715 162691 93781 162692
rect 94451 162756 94517 162757
rect 94451 162692 94452 162756
rect 94516 162692 94517 162756
rect 94451 162691 94517 162692
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 92414 148394
rect 91794 148074 92414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 92414 148074
rect 91794 145308 92414 147838
rect 95514 152114 96134 163000
rect 97030 162757 97090 164870
rect 98134 162757 98194 164870
rect 98502 164253 98562 164870
rect 99422 164870 99508 164930
rect 100672 164930 100732 165106
rect 101080 164930 101140 165106
rect 100672 164870 100770 164930
rect 98499 164252 98565 164253
rect 98499 164188 98500 164252
rect 98564 164188 98565 164252
rect 98499 164187 98565 164188
rect 99422 163165 99482 164870
rect 99419 163164 99485 163165
rect 99419 163100 99420 163164
rect 99484 163100 99485 163164
rect 99419 163099 99485 163100
rect 97027 162756 97093 162757
rect 97027 162692 97028 162756
rect 97092 162692 97093 162756
rect 97027 162691 97093 162692
rect 98131 162756 98197 162757
rect 98131 162692 98132 162756
rect 98196 162692 98197 162756
rect 98131 162691 98197 162692
rect 95514 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 96134 152114
rect 95514 151794 96134 151878
rect 95514 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 96134 151794
rect 95514 145308 96134 151558
rect 99234 153954 99854 163000
rect 100710 162757 100770 164870
rect 101078 164870 101140 164930
rect 101760 164930 101820 165106
rect 102848 164930 102908 165106
rect 101760 164870 101874 164930
rect 101078 164253 101138 164870
rect 101075 164252 101141 164253
rect 101075 164188 101076 164252
rect 101140 164188 101141 164252
rect 101075 164187 101141 164188
rect 100707 162756 100773 162757
rect 100707 162692 100708 162756
rect 100772 162692 100773 162756
rect 100707 162691 100773 162692
rect 101814 162213 101874 164870
rect 102734 164870 102908 164930
rect 102734 162757 102794 164870
rect 103528 164661 103588 165106
rect 103936 164930 103996 165106
rect 103838 164870 103996 164930
rect 105296 164930 105356 165106
rect 105296 164870 105370 164930
rect 103525 164660 103591 164661
rect 103525 164596 103526 164660
rect 103590 164596 103591 164660
rect 103525 164595 103591 164596
rect 102731 162756 102797 162757
rect 102731 162692 102732 162756
rect 102796 162692 102797 162756
rect 102731 162691 102797 162692
rect 101811 162212 101877 162213
rect 101811 162148 101812 162212
rect 101876 162148 101877 162212
rect 101811 162147 101877 162148
rect 99234 153718 99266 153954
rect 99502 153718 99586 153954
rect 99822 153718 99854 153954
rect 99234 153634 99854 153718
rect 99234 153398 99266 153634
rect 99502 153398 99586 153634
rect 99822 153398 99854 153634
rect 99234 145308 99854 153398
rect 102954 157674 103574 163000
rect 103838 162757 103898 164870
rect 105310 162757 105370 164870
rect 105976 164661 106036 165106
rect 106384 164930 106444 165106
rect 107608 164930 107668 165106
rect 108288 164930 108348 165106
rect 108696 164930 108756 165106
rect 109784 164930 109844 165106
rect 106384 164870 106474 164930
rect 105973 164660 106039 164661
rect 105973 164596 105974 164660
rect 106038 164596 106039 164660
rect 105973 164595 106039 164596
rect 106414 162757 106474 164870
rect 107518 164870 107668 164930
rect 108254 164870 108348 164930
rect 108622 164870 108756 164930
rect 109542 164870 109844 164930
rect 111008 164930 111068 165106
rect 111144 164930 111204 165106
rect 112232 164930 112292 165106
rect 113320 164930 113380 165106
rect 113592 164930 113652 165106
rect 111008 164870 111074 164930
rect 111144 164870 111258 164930
rect 103835 162756 103901 162757
rect 103835 162692 103836 162756
rect 103900 162692 103901 162756
rect 103835 162691 103901 162692
rect 105307 162756 105373 162757
rect 105307 162692 105308 162756
rect 105372 162692 105373 162756
rect 105307 162691 105373 162692
rect 106411 162756 106477 162757
rect 106411 162692 106412 162756
rect 106476 162692 106477 162756
rect 106411 162691 106477 162692
rect 107518 162213 107578 164870
rect 108254 164253 108314 164870
rect 108251 164252 108317 164253
rect 108251 164188 108252 164252
rect 108316 164188 108317 164252
rect 108251 164187 108317 164188
rect 108622 162757 108682 164870
rect 109542 162757 109602 164870
rect 108619 162756 108685 162757
rect 108619 162692 108620 162756
rect 108684 162692 108685 162756
rect 108619 162691 108685 162692
rect 109539 162756 109605 162757
rect 109539 162692 109540 162756
rect 109604 162692 109605 162756
rect 109539 162691 109605 162692
rect 107515 162212 107581 162213
rect 107515 162148 107516 162212
rect 107580 162148 107581 162212
rect 107515 162147 107581 162148
rect 102954 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 103574 157674
rect 102954 157354 103574 157438
rect 102954 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 103574 157354
rect 102954 145308 103574 157118
rect 109794 147454 110414 163000
rect 111014 162213 111074 164870
rect 111198 162757 111258 164870
rect 112118 164870 112292 164930
rect 113222 164870 113380 164930
rect 113590 164870 113652 164930
rect 114408 164930 114468 165106
rect 115768 164930 115828 165106
rect 116040 164930 116100 165106
rect 114408 164870 114570 164930
rect 115768 164870 115858 164930
rect 112118 162757 112178 164870
rect 113222 162757 113282 164870
rect 113590 163165 113650 164870
rect 113587 163164 113653 163165
rect 113587 163100 113588 163164
rect 113652 163100 113653 163164
rect 113587 163099 113653 163100
rect 111195 162756 111261 162757
rect 111195 162692 111196 162756
rect 111260 162692 111261 162756
rect 111195 162691 111261 162692
rect 112115 162756 112181 162757
rect 112115 162692 112116 162756
rect 112180 162692 112181 162756
rect 112115 162691 112181 162692
rect 113219 162756 113285 162757
rect 113219 162692 113220 162756
rect 113284 162692 113285 162756
rect 113219 162691 113285 162692
rect 111011 162212 111077 162213
rect 111011 162148 111012 162212
rect 111076 162148 111077 162212
rect 111011 162147 111077 162148
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 145308 110414 146898
rect 113514 151174 114134 163000
rect 114510 162077 114570 164870
rect 115798 162757 115858 164870
rect 115982 164870 116100 164930
rect 115982 162757 116042 164870
rect 116992 164661 117052 165106
rect 118080 164930 118140 165106
rect 118488 164930 118548 165106
rect 119168 164930 119228 165106
rect 120936 164930 120996 165106
rect 123520 164930 123580 165106
rect 125968 164930 126028 165106
rect 118006 164870 118140 164930
rect 118374 164870 118548 164930
rect 119110 164870 119228 164930
rect 120766 164870 120996 164930
rect 123342 164870 123580 164930
rect 125918 164870 126028 164930
rect 128280 164930 128340 165106
rect 131000 164930 131060 165106
rect 128280 164870 128370 164930
rect 116989 164660 117055 164661
rect 116989 164596 116990 164660
rect 117054 164596 117055 164660
rect 116989 164595 117055 164596
rect 115795 162756 115861 162757
rect 115795 162692 115796 162756
rect 115860 162692 115861 162756
rect 115795 162691 115861 162692
rect 115979 162756 116045 162757
rect 115979 162692 115980 162756
rect 116044 162692 116045 162756
rect 115979 162691 116045 162692
rect 114507 162076 114573 162077
rect 114507 162012 114508 162076
rect 114572 162012 114573 162076
rect 114507 162011 114573 162012
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 145308 114134 150618
rect 117234 154894 117854 163000
rect 118006 162757 118066 164870
rect 118374 162757 118434 164870
rect 119110 162757 119170 164870
rect 120766 162757 120826 164870
rect 123342 164250 123402 164870
rect 122606 164190 123402 164250
rect 118003 162756 118069 162757
rect 118003 162692 118004 162756
rect 118068 162692 118069 162756
rect 118003 162691 118069 162692
rect 118371 162756 118437 162757
rect 118371 162692 118372 162756
rect 118436 162692 118437 162756
rect 118371 162691 118437 162692
rect 119107 162756 119173 162757
rect 119107 162692 119108 162756
rect 119172 162692 119173 162756
rect 119107 162691 119173 162692
rect 120763 162756 120829 162757
rect 120763 162692 120764 162756
rect 120828 162692 120829 162756
rect 120763 162691 120829 162692
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 145308 117854 154338
rect 120954 158614 121574 163000
rect 122606 162757 122666 164190
rect 125918 162757 125978 164870
rect 128310 163165 128370 164870
rect 130886 164870 131060 164930
rect 133448 164930 133508 165106
rect 135896 164930 135956 165106
rect 138480 164930 138540 165106
rect 133448 164870 133522 164930
rect 135896 164870 136098 164930
rect 128307 163164 128373 163165
rect 128307 163100 128308 163164
rect 128372 163100 128373 163164
rect 128307 163099 128373 163100
rect 122603 162756 122669 162757
rect 122603 162692 122604 162756
rect 122668 162692 122669 162756
rect 122603 162691 122669 162692
rect 125915 162756 125981 162757
rect 125915 162692 125916 162756
rect 125980 162692 125981 162756
rect 125915 162691 125981 162692
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 145308 121574 158058
rect 127794 148394 128414 163000
rect 130886 162757 130946 164870
rect 130883 162756 130949 162757
rect 130883 162692 130884 162756
rect 130948 162692 130949 162756
rect 130883 162691 130949 162692
rect 127794 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 128414 148394
rect 127794 148074 128414 148158
rect 127794 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 128414 148074
rect 127794 145308 128414 147838
rect 131514 152114 132134 163000
rect 133462 162757 133522 164870
rect 133459 162756 133525 162757
rect 133459 162692 133460 162756
rect 133524 162692 133525 162756
rect 133459 162691 133525 162692
rect 131514 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 132134 152114
rect 131514 151794 132134 151878
rect 131514 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 132134 151794
rect 131514 145308 132134 151558
rect 135234 153954 135854 163000
rect 136038 162349 136098 164870
rect 138430 164870 138540 164930
rect 138430 164389 138490 164870
rect 140928 164797 140988 165106
rect 143512 164930 143572 165106
rect 145960 164930 146020 165106
rect 148544 164930 148604 165106
rect 150992 164930 151052 165106
rect 143512 164870 143642 164930
rect 145960 164870 146034 164930
rect 148544 164870 148610 164930
rect 140925 164796 140991 164797
rect 140925 164732 140926 164796
rect 140990 164732 140991 164796
rect 140925 164731 140991 164732
rect 138427 164388 138493 164389
rect 138427 164324 138428 164388
rect 138492 164324 138493 164388
rect 138427 164323 138493 164324
rect 143582 164117 143642 164870
rect 145974 164253 146034 164870
rect 148550 164253 148610 164870
rect 150942 164870 151052 164930
rect 150942 164253 151002 164870
rect 153440 164661 153500 165106
rect 155888 164930 155948 165106
rect 158472 164930 158532 165106
rect 160920 164930 160980 165106
rect 155888 164870 155970 164930
rect 158472 164870 158546 164930
rect 153437 164660 153503 164661
rect 153437 164596 153438 164660
rect 153502 164596 153503 164660
rect 153437 164595 153503 164596
rect 145971 164252 146037 164253
rect 145971 164188 145972 164252
rect 146036 164188 146037 164252
rect 145971 164187 146037 164188
rect 148547 164252 148613 164253
rect 148547 164188 148548 164252
rect 148612 164188 148613 164252
rect 148547 164187 148613 164188
rect 150939 164252 151005 164253
rect 150939 164188 150940 164252
rect 151004 164188 151005 164252
rect 150939 164187 151005 164188
rect 143579 164116 143645 164117
rect 143579 164052 143580 164116
rect 143644 164052 143645 164116
rect 143579 164051 143645 164052
rect 136035 162348 136101 162349
rect 136035 162284 136036 162348
rect 136100 162284 136101 162348
rect 136035 162283 136101 162284
rect 135234 153718 135266 153954
rect 135502 153718 135586 153954
rect 135822 153718 135854 153954
rect 135234 153634 135854 153718
rect 135234 153398 135266 153634
rect 135502 153398 135586 153634
rect 135822 153398 135854 153634
rect 135234 145308 135854 153398
rect 138954 157674 139574 163000
rect 138954 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 139574 157674
rect 138954 157354 139574 157438
rect 138954 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 139574 157354
rect 138954 145308 139574 157118
rect 145794 147454 146414 163000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 145308 146414 146898
rect 149514 151174 150134 163000
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 145308 150134 150618
rect 153234 154894 153854 163000
rect 155910 162485 155970 164870
rect 155907 162484 155973 162485
rect 155907 162420 155908 162484
rect 155972 162420 155973 162484
rect 155907 162419 155973 162420
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 145308 153854 154338
rect 156954 158614 157574 163000
rect 158486 162621 158546 164870
rect 160878 164870 160980 164930
rect 158483 162620 158549 162621
rect 158483 162556 158484 162620
rect 158548 162556 158549 162620
rect 158483 162555 158549 162556
rect 160878 161941 160938 164870
rect 163368 164661 163428 165106
rect 165952 164930 166012 165106
rect 183224 164930 183284 165106
rect 165952 164870 166090 164930
rect 163365 164660 163431 164661
rect 163365 164596 163366 164660
rect 163430 164596 163431 164660
rect 163365 164595 163431 164596
rect 160875 161940 160941 161941
rect 160875 161876 160876 161940
rect 160940 161876 160941 161940
rect 160875 161875 160941 161876
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 145308 157574 158058
rect 163794 148394 164414 163000
rect 166030 162621 166090 164870
rect 183142 164870 183284 164930
rect 183360 164930 183420 165106
rect 183360 164870 183570 164930
rect 166027 162620 166093 162621
rect 166027 162556 166028 162620
rect 166092 162556 166093 162620
rect 166027 162555 166093 162556
rect 163794 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 164414 148394
rect 163794 148074 164414 148158
rect 163794 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 164414 148074
rect 163794 145308 164414 147838
rect 167514 152114 168134 163000
rect 167514 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 168134 152114
rect 167514 151794 168134 151878
rect 167514 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 168134 151794
rect 167514 145308 168134 151558
rect 171234 153954 171854 163000
rect 171234 153718 171266 153954
rect 171502 153718 171586 153954
rect 171822 153718 171854 153954
rect 171234 153634 171854 153718
rect 171234 153398 171266 153634
rect 171502 153398 171586 153634
rect 171822 153398 171854 153634
rect 171234 145308 171854 153398
rect 174954 157674 175574 163000
rect 174954 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 175574 157674
rect 174954 157354 175574 157438
rect 174954 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 175574 157354
rect 174954 145308 175574 157118
rect 181794 147454 182414 163000
rect 183142 162485 183202 164870
rect 183510 162757 183570 164870
rect 196574 163437 196634 478483
rect 197859 478412 197925 478413
rect 197859 478348 197860 478412
rect 197924 478348 197925 478412
rect 197859 478347 197925 478348
rect 196755 468484 196821 468485
rect 196755 468420 196756 468484
rect 196820 468420 196821 468484
rect 196755 468419 196821 468420
rect 196758 266253 196818 468419
rect 196755 266252 196821 266253
rect 196755 266188 196756 266252
rect 196820 266188 196821 266252
rect 196755 266187 196821 266188
rect 196571 163436 196637 163437
rect 196571 163372 196572 163436
rect 196636 163372 196637 163436
rect 196571 163371 196637 163372
rect 183507 162756 183573 162757
rect 183507 162692 183508 162756
rect 183572 162692 183573 162756
rect 183507 162691 183573 162692
rect 183139 162484 183205 162485
rect 183139 162420 183140 162484
rect 183204 162420 183205 162484
rect 183139 162419 183205 162420
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 145308 182414 146898
rect 185514 151174 186134 163000
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 145308 186134 150618
rect 189234 154894 189854 163000
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 145308 189854 154338
rect 192954 158614 193574 163000
rect 196758 162077 196818 266187
rect 196755 162076 196821 162077
rect 196755 162012 196756 162076
rect 196820 162012 196821 162076
rect 196755 162011 196821 162012
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 190867 145484 190933 145485
rect 190867 145420 190868 145484
rect 190932 145420 190933 145484
rect 190867 145419 190933 145420
rect 178539 144940 178605 144941
rect 178539 144876 178540 144940
rect 178604 144876 178605 144940
rect 178539 144875 178605 144876
rect 179643 144940 179709 144941
rect 179643 144876 179644 144940
rect 179708 144876 179709 144940
rect 179643 144875 179709 144876
rect 178542 143850 178602 144875
rect 178464 143790 178602 143850
rect 179646 143850 179706 144875
rect 190870 143850 190930 145419
rect 192954 145308 193574 158058
rect 179646 143790 179748 143850
rect 178464 143202 178524 143790
rect 179688 143202 179748 143790
rect 190840 143790 190930 143850
rect 190840 143202 190900 143790
rect 60272 129454 60620 129486
rect 60272 129218 60328 129454
rect 60564 129218 60620 129454
rect 60272 129134 60620 129218
rect 60272 128898 60328 129134
rect 60564 128898 60620 129134
rect 60272 128866 60620 128898
rect 196000 129454 196348 129486
rect 196000 129218 196056 129454
rect 196292 129218 196348 129454
rect 196000 129134 196348 129218
rect 196000 128898 196056 129134
rect 196292 128898 196348 129134
rect 196000 128866 196348 128898
rect 60952 111454 61300 111486
rect 60952 111218 61008 111454
rect 61244 111218 61300 111454
rect 60952 111134 61300 111218
rect 60952 110898 61008 111134
rect 61244 110898 61300 111134
rect 60952 110866 61300 110898
rect 195320 111454 195668 111486
rect 195320 111218 195376 111454
rect 195612 111218 195668 111454
rect 195320 111134 195668 111218
rect 195320 110898 195376 111134
rect 195612 110898 195668 111134
rect 195320 110866 195668 110898
rect 60272 93454 60620 93486
rect 60272 93218 60328 93454
rect 60564 93218 60620 93454
rect 60272 93134 60620 93218
rect 60272 92898 60328 93134
rect 60564 92898 60620 93134
rect 60272 92866 60620 92898
rect 196000 93454 196348 93486
rect 196000 93218 196056 93454
rect 196292 93218 196348 93454
rect 196000 93134 196348 93218
rect 196000 92898 196056 93134
rect 196292 92898 196348 93134
rect 196000 92866 196348 92898
rect 60952 75454 61300 75486
rect 60952 75218 61008 75454
rect 61244 75218 61300 75454
rect 60952 75134 61300 75218
rect 60952 74898 61008 75134
rect 61244 74898 61300 75134
rect 60952 74866 61300 74898
rect 195320 75454 195668 75486
rect 195320 75218 195376 75454
rect 195612 75218 195668 75454
rect 195320 75134 195668 75218
rect 195320 74898 195376 75134
rect 195612 74898 195668 75134
rect 195320 74866 195668 74898
rect 76056 59530 76116 60106
rect 77144 59805 77204 60106
rect 77141 59804 77207 59805
rect 77141 59740 77142 59804
rect 77206 59740 77207 59804
rect 77141 59739 77207 59740
rect 76054 59470 76116 59530
rect 78232 59530 78292 60106
rect 79592 59530 79652 60106
rect 80544 59530 80604 60106
rect 78232 59470 78322 59530
rect 59307 58444 59373 58445
rect 59307 58380 59308 58444
rect 59372 58380 59373 58444
rect 59307 58379 59373 58380
rect 59123 57220 59189 57221
rect 59123 57156 59124 57220
rect 59188 57156 59189 57220
rect 59123 57155 59189 57156
rect 58939 57084 59005 57085
rect 58939 57020 58940 57084
rect 59004 57020 59005 57084
rect 58939 57019 59005 57020
rect 57467 54772 57533 54773
rect 57467 54708 57468 54772
rect 57532 54708 57533 54772
rect 57467 54707 57533 54708
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 76054 57901 76114 59470
rect 76051 57900 76117 57901
rect 76051 57836 76052 57900
rect 76116 57836 76117 57900
rect 76051 57835 76117 57836
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 78262 57901 78322 59470
rect 79550 59470 79652 59530
rect 80470 59470 80604 59530
rect 81768 59530 81828 60106
rect 83128 59805 83188 60106
rect 83125 59804 83191 59805
rect 83125 59740 83126 59804
rect 83190 59740 83191 59804
rect 83125 59739 83191 59740
rect 84216 59530 84276 60106
rect 85440 59530 85500 60106
rect 81768 59470 82002 59530
rect 79550 57901 79610 59470
rect 80470 57901 80530 59470
rect 78259 57900 78325 57901
rect 78259 57836 78260 57900
rect 78324 57836 78325 57900
rect 78259 57835 78325 57836
rect 79547 57900 79613 57901
rect 79547 57836 79548 57900
rect 79612 57836 79613 57900
rect 79547 57835 79613 57836
rect 80467 57900 80533 57901
rect 80467 57836 80468 57900
rect 80532 57836 80533 57900
rect 80467 57835 80533 57836
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81942 57901 82002 59470
rect 83966 59470 84276 59530
rect 85438 59470 85500 59530
rect 86528 59530 86588 60106
rect 87616 59530 87676 60106
rect 88296 59530 88356 60106
rect 88704 59530 88764 60106
rect 90064 59530 90124 60106
rect 86528 59470 86602 59530
rect 87616 59470 87706 59530
rect 88296 59470 88442 59530
rect 88704 59470 88810 59530
rect 83966 58037 84026 59470
rect 85438 58173 85498 59470
rect 85435 58172 85501 58173
rect 85435 58108 85436 58172
rect 85500 58108 85501 58172
rect 85435 58107 85501 58108
rect 83963 58036 84029 58037
rect 83963 57972 83964 58036
rect 84028 57972 84029 58036
rect 83963 57971 84029 57972
rect 81939 57900 82005 57901
rect 81939 57836 81940 57900
rect 82004 57836 82005 57900
rect 81939 57835 82005 57836
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 86542 57901 86602 59470
rect 87646 57901 87706 59470
rect 88382 57901 88442 59470
rect 88750 57901 88810 59470
rect 90038 59470 90124 59530
rect 90744 59530 90804 60106
rect 91288 59530 91348 60106
rect 92376 59530 92436 60106
rect 93464 59530 93524 60106
rect 90744 59470 90834 59530
rect 91288 59470 91386 59530
rect 90038 57901 90098 59470
rect 90774 57901 90834 59470
rect 91326 57901 91386 59470
rect 92246 59470 92436 59530
rect 93350 59470 93524 59530
rect 93600 59530 93660 60106
rect 94552 59669 94612 60106
rect 94549 59668 94615 59669
rect 94549 59604 94550 59668
rect 94614 59604 94615 59668
rect 95912 59666 95972 60106
rect 95912 59606 95986 59666
rect 94549 59603 94615 59604
rect 93600 59470 93778 59530
rect 92246 58173 92306 59470
rect 92243 58172 92309 58173
rect 92243 58108 92244 58172
rect 92308 58108 92309 58172
rect 92243 58107 92309 58108
rect 86539 57900 86605 57901
rect 86539 57836 86540 57900
rect 86604 57836 86605 57900
rect 86539 57835 86605 57836
rect 87643 57900 87709 57901
rect 87643 57836 87644 57900
rect 87708 57836 87709 57900
rect 87643 57835 87709 57836
rect 88379 57900 88445 57901
rect 88379 57836 88380 57900
rect 88444 57836 88445 57900
rect 88379 57835 88445 57836
rect 88747 57900 88813 57901
rect 88747 57836 88748 57900
rect 88812 57836 88813 57900
rect 88747 57835 88813 57836
rect 90035 57900 90101 57901
rect 90035 57836 90036 57900
rect 90100 57836 90101 57900
rect 90035 57835 90101 57836
rect 90771 57900 90837 57901
rect 90771 57836 90772 57900
rect 90836 57836 90837 57900
rect 90771 57835 90837 57836
rect 91323 57900 91389 57901
rect 91323 57836 91324 57900
rect 91388 57836 91389 57900
rect 91323 57835 91389 57836
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 93350 57901 93410 59470
rect 93347 57900 93413 57901
rect 93347 57836 93348 57900
rect 93412 57836 93413 57900
rect 93347 57835 93413 57836
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 93718 57085 93778 59470
rect 95926 59397 95986 59606
rect 96048 59530 96108 60106
rect 97000 59530 97060 60106
rect 98088 59666 98148 60106
rect 98088 59606 98194 59666
rect 96048 59470 96354 59530
rect 97000 59470 97090 59530
rect 95923 59396 95989 59397
rect 95923 59332 95924 59396
rect 95988 59332 95989 59396
rect 95923 59331 95989 59332
rect 93715 57084 93781 57085
rect 93715 57020 93716 57084
rect 93780 57020 93781 57084
rect 93715 57019 93781 57020
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 96294 57221 96354 59470
rect 97030 57357 97090 59470
rect 98134 59397 98194 59606
rect 98496 59530 98556 60106
rect 99448 59805 99508 60106
rect 99445 59804 99511 59805
rect 99445 59740 99446 59804
rect 99510 59740 99511 59804
rect 99445 59739 99511 59740
rect 100672 59666 100732 60106
rect 100672 59606 100770 59666
rect 98496 59470 98562 59530
rect 98131 59396 98197 59397
rect 98131 59332 98132 59396
rect 98196 59332 98197 59396
rect 98131 59331 98197 59332
rect 98502 57629 98562 59470
rect 100710 59397 100770 59606
rect 101080 59530 101140 60106
rect 101078 59470 101140 59530
rect 101760 59530 101820 60106
rect 102848 59669 102908 60106
rect 102845 59668 102911 59669
rect 102845 59604 102846 59668
rect 102910 59604 102911 59668
rect 102845 59603 102911 59604
rect 103528 59530 103588 60106
rect 103936 59666 103996 60106
rect 103838 59606 103996 59666
rect 101760 59470 101874 59530
rect 103528 59470 103714 59530
rect 100707 59396 100773 59397
rect 100707 59332 100708 59396
rect 100772 59332 100773 59396
rect 100707 59331 100773 59332
rect 101078 58445 101138 59470
rect 101814 59397 101874 59470
rect 101811 59396 101877 59397
rect 101811 59332 101812 59396
rect 101876 59332 101877 59396
rect 101811 59331 101877 59332
rect 101075 58444 101141 58445
rect 101075 58380 101076 58444
rect 101140 58380 101141 58444
rect 101075 58379 101141 58380
rect 98499 57628 98565 57629
rect 98499 57564 98500 57628
rect 98564 57564 98565 57628
rect 98499 57563 98565 57564
rect 97027 57356 97093 57357
rect 97027 57292 97028 57356
rect 97092 57292 97093 57356
rect 97027 57291 97093 57292
rect 96291 57220 96357 57221
rect 96291 57156 96292 57220
rect 96356 57156 96357 57220
rect 96291 57155 96357 57156
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 103654 57490 103714 59470
rect 103838 57901 103898 59606
rect 105296 59530 105356 60106
rect 105976 59669 106036 60106
rect 105973 59668 106039 59669
rect 105973 59604 105974 59668
rect 106038 59604 106039 59668
rect 105973 59603 106039 59604
rect 106384 59530 106444 60106
rect 107608 59666 107668 60106
rect 107518 59606 107668 59666
rect 105296 59470 105370 59530
rect 106384 59470 106474 59530
rect 105310 57901 105370 59470
rect 106414 57901 106474 59470
rect 107518 57901 107578 59606
rect 108288 59530 108348 60106
rect 108696 59666 108756 60106
rect 108254 59470 108348 59530
rect 108622 59606 108756 59666
rect 108254 58717 108314 59470
rect 108251 58716 108317 58717
rect 108251 58652 108252 58716
rect 108316 58652 108317 58716
rect 108251 58651 108317 58652
rect 108622 57901 108682 59606
rect 109784 59530 109844 60106
rect 109542 59470 109844 59530
rect 111008 59530 111068 60106
rect 111144 59530 111204 60106
rect 112232 59666 112292 60106
rect 113320 59669 113380 60106
rect 113592 59805 113652 60106
rect 113589 59804 113655 59805
rect 113589 59740 113590 59804
rect 113654 59740 113655 59804
rect 113589 59739 113655 59740
rect 112118 59606 112292 59666
rect 113317 59668 113383 59669
rect 111008 59470 111074 59530
rect 111144 59470 111258 59530
rect 109542 57901 109602 59470
rect 111014 58581 111074 59470
rect 111011 58580 111077 58581
rect 111011 58516 111012 58580
rect 111076 58516 111077 58580
rect 111011 58515 111077 58516
rect 103835 57900 103901 57901
rect 103835 57836 103836 57900
rect 103900 57836 103901 57900
rect 103835 57835 103901 57836
rect 105307 57900 105373 57901
rect 105307 57836 105308 57900
rect 105372 57836 105373 57900
rect 105307 57835 105373 57836
rect 106411 57900 106477 57901
rect 106411 57836 106412 57900
rect 106476 57836 106477 57900
rect 106411 57835 106477 57836
rect 107515 57900 107581 57901
rect 107515 57836 107516 57900
rect 107580 57836 107581 57900
rect 107515 57835 107581 57836
rect 108619 57900 108685 57901
rect 108619 57836 108620 57900
rect 108684 57836 108685 57900
rect 108619 57835 108685 57836
rect 109539 57900 109605 57901
rect 109539 57836 109540 57900
rect 109604 57836 109605 57900
rect 109539 57835 109605 57836
rect 103835 57492 103901 57493
rect 103835 57490 103836 57492
rect 103654 57430 103836 57490
rect 103835 57428 103836 57430
rect 103900 57428 103901 57492
rect 103835 57427 103901 57428
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 111198 57901 111258 59470
rect 111195 57900 111261 57901
rect 111195 57836 111196 57900
rect 111260 57836 111261 57900
rect 111195 57835 111261 57836
rect 112118 57629 112178 59606
rect 113317 59604 113318 59668
rect 113382 59604 113383 59668
rect 113317 59603 113383 59604
rect 114408 59530 114468 60106
rect 114326 59470 114468 59530
rect 115768 59530 115828 60106
rect 116040 59530 116100 60106
rect 116992 59669 117052 60106
rect 116989 59668 117055 59669
rect 116989 59604 116990 59668
rect 117054 59604 117055 59668
rect 116989 59603 117055 59604
rect 118080 59530 118140 60106
rect 118488 59530 118548 60106
rect 119168 59530 119228 60106
rect 120936 59805 120996 60106
rect 120933 59804 120999 59805
rect 120933 59740 120934 59804
rect 120998 59740 120999 59804
rect 120933 59739 120999 59740
rect 115768 59470 115858 59530
rect 112115 57628 112181 57629
rect 112115 57564 112116 57628
rect 112180 57564 112181 57628
rect 112115 57563 112181 57564
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 114326 57629 114386 59470
rect 115798 57901 115858 59470
rect 115982 59470 116100 59530
rect 118006 59470 118140 59530
rect 118374 59470 118548 59530
rect 119110 59470 119228 59530
rect 123520 59530 123580 60106
rect 125968 59530 126028 60106
rect 123520 59470 123586 59530
rect 115795 57900 115861 57901
rect 115795 57836 115796 57900
rect 115860 57836 115861 57900
rect 115795 57835 115861 57836
rect 115982 57629 116042 59470
rect 114323 57628 114389 57629
rect 114323 57564 114324 57628
rect 114388 57564 114389 57628
rect 114323 57563 114389 57564
rect 115979 57628 116045 57629
rect 115979 57564 115980 57628
rect 116044 57564 116045 57628
rect 115979 57563 116045 57564
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 118006 57765 118066 59470
rect 118003 57764 118069 57765
rect 118003 57700 118004 57764
rect 118068 57700 118069 57764
rect 118003 57699 118069 57700
rect 118374 56677 118434 59470
rect 119110 57629 119170 59470
rect 119107 57628 119173 57629
rect 119107 57564 119108 57628
rect 119172 57564 119173 57628
rect 119107 57563 119173 57564
rect 118371 56676 118437 56677
rect 118371 56612 118372 56676
rect 118436 56612 118437 56676
rect 118371 56611 118437 56612
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 123526 57901 123586 59470
rect 125918 59470 126028 59530
rect 128280 59530 128340 60106
rect 131000 59530 131060 60106
rect 128280 59470 128370 59530
rect 125918 57901 125978 59470
rect 128310 58173 128370 59470
rect 130886 59470 131060 59530
rect 133448 59530 133508 60106
rect 135896 59530 135956 60106
rect 138480 59530 138540 60106
rect 140928 59530 140988 60106
rect 133448 59470 133522 59530
rect 128307 58172 128373 58173
rect 128307 58108 128308 58172
rect 128372 58108 128373 58172
rect 128307 58107 128373 58108
rect 123523 57900 123589 57901
rect 123523 57836 123524 57900
rect 123588 57836 123589 57900
rect 123523 57835 123589 57836
rect 125915 57900 125981 57901
rect 125915 57836 125916 57900
rect 125980 57836 125981 57900
rect 125915 57835 125981 57836
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 130886 57901 130946 59470
rect 130883 57900 130949 57901
rect 130883 57836 130884 57900
rect 130948 57836 130949 57900
rect 130883 57835 130949 57836
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 133462 57901 133522 59470
rect 135854 59470 135956 59530
rect 138430 59470 138540 59530
rect 140822 59470 140988 59530
rect 143512 59530 143572 60106
rect 145960 59530 146020 60106
rect 143512 59470 143642 59530
rect 135854 58853 135914 59470
rect 138430 58989 138490 59470
rect 140822 59125 140882 59470
rect 143582 59261 143642 59470
rect 145606 59470 146020 59530
rect 148544 59530 148604 60106
rect 150992 59530 151052 60106
rect 153440 59530 153500 60106
rect 148544 59470 148610 59530
rect 143579 59260 143645 59261
rect 143579 59196 143580 59260
rect 143644 59196 143645 59260
rect 143579 59195 143645 59196
rect 140819 59124 140885 59125
rect 140819 59060 140820 59124
rect 140884 59060 140885 59124
rect 140819 59059 140885 59060
rect 138427 58988 138493 58989
rect 138427 58924 138428 58988
rect 138492 58924 138493 58988
rect 138427 58923 138493 58924
rect 135851 58852 135917 58853
rect 135851 58788 135852 58852
rect 135916 58788 135917 58852
rect 135851 58787 135917 58788
rect 133459 57900 133525 57901
rect 133459 57836 133460 57900
rect 133524 57836 133525 57900
rect 133459 57835 133525 57836
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 145606 57901 145666 59470
rect 148550 59261 148610 59470
rect 150942 59470 151052 59530
rect 153334 59470 153500 59530
rect 155888 59530 155948 60106
rect 158472 59530 158532 60106
rect 160920 59530 160980 60106
rect 163368 59530 163428 60106
rect 165952 59530 166012 60106
rect 183224 59530 183284 60106
rect 155888 59470 155970 59530
rect 158472 59470 158546 59530
rect 150942 59261 151002 59470
rect 148547 59260 148613 59261
rect 148547 59196 148548 59260
rect 148612 59196 148613 59260
rect 148547 59195 148613 59196
rect 150939 59260 151005 59261
rect 150939 59196 150940 59260
rect 151004 59196 151005 59260
rect 150939 59195 151005 59196
rect 153334 58173 153394 59470
rect 153331 58172 153397 58173
rect 153331 58108 153332 58172
rect 153396 58108 153397 58172
rect 153331 58107 153397 58108
rect 145603 57900 145669 57901
rect 145603 57836 145604 57900
rect 145668 57836 145669 57900
rect 145603 57835 145669 57836
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 155910 57629 155970 59470
rect 155907 57628 155973 57629
rect 155907 57564 155908 57628
rect 155972 57564 155973 57628
rect 155907 57563 155973 57564
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 158486 56405 158546 59470
rect 160878 59470 160980 59530
rect 163270 59470 163428 59530
rect 165846 59470 166012 59530
rect 183142 59470 183284 59530
rect 183360 59530 183420 60106
rect 183360 59470 183570 59530
rect 160878 57629 160938 59470
rect 160875 57628 160941 57629
rect 160875 57564 160876 57628
rect 160940 57564 160941 57628
rect 160875 57563 160941 57564
rect 163270 56677 163330 59470
rect 163794 57454 164414 58000
rect 165846 57629 165906 59470
rect 165843 57628 165909 57629
rect 165843 57564 165844 57628
rect 165908 57564 165909 57628
rect 165843 57563 165909 57564
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163267 56676 163333 56677
rect 163267 56612 163268 56676
rect 163332 56612 163333 56676
rect 163267 56611 163333 56612
rect 158483 56404 158549 56405
rect 158483 56340 158484 56404
rect 158548 56340 158549 56404
rect 158483 56339 158549 56340
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 183142 57901 183202 59470
rect 183139 57900 183205 57901
rect 183139 57836 183140 57900
rect 183204 57836 183205 57900
rect 183139 57835 183205 57836
rect 183510 57765 183570 59470
rect 197862 59397 197922 478347
rect 198046 163573 198106 478619
rect 201355 478548 201421 478549
rect 201355 478484 201356 478548
rect 201420 478484 201421 478548
rect 201355 478483 201421 478484
rect 200619 478140 200685 478141
rect 200619 478076 200620 478140
rect 200684 478076 200685 478140
rect 200619 478075 200685 478076
rect 198227 478004 198293 478005
rect 198227 477940 198228 478004
rect 198292 477940 198293 478004
rect 198227 477939 198293 477940
rect 198230 375325 198290 477939
rect 198595 477868 198661 477869
rect 198595 477804 198596 477868
rect 198660 477804 198661 477868
rect 198595 477803 198661 477804
rect 198227 375324 198293 375325
rect 198227 375260 198228 375324
rect 198292 375260 198293 375324
rect 198227 375259 198293 375260
rect 198043 163572 198109 163573
rect 198043 163508 198044 163572
rect 198108 163508 198109 163572
rect 198043 163507 198109 163508
rect 197859 59396 197925 59397
rect 197859 59332 197860 59396
rect 197924 59332 197925 59396
rect 197859 59331 197925 59332
rect 198598 59125 198658 477803
rect 199331 477732 199397 477733
rect 199331 477668 199332 477732
rect 199396 477668 199397 477732
rect 199331 477667 199397 477668
rect 199147 471204 199213 471205
rect 199147 471140 199148 471204
rect 199212 471140 199213 471204
rect 199147 471139 199213 471140
rect 198963 462908 199029 462909
rect 198963 462844 198964 462908
rect 199028 462844 199029 462908
rect 198963 462843 199029 462844
rect 198779 460052 198845 460053
rect 198779 459988 198780 460052
rect 198844 459988 198845 460052
rect 198779 459987 198845 459988
rect 198782 162621 198842 459987
rect 198966 267613 199026 462843
rect 199150 392733 199210 471139
rect 199147 392732 199213 392733
rect 199147 392668 199148 392732
rect 199212 392668 199213 392732
rect 199147 392667 199213 392668
rect 199150 392053 199210 392667
rect 199147 392052 199213 392053
rect 199147 391988 199148 392052
rect 199212 391988 199213 392052
rect 199147 391987 199213 391988
rect 199334 268973 199394 477667
rect 199794 470514 200414 478000
rect 199794 470278 199826 470514
rect 200062 470278 200146 470514
rect 200382 470278 200414 470514
rect 199794 470194 200414 470278
rect 199794 469958 199826 470194
rect 200062 469958 200146 470194
rect 200382 469958 200414 470194
rect 199794 453454 200414 469958
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199515 392052 199581 392053
rect 199515 391988 199516 392052
rect 199580 391988 199581 392052
rect 199515 391987 199581 391988
rect 199518 358053 199578 391987
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 364394 200414 380898
rect 199794 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 200414 364394
rect 199794 364074 200414 364158
rect 199794 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 200414 364074
rect 199515 358052 199581 358053
rect 199515 357988 199516 358052
rect 199580 357988 199581 358052
rect 199515 357987 199581 357988
rect 199794 345454 200414 363838
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199331 268972 199397 268973
rect 199331 268908 199332 268972
rect 199396 268908 199397 268972
rect 199331 268907 199397 268908
rect 198963 267612 199029 267613
rect 198963 267548 198964 267612
rect 199028 267548 199029 267612
rect 198963 267547 199029 267548
rect 199794 256394 200414 272898
rect 199794 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 200414 256394
rect 199794 256074 200414 256158
rect 199794 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 200414 256074
rect 199794 237454 200414 255838
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 198779 162620 198845 162621
rect 198779 162556 198780 162620
rect 198844 162556 198845 162620
rect 198779 162555 198845 162556
rect 199794 148394 200414 164898
rect 199794 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 200414 148394
rect 199794 148074 200414 148158
rect 199794 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 200414 148074
rect 199794 129454 200414 147838
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 198595 59124 198661 59125
rect 198595 59060 198596 59124
rect 198660 59060 198661 59124
rect 198595 59059 198661 59060
rect 183507 57764 183573 57765
rect 183507 57700 183508 57764
rect 183572 57700 183573 57764
rect 183507 57699 183573 57700
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 92898
rect 200622 58445 200682 478075
rect 200987 477596 201053 477597
rect 200987 477532 200988 477596
rect 201052 477532 201053 477596
rect 200987 477531 201053 477532
rect 200803 461548 200869 461549
rect 200803 461484 200804 461548
rect 200868 461484 200869 461548
rect 200803 461483 200869 461484
rect 200806 161941 200866 461483
rect 200990 375325 201050 477531
rect 200987 375324 201053 375325
rect 200987 375260 200988 375324
rect 201052 375260 201053 375324
rect 200987 375259 201053 375260
rect 200803 161940 200869 161941
rect 200803 161876 200804 161940
rect 200868 161876 200869 161940
rect 200803 161875 200869 161876
rect 201358 58853 201418 478483
rect 202091 478276 202157 478277
rect 202091 478212 202092 478276
rect 202156 478212 202157 478276
rect 202091 478211 202157 478212
rect 201355 58852 201421 58853
rect 201355 58788 201356 58852
rect 201420 58788 201421 58852
rect 201355 58787 201421 58788
rect 202094 58581 202154 478211
rect 202275 471612 202341 471613
rect 202275 471548 202276 471612
rect 202340 471548 202341 471612
rect 202275 471547 202341 471548
rect 202091 58580 202157 58581
rect 202091 58516 202092 58580
rect 202156 58516 202157 58580
rect 202091 58515 202157 58516
rect 200619 58444 200685 58445
rect 200619 58380 200620 58444
rect 200684 58380 200685 58444
rect 200619 58379 200685 58380
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 202278 56677 202338 471547
rect 202462 164117 202522 478755
rect 211843 478684 211909 478685
rect 211843 478620 211844 478684
rect 211908 478620 211909 478684
rect 211843 478619 211909 478620
rect 206691 478548 206757 478549
rect 206691 478484 206692 478548
rect 206756 478484 206757 478548
rect 206691 478483 206757 478484
rect 202643 478412 202709 478413
rect 202643 478348 202644 478412
rect 202708 478348 202709 478412
rect 202643 478347 202709 478348
rect 202459 164116 202525 164117
rect 202459 164052 202460 164116
rect 202524 164052 202525 164116
rect 202459 164051 202525 164052
rect 202646 59261 202706 478347
rect 203514 474234 204134 478000
rect 206507 477732 206573 477733
rect 206507 477668 206508 477732
rect 206572 477668 206573 477732
rect 206507 477667 206573 477668
rect 204851 474332 204917 474333
rect 204851 474268 204852 474332
rect 204916 474268 204917 474332
rect 204851 474267 204917 474268
rect 203514 473998 203546 474234
rect 203782 473998 203866 474234
rect 204102 473998 204134 474234
rect 203514 473914 204134 473998
rect 203514 473678 203546 473914
rect 203782 473678 203866 473914
rect 204102 473678 204134 473914
rect 203195 467260 203261 467261
rect 203195 467196 203196 467260
rect 203260 467196 203261 467260
rect 203195 467195 203261 467196
rect 203011 463452 203077 463453
rect 203011 463388 203012 463452
rect 203076 463388 203077 463452
rect 203011 463387 203077 463388
rect 203014 163981 203074 463387
rect 203011 163980 203077 163981
rect 203011 163916 203012 163980
rect 203076 163916 203077 163980
rect 203011 163915 203077 163916
rect 203198 162485 203258 467195
rect 203514 457174 204134 473678
rect 204299 463180 204365 463181
rect 204299 463116 204300 463180
rect 204364 463116 204365 463180
rect 204299 463115 204365 463116
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 366234 204134 384618
rect 204302 375325 204362 463115
rect 204299 375324 204365 375325
rect 204299 375260 204300 375324
rect 204364 375260 204365 375324
rect 204299 375259 204365 375260
rect 203514 365998 203546 366234
rect 203782 365998 203866 366234
rect 204102 365998 204134 366234
rect 203514 365914 204134 365998
rect 203514 365678 203546 365914
rect 203782 365678 203866 365914
rect 204102 365678 204134 365914
rect 203514 349174 204134 365678
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 260114 204134 276618
rect 203514 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 204134 260114
rect 203514 259794 204134 259878
rect 203514 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 204134 259794
rect 203514 241174 204134 259558
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203195 162484 203261 162485
rect 203195 162420 203196 162484
rect 203260 162420 203261 162484
rect 203195 162419 203261 162420
rect 203514 152114 204134 168618
rect 203514 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 204134 152114
rect 203514 151794 204134 151878
rect 203514 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 204134 151794
rect 203514 133174 204134 151558
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 202643 59260 202709 59261
rect 202643 59196 202644 59260
rect 202708 59196 202709 59260
rect 202643 59195 202709 59196
rect 202275 56676 202341 56677
rect 202275 56612 202276 56676
rect 202340 56612 202341 56676
rect 202275 56611 202341 56612
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 60618
rect 204854 57629 204914 474267
rect 205035 474196 205101 474197
rect 205035 474132 205036 474196
rect 205100 474132 205101 474196
rect 205035 474131 205101 474132
rect 204851 57628 204917 57629
rect 204851 57564 204852 57628
rect 204916 57564 204917 57628
rect 204851 57563 204917 57564
rect 205038 57357 205098 474131
rect 206323 460868 206389 460869
rect 206323 460804 206324 460868
rect 206388 460804 206389 460868
rect 206323 460803 206389 460804
rect 205219 460460 205285 460461
rect 205219 460396 205220 460460
rect 205284 460396 205285 460460
rect 205219 460395 205285 460396
rect 205035 57356 205101 57357
rect 205035 57292 205036 57356
rect 205100 57292 205101 57356
rect 205035 57291 205101 57292
rect 205222 55181 205282 460395
rect 206139 460324 206205 460325
rect 206139 460260 206140 460324
rect 206204 460260 206205 460324
rect 206139 460259 206205 460260
rect 206142 68101 206202 460259
rect 206326 163845 206386 460803
rect 206510 374645 206570 477667
rect 206694 408645 206754 478483
rect 210739 478276 210805 478277
rect 210739 478212 210740 478276
rect 210804 478212 210805 478276
rect 210739 478211 210805 478212
rect 209635 478004 209701 478005
rect 207234 470078 207854 478000
rect 209635 477940 209636 478004
rect 209700 477940 209701 478004
rect 209635 477939 209701 477940
rect 208347 476780 208413 476781
rect 208347 476716 208348 476780
rect 208412 476716 208413 476780
rect 208347 476715 208413 476716
rect 207234 469842 207266 470078
rect 207502 469842 207586 470078
rect 207822 469842 207854 470078
rect 207234 469758 207854 469842
rect 207234 469522 207266 469758
rect 207502 469522 207586 469758
rect 207822 469522 207854 469758
rect 207059 467124 207125 467125
rect 207059 467060 207060 467124
rect 207124 467060 207125 467124
rect 207059 467059 207125 467060
rect 206691 408644 206757 408645
rect 206691 408580 206692 408644
rect 206756 408580 206757 408644
rect 206691 408579 206757 408580
rect 207062 382397 207122 467059
rect 207234 460894 207854 469522
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207979 459100 208045 459101
rect 207979 459036 207980 459100
rect 208044 459036 208045 459100
rect 207979 459035 208045 459036
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207059 382396 207125 382397
rect 207059 382332 207060 382396
rect 207124 382332 207125 382396
rect 207059 382331 207125 382332
rect 206507 374644 206573 374645
rect 206507 374580 206508 374644
rect 206572 374580 206573 374644
rect 206507 374579 206573 374580
rect 207234 369954 207854 388338
rect 207234 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 207854 369954
rect 207234 369634 207854 369718
rect 207234 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 207854 369634
rect 207234 352894 207854 369398
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 261954 207854 280338
rect 207234 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 207854 261954
rect 207234 261634 207854 261718
rect 207234 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 207854 261634
rect 207234 244894 207854 261398
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 206323 163844 206389 163845
rect 206323 163780 206324 163844
rect 206388 163780 206389 163844
rect 206323 163779 206389 163780
rect 207234 153954 207854 172338
rect 207982 163709 208042 459035
rect 208350 374645 208410 476715
rect 208899 472836 208965 472837
rect 208899 472772 208900 472836
rect 208964 472772 208965 472836
rect 208899 472771 208965 472772
rect 208347 374644 208413 374645
rect 208347 374580 208348 374644
rect 208412 374580 208413 374644
rect 208347 374579 208413 374580
rect 207979 163708 208045 163709
rect 207979 163644 207980 163708
rect 208044 163644 208045 163708
rect 207979 163643 208045 163644
rect 207234 153718 207266 153954
rect 207502 153718 207586 153954
rect 207822 153718 207854 153954
rect 207234 153634 207854 153718
rect 207234 153398 207266 153634
rect 207502 153398 207586 153634
rect 207822 153398 207854 153634
rect 207234 136894 207854 153398
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 206139 68100 206205 68101
rect 206139 68036 206140 68100
rect 206204 68036 206205 68100
rect 206139 68035 206205 68036
rect 207234 64894 207854 100338
rect 208902 70005 208962 472771
rect 208899 70004 208965 70005
rect 208899 69940 208900 70004
rect 208964 69940 208965 70004
rect 208899 69939 208965 69940
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 205219 55180 205285 55181
rect 205219 55116 205220 55180
rect 205284 55116 205285 55180
rect 205219 55115 205285 55116
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 64338
rect 209638 58717 209698 477939
rect 209819 469980 209885 469981
rect 209819 469916 209820 469980
rect 209884 469916 209885 469980
rect 209819 469915 209885 469916
rect 209822 374645 209882 469915
rect 210371 460732 210437 460733
rect 210371 460668 210372 460732
rect 210436 460668 210437 460732
rect 210371 460667 210437 460668
rect 209819 374644 209885 374645
rect 209819 374580 209820 374644
rect 209884 374580 209885 374644
rect 209819 374579 209885 374580
rect 210374 164253 210434 460667
rect 210371 164252 210437 164253
rect 210371 164188 210372 164252
rect 210436 164188 210437 164252
rect 210371 164187 210437 164188
rect 210742 58989 210802 478211
rect 210954 464614 211574 478000
rect 211659 475692 211725 475693
rect 211659 475628 211660 475692
rect 211724 475628 211725 475692
rect 211659 475627 211725 475628
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 265674 211574 284058
rect 210954 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 211574 265674
rect 210954 265354 211574 265438
rect 210954 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 211574 265354
rect 210954 248614 211574 265118
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 157674 211574 176058
rect 210954 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 211574 157674
rect 210954 157354 211574 157438
rect 210954 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 211574 157354
rect 210954 140614 211574 157118
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210739 58988 210805 58989
rect 210739 58924 210740 58988
rect 210804 58924 210805 58988
rect 210739 58923 210805 58924
rect 209635 58716 209701 58717
rect 209635 58652 209636 58716
rect 209700 58652 209701 58716
rect 209635 58651 209701 58652
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 68058
rect 211662 57765 211722 475627
rect 211846 270469 211906 478619
rect 219203 478276 219269 478277
rect 219203 478212 219204 478276
rect 219268 478212 219269 478276
rect 219203 478211 219269 478212
rect 216995 477596 217061 477597
rect 216995 477532 216996 477596
rect 217060 477532 217061 477596
rect 216995 477531 217061 477532
rect 217363 477596 217429 477597
rect 217363 477532 217364 477596
rect 217428 477532 217429 477596
rect 217363 477531 217429 477532
rect 217547 477596 217613 477597
rect 217547 477532 217548 477596
rect 217612 477532 217613 477596
rect 217547 477531 217613 477532
rect 214419 475556 214485 475557
rect 214419 475492 214420 475556
rect 214484 475492 214485 475556
rect 214419 475491 214485 475492
rect 212763 469844 212829 469845
rect 212763 469780 212764 469844
rect 212828 469780 212829 469844
rect 212763 469779 212829 469780
rect 212579 468620 212645 468621
rect 212579 468556 212580 468620
rect 212644 468556 212645 468620
rect 212579 468555 212645 468556
rect 211843 270468 211909 270469
rect 211843 270404 211844 270468
rect 211908 270404 211909 270468
rect 211843 270403 211909 270404
rect 212582 269109 212642 468555
rect 212766 369205 212826 469779
rect 213131 460596 213197 460597
rect 213131 460532 213132 460596
rect 213196 460532 213197 460596
rect 213131 460531 213197 460532
rect 212763 369204 212829 369205
rect 212763 369140 212764 369204
rect 212828 369140 212829 369204
rect 212763 369139 212829 369140
rect 212579 269108 212645 269109
rect 212579 269044 212580 269108
rect 212644 269044 212645 269108
rect 212579 269043 212645 269044
rect 213134 164389 213194 460531
rect 213131 164388 213197 164389
rect 213131 164324 213132 164388
rect 213196 164324 213197 164388
rect 213131 164323 213197 164324
rect 211659 57764 211725 57765
rect 211659 57700 211660 57764
rect 211724 57700 211725 57764
rect 211659 57699 211725 57700
rect 214422 57493 214482 475491
rect 214603 475420 214669 475421
rect 214603 475356 214604 475420
rect 214668 475356 214669 475420
rect 214603 475355 214669 475356
rect 214419 57492 214485 57493
rect 214419 57428 214420 57492
rect 214484 57428 214485 57492
rect 214419 57427 214485 57428
rect 214606 57085 214666 475355
rect 215339 474060 215405 474061
rect 215339 473996 215340 474060
rect 215404 473996 215405 474060
rect 215339 473995 215405 473996
rect 214787 472700 214853 472701
rect 214787 472636 214788 472700
rect 214852 472636 214853 472700
rect 214787 472635 214853 472636
rect 214790 162621 214850 472635
rect 214971 471476 215037 471477
rect 214971 471412 214972 471476
rect 215036 471412 215037 471476
rect 214971 471411 215037 471412
rect 214787 162620 214853 162621
rect 214787 162556 214788 162620
rect 214852 162556 214853 162620
rect 214787 162555 214853 162556
rect 214974 162349 215034 471411
rect 215342 251157 215402 473995
rect 215891 471340 215957 471341
rect 215891 471276 215892 471340
rect 215956 471276 215957 471340
rect 215891 471275 215957 471276
rect 215523 460188 215589 460189
rect 215523 460124 215524 460188
rect 215588 460124 215589 460188
rect 215523 460123 215589 460124
rect 215526 369205 215586 460123
rect 215523 369204 215589 369205
rect 215523 369140 215524 369204
rect 215588 369140 215589 369204
rect 215523 369139 215589 369140
rect 215339 251156 215405 251157
rect 215339 251092 215340 251156
rect 215404 251092 215405 251156
rect 215339 251091 215405 251092
rect 214971 162348 215037 162349
rect 214971 162284 214972 162348
rect 215036 162284 215037 162348
rect 214971 162283 215037 162284
rect 215894 57221 215954 471275
rect 216998 372741 217058 477531
rect 217179 466308 217245 466309
rect 217179 466244 217180 466308
rect 217244 466244 217245 466308
rect 217179 466243 217245 466244
rect 216995 372740 217061 372741
rect 216995 372676 216996 372740
rect 217060 372676 217061 372740
rect 216995 372675 217061 372676
rect 216998 371109 217058 372675
rect 216995 371108 217061 371109
rect 216995 371044 216996 371108
rect 217060 371044 217061 371108
rect 216995 371043 217061 371044
rect 216627 270604 216693 270605
rect 216627 270540 216628 270604
rect 216692 270540 216693 270604
rect 216627 270539 216693 270540
rect 216630 269789 216690 270539
rect 216627 269788 216693 269789
rect 216627 269724 216628 269788
rect 216692 269724 216693 269788
rect 216627 269723 216693 269724
rect 217182 269109 217242 466243
rect 217366 368389 217426 477531
rect 217550 371653 217610 477531
rect 217794 471454 218414 478000
rect 218835 472564 218901 472565
rect 218835 472500 218836 472564
rect 218900 472500 218901 472564
rect 218835 472499 218901 472500
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 460308 218414 470898
rect 218651 459780 218717 459781
rect 218651 459716 218652 459780
rect 218716 459716 218717 459780
rect 218651 459715 218717 459716
rect 217547 371652 217613 371653
rect 217547 371588 217548 371652
rect 217612 371588 217613 371652
rect 217547 371587 217613 371588
rect 217363 368388 217429 368389
rect 217363 368324 217364 368388
rect 217428 368324 217429 368388
rect 217363 368323 217429 368324
rect 217794 363454 218414 373000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 355308 218414 362898
rect 217363 353428 217429 353429
rect 217363 353364 217364 353428
rect 217428 353364 217429 353428
rect 217363 353363 217429 353364
rect 217366 270605 217426 353363
rect 217363 270604 217429 270605
rect 217363 270540 217364 270604
rect 217428 270540 217429 270604
rect 217363 270539 217429 270540
rect 217179 269108 217245 269109
rect 217179 269044 217180 269108
rect 217244 269044 217245 269108
rect 217179 269043 217245 269044
rect 217547 265980 217613 265981
rect 217547 265916 217548 265980
rect 217612 265916 217613 265980
rect 217547 265915 217613 265916
rect 217363 148340 217429 148341
rect 217363 148276 217364 148340
rect 217428 148276 217429 148340
rect 217363 148275 217429 148276
rect 217179 146436 217245 146437
rect 217179 146372 217180 146436
rect 217244 146372 217245 146436
rect 217179 146371 217245 146372
rect 215891 57220 215957 57221
rect 215891 57156 215892 57220
rect 215956 57156 215957 57220
rect 215891 57155 215957 57156
rect 214603 57084 214669 57085
rect 214603 57020 214604 57084
rect 214668 57020 214669 57084
rect 214603 57019 214669 57020
rect 217182 56405 217242 146371
rect 217179 56404 217245 56405
rect 217179 56340 217180 56404
rect 217244 56340 217245 56404
rect 217179 56339 217245 56340
rect 217366 55045 217426 148275
rect 217550 146029 217610 265915
rect 217794 255454 218414 268000
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 250308 218414 254898
rect 217794 147454 218414 163000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217547 146028 217613 146029
rect 217547 145964 217548 146028
rect 217612 145964 217613 146028
rect 217547 145963 217613 145964
rect 217363 55044 217429 55045
rect 217363 54980 217364 55044
rect 217428 54980 217429 55044
rect 217363 54979 217429 54980
rect 217550 54909 217610 145963
rect 217794 145308 218414 146898
rect 218654 60621 218714 459715
rect 218838 270469 218898 472499
rect 218835 270468 218901 270469
rect 218835 270404 218836 270468
rect 218900 270404 218901 270468
rect 218835 270403 218901 270404
rect 219206 60621 219266 478211
rect 219939 477596 220005 477597
rect 219939 477532 219940 477596
rect 220004 477532 220005 477596
rect 219939 477531 220005 477532
rect 218651 60620 218717 60621
rect 218651 60556 218652 60620
rect 218716 60556 218717 60620
rect 218651 60555 218717 60556
rect 219203 60620 219269 60621
rect 219203 60556 219204 60620
rect 219268 60556 219269 60620
rect 219203 60555 219269 60556
rect 217547 54908 217613 54909
rect 217547 54844 217548 54908
rect 217612 54844 217613 54908
rect 217547 54843 217613 54844
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 219942 56541 220002 477531
rect 221514 475174 222134 478000
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 460308 222134 474618
rect 225234 469138 225854 478000
rect 225234 468902 225266 469138
rect 225502 468902 225586 469138
rect 225822 468902 225854 469138
rect 225234 468818 225854 468902
rect 225234 468582 225266 468818
rect 225502 468582 225586 468818
rect 225822 468582 225854 468818
rect 225234 460308 225854 468582
rect 228954 465554 229574 478000
rect 228954 465318 228986 465554
rect 229222 465318 229306 465554
rect 229542 465318 229574 465554
rect 228954 465234 229574 465318
rect 228954 464998 228986 465234
rect 229222 464998 229306 465234
rect 229542 464998 229574 465234
rect 228954 460308 229574 464998
rect 235794 470514 236414 478000
rect 235794 470278 235826 470514
rect 236062 470278 236146 470514
rect 236382 470278 236414 470514
rect 235794 470194 236414 470278
rect 235794 469958 235826 470194
rect 236062 469958 236146 470194
rect 236382 469958 236414 470194
rect 235794 460308 236414 469958
rect 239514 474234 240134 478000
rect 239514 473998 239546 474234
rect 239782 473998 239866 474234
rect 240102 473998 240134 474234
rect 239514 473914 240134 473998
rect 239514 473678 239546 473914
rect 239782 473678 239866 473914
rect 240102 473678 240134 473914
rect 239514 460308 240134 473678
rect 243234 470078 243854 478000
rect 243234 469842 243266 470078
rect 243502 469842 243586 470078
rect 243822 469842 243854 470078
rect 243234 469758 243854 469842
rect 243234 469522 243266 469758
rect 243502 469522 243586 469758
rect 243822 469522 243854 469758
rect 243234 460308 243854 469522
rect 246954 464614 247574 478000
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 460308 247574 464058
rect 253794 471454 254414 478000
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 460308 254414 470898
rect 257514 475174 258134 478000
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 460308 258134 474618
rect 261234 469138 261854 478000
rect 261234 468902 261266 469138
rect 261502 468902 261586 469138
rect 261822 468902 261854 469138
rect 261234 468818 261854 468902
rect 261234 468582 261266 468818
rect 261502 468582 261586 468818
rect 261822 468582 261854 468818
rect 261234 460308 261854 468582
rect 264954 465554 265574 478000
rect 264954 465318 264986 465554
rect 265222 465318 265306 465554
rect 265542 465318 265574 465554
rect 264954 465234 265574 465318
rect 264954 464998 264986 465234
rect 265222 464998 265306 465234
rect 265542 464998 265574 465234
rect 264954 460308 265574 464998
rect 271794 470514 272414 478000
rect 271794 470278 271826 470514
rect 272062 470278 272146 470514
rect 272382 470278 272414 470514
rect 271794 470194 272414 470278
rect 271794 469958 271826 470194
rect 272062 469958 272146 470194
rect 272382 469958 272414 470194
rect 271794 460308 272414 469958
rect 275514 474234 276134 478000
rect 275514 473998 275546 474234
rect 275782 473998 275866 474234
rect 276102 473998 276134 474234
rect 275514 473914 276134 473998
rect 275514 473678 275546 473914
rect 275782 473678 275866 473914
rect 276102 473678 276134 473914
rect 275514 460308 276134 473678
rect 279234 470078 279854 478000
rect 279234 469842 279266 470078
rect 279502 469842 279586 470078
rect 279822 469842 279854 470078
rect 279234 469758 279854 469842
rect 279234 469522 279266 469758
rect 279502 469522 279586 469758
rect 279822 469522 279854 469758
rect 279234 460308 279854 469522
rect 282954 464614 283574 478000
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 460308 283574 464058
rect 289794 471454 290414 478000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 460308 290414 470898
rect 293514 475174 294134 478000
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 460308 294134 474618
rect 297234 469138 297854 478000
rect 297234 468902 297266 469138
rect 297502 468902 297586 469138
rect 297822 468902 297854 469138
rect 297234 468818 297854 468902
rect 297234 468582 297266 468818
rect 297502 468582 297586 468818
rect 297822 468582 297854 468818
rect 297234 460308 297854 468582
rect 300954 465554 301574 478000
rect 300954 465318 300986 465554
rect 301222 465318 301306 465554
rect 301542 465318 301574 465554
rect 300954 465234 301574 465318
rect 300954 464998 300986 465234
rect 301222 464998 301306 465234
rect 301542 464998 301574 465234
rect 300954 460308 301574 464998
rect 307794 460308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 460308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 633033 319574 644058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 633033 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 633033 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 633033 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 633033 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633033 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 633033 348134 636618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 633033 351854 640338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 633033 355574 644058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 633033 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 633033 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 633033 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 633033 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633033 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 633033 384134 636618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 633033 387854 640338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 633033 391574 644058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 633033 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 633033 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 633033 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 633033 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633033 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 633033 420134 636618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 633033 423854 640338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 633033 427574 644058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 324208 615454 324528 615486
rect 324208 615218 324250 615454
rect 324486 615218 324528 615454
rect 324208 615134 324528 615218
rect 324208 614898 324250 615134
rect 324486 614898 324528 615134
rect 324208 614866 324528 614898
rect 354928 615454 355248 615486
rect 354928 615218 354970 615454
rect 355206 615218 355248 615454
rect 354928 615134 355248 615218
rect 354928 614898 354970 615134
rect 355206 614898 355248 615134
rect 354928 614866 355248 614898
rect 385648 615454 385968 615486
rect 385648 615218 385690 615454
rect 385926 615218 385968 615454
rect 385648 615134 385968 615218
rect 385648 614898 385690 615134
rect 385926 614898 385968 615134
rect 385648 614866 385968 614898
rect 416368 615454 416688 615486
rect 416368 615218 416410 615454
rect 416646 615218 416688 615454
rect 416368 615134 416688 615218
rect 416368 614898 416410 615134
rect 416646 614898 416688 615134
rect 416368 614866 416688 614898
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 430619 597684 430685 597685
rect 430619 597620 430620 597684
rect 430684 597620 430685 597684
rect 430619 597619 430685 597620
rect 339568 597454 339888 597486
rect 339568 597218 339610 597454
rect 339846 597218 339888 597454
rect 339568 597134 339888 597218
rect 339568 596898 339610 597134
rect 339846 596898 339888 597134
rect 339568 596866 339888 596898
rect 370288 597454 370608 597486
rect 370288 597218 370330 597454
rect 370566 597218 370608 597454
rect 370288 597134 370608 597218
rect 370288 596898 370330 597134
rect 370566 596898 370608 597134
rect 370288 596866 370608 596898
rect 401008 597454 401328 597486
rect 401008 597218 401050 597454
rect 401286 597218 401328 597454
rect 401008 597134 401328 597218
rect 401008 596898 401050 597134
rect 401286 596898 401328 597134
rect 401008 596866 401328 596898
rect 324208 579454 324528 579486
rect 324208 579218 324250 579454
rect 324486 579218 324528 579454
rect 324208 579134 324528 579218
rect 324208 578898 324250 579134
rect 324486 578898 324528 579134
rect 324208 578866 324528 578898
rect 354928 579454 355248 579486
rect 354928 579218 354970 579454
rect 355206 579218 355248 579454
rect 354928 579134 355248 579218
rect 354928 578898 354970 579134
rect 355206 578898 355248 579134
rect 354928 578866 355248 578898
rect 385648 579454 385968 579486
rect 385648 579218 385690 579454
rect 385926 579218 385968 579454
rect 385648 579134 385968 579218
rect 385648 578898 385690 579134
rect 385926 578898 385968 579134
rect 385648 578866 385968 578898
rect 416368 579454 416688 579486
rect 416368 579218 416410 579454
rect 416646 579218 416688 579454
rect 416368 579134 416688 579218
rect 416368 578898 416410 579134
rect 416646 578898 416688 579134
rect 416368 578866 416688 578898
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 339568 561454 339888 561486
rect 339568 561218 339610 561454
rect 339846 561218 339888 561454
rect 339568 561134 339888 561218
rect 339568 560898 339610 561134
rect 339846 560898 339888 561134
rect 339568 560866 339888 560898
rect 370288 561454 370608 561486
rect 370288 561218 370330 561454
rect 370566 561218 370608 561454
rect 370288 561134 370608 561218
rect 370288 560898 370330 561134
rect 370566 560898 370608 561134
rect 370288 560866 370608 560898
rect 401008 561454 401328 561486
rect 401008 561218 401050 561454
rect 401286 561218 401328 561454
rect 401008 561134 401328 561218
rect 401008 560898 401050 561134
rect 401286 560898 401328 561134
rect 401008 560866 401328 560898
rect 324208 543454 324528 543486
rect 324208 543218 324250 543454
rect 324486 543218 324528 543454
rect 324208 543134 324528 543218
rect 324208 542898 324250 543134
rect 324486 542898 324528 543134
rect 324208 542866 324528 542898
rect 354928 543454 355248 543486
rect 354928 543218 354970 543454
rect 355206 543218 355248 543454
rect 354928 543134 355248 543218
rect 354928 542898 354970 543134
rect 355206 542898 355248 543134
rect 354928 542866 355248 542898
rect 385648 543454 385968 543486
rect 385648 543218 385690 543454
rect 385926 543218 385968 543454
rect 385648 543134 385968 543218
rect 385648 542898 385690 543134
rect 385926 542898 385968 543134
rect 385648 542866 385968 542898
rect 416368 543454 416688 543486
rect 416368 543218 416410 543454
rect 416646 543218 416688 543454
rect 416368 543134 416688 543218
rect 416368 542898 416410 543134
rect 416646 542898 416688 543134
rect 416368 542866 416688 542898
rect 320587 541108 320653 541109
rect 320587 541044 320588 541108
rect 320652 541044 320653 541108
rect 320587 541043 320653 541044
rect 320590 538230 320650 541043
rect 320590 538170 320834 538230
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 320774 518669 320834 538170
rect 339568 525454 339888 525486
rect 339568 525218 339610 525454
rect 339846 525218 339888 525454
rect 339568 525134 339888 525218
rect 339568 524898 339610 525134
rect 339846 524898 339888 525134
rect 339568 524866 339888 524898
rect 370288 525454 370608 525486
rect 370288 525218 370330 525454
rect 370566 525218 370608 525454
rect 370288 525134 370608 525218
rect 370288 524898 370330 525134
rect 370566 524898 370608 525134
rect 370288 524866 370608 524898
rect 401008 525454 401328 525486
rect 401008 525218 401050 525454
rect 401286 525218 401328 525454
rect 401008 525134 401328 525218
rect 401008 524898 401050 525134
rect 401286 524898 401328 525134
rect 401008 524866 401328 524898
rect 430622 518805 430682 597619
rect 430803 592244 430869 592245
rect 430803 592180 430804 592244
rect 430868 592180 430869 592244
rect 430803 592179 430869 592180
rect 430619 518804 430685 518805
rect 430619 518740 430620 518804
rect 430684 518740 430685 518804
rect 430619 518739 430685 518740
rect 320771 518668 320837 518669
rect 320771 518604 320772 518668
rect 320836 518604 320837 518668
rect 320771 518603 320837 518604
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460308 315854 496338
rect 318954 500614 319574 518000
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 460308 319574 464058
rect 325794 507454 326414 518000
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 460308 326414 470898
rect 329514 511174 330134 518000
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 460308 330134 474618
rect 333234 514894 333854 518000
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 460308 333854 478338
rect 336954 482614 337574 518000
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 460308 337574 482058
rect 343794 489454 344414 518000
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 338251 461004 338317 461005
rect 338251 460940 338252 461004
rect 338316 460950 338317 461004
rect 339723 461004 339789 461005
rect 338316 460940 338498 460950
rect 338251 460939 338498 460940
rect 339723 460940 339724 461004
rect 339788 460940 339789 461004
rect 339723 460939 339789 460940
rect 338254 460890 338498 460939
rect 338438 458690 338498 460890
rect 339726 458690 339786 460939
rect 343794 460308 344414 488898
rect 347514 493174 348134 518000
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 460308 348134 492618
rect 351234 496894 351854 518000
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350947 461004 351013 461005
rect 350947 460940 350948 461004
rect 351012 460940 351013 461004
rect 350947 460939 351013 460940
rect 350950 458690 351010 460939
rect 351234 460308 351854 496338
rect 354954 500614 355574 518000
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 361794 507454 362414 518000
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 360699 485076 360765 485077
rect 360699 485012 360700 485076
rect 360764 485012 360765 485076
rect 360699 485011 360765 485012
rect 357939 478820 358005 478821
rect 357939 478756 357940 478820
rect 358004 478756 358005 478820
rect 357939 478755 358005 478756
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 460308 355574 464058
rect 338438 458630 338524 458690
rect 338464 458202 338524 458630
rect 339688 458630 339786 458690
rect 350840 458630 351010 458690
rect 339688 458202 339748 458630
rect 350840 458202 350900 458630
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 220952 399454 221300 399486
rect 220952 399218 221008 399454
rect 221244 399218 221300 399454
rect 220952 399134 221300 399218
rect 220952 398898 221008 399134
rect 221244 398898 221300 399134
rect 220952 398866 221300 398898
rect 355320 399454 355668 399486
rect 355320 399218 355376 399454
rect 355612 399218 355668 399454
rect 355320 399134 355668 399218
rect 355320 398898 355376 399134
rect 355612 398898 355668 399134
rect 355320 398866 355668 398898
rect 220272 381454 220620 381486
rect 220272 381218 220328 381454
rect 220564 381218 220620 381454
rect 220272 381134 220620 381218
rect 220272 380898 220328 381134
rect 220564 380898 220620 381134
rect 220272 380866 220620 380898
rect 356000 381454 356348 381486
rect 356000 381218 356056 381454
rect 356292 381218 356348 381454
rect 356000 381134 356348 381218
rect 356000 380898 356056 381134
rect 356292 380898 356348 381134
rect 356000 380866 356348 380898
rect 236056 374509 236116 375020
rect 236502 374990 237174 375050
rect 238158 374990 238262 375050
rect 239262 374990 239622 375050
rect 240366 374990 240574 375050
rect 241654 374990 241798 375050
rect 242942 374990 243158 375050
rect 236053 374508 236119 374509
rect 236053 374444 236054 374508
rect 236118 374444 236119 374508
rect 236053 374443 236119 374444
rect 236502 373421 236562 374990
rect 236499 373420 236565 373421
rect 236499 373356 236500 373420
rect 236564 373356 236565 373420
rect 236499 373355 236565 373356
rect 221514 367174 222134 373000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 355308 222134 366618
rect 225234 370894 225854 373000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 355308 225854 370338
rect 228954 357554 229574 373000
rect 228954 357318 228986 357554
rect 229222 357318 229306 357554
rect 229542 357318 229574 357554
rect 228954 357234 229574 357318
rect 228954 356998 228986 357234
rect 229222 356998 229306 357234
rect 229542 356998 229574 357234
rect 228954 355308 229574 356998
rect 235794 364394 236414 373000
rect 238158 372605 238218 374990
rect 239262 372605 239322 374990
rect 238155 372604 238221 372605
rect 238155 372540 238156 372604
rect 238220 372540 238221 372604
rect 238155 372539 238221 372540
rect 239259 372604 239325 372605
rect 239259 372540 239260 372604
rect 239324 372540 239325 372604
rect 239259 372539 239325 372540
rect 235794 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 236414 364394
rect 235794 364074 236414 364158
rect 235794 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 236414 364074
rect 235794 355308 236414 363838
rect 239514 366234 240134 373000
rect 240366 372605 240426 374990
rect 241654 372605 241714 374990
rect 242942 373421 243002 374990
rect 244230 374509 244290 375050
rect 244782 374990 245470 375050
rect 245886 374990 246558 375050
rect 247174 374990 247646 375050
rect 247910 374990 248326 375050
rect 248462 374990 248734 375050
rect 244227 374508 244293 374509
rect 244227 374444 244228 374508
rect 244292 374444 244293 374508
rect 244227 374443 244293 374444
rect 242939 373420 243005 373421
rect 242939 373356 242940 373420
rect 243004 373356 243005 373420
rect 242939 373355 243005 373356
rect 240363 372604 240429 372605
rect 240363 372540 240364 372604
rect 240428 372540 240429 372604
rect 240363 372539 240429 372540
rect 241651 372604 241717 372605
rect 241651 372540 241652 372604
rect 241716 372540 241717 372604
rect 241651 372539 241717 372540
rect 239514 365998 239546 366234
rect 239782 365998 239866 366234
rect 240102 365998 240134 366234
rect 239514 365914 240134 365998
rect 239514 365678 239546 365914
rect 239782 365678 239866 365914
rect 240102 365678 240134 365914
rect 239514 355308 240134 365678
rect 243234 369954 243854 373000
rect 244782 372605 244842 374990
rect 244779 372604 244845 372605
rect 244779 372540 244780 372604
rect 244844 372540 244845 372604
rect 244779 372539 244845 372540
rect 245886 371789 245946 374990
rect 247174 373149 247234 374990
rect 247171 373148 247237 373149
rect 247171 373084 247172 373148
rect 247236 373084 247237 373148
rect 247171 373083 247237 373084
rect 245883 371788 245949 371789
rect 245883 371724 245884 371788
rect 245948 371724 245949 371788
rect 245883 371723 245949 371724
rect 243234 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 243854 369954
rect 243234 369634 243854 369718
rect 243234 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 243854 369634
rect 243234 355308 243854 369398
rect 246954 356614 247574 373000
rect 247910 371381 247970 374990
rect 248462 372605 248522 374990
rect 250064 374509 250124 375020
rect 250744 374509 250804 375020
rect 251288 374509 251348 375020
rect 251774 374990 252406 375050
rect 252878 374990 253494 375050
rect 250061 374508 250127 374509
rect 250061 374444 250062 374508
rect 250126 374444 250127 374508
rect 250061 374443 250127 374444
rect 250741 374508 250807 374509
rect 250741 374444 250742 374508
rect 250806 374444 250807 374508
rect 250741 374443 250807 374444
rect 251285 374508 251351 374509
rect 251285 374444 251286 374508
rect 251350 374444 251351 374508
rect 251285 374443 251351 374444
rect 251774 372605 251834 374990
rect 252878 372741 252938 374990
rect 252875 372740 252941 372741
rect 252875 372676 252876 372740
rect 252940 372676 252941 372740
rect 252875 372675 252941 372676
rect 248459 372604 248525 372605
rect 248459 372540 248460 372604
rect 248524 372540 248525 372604
rect 248459 372539 248525 372540
rect 251771 372604 251837 372605
rect 251771 372540 251772 372604
rect 251836 372540 251837 372604
rect 251771 372539 251837 372540
rect 253614 371381 253674 375050
rect 253982 374990 254582 375050
rect 255454 374990 255942 375050
rect 253982 373149 254042 374990
rect 255454 373557 255514 374990
rect 256048 374509 256108 375020
rect 256742 374990 257030 375050
rect 257846 374990 258118 375050
rect 258398 374990 258526 375050
rect 259478 374990 259562 375050
rect 256045 374508 256111 374509
rect 256045 374444 256046 374508
rect 256110 374444 256111 374508
rect 256045 374443 256111 374444
rect 256742 373557 256802 374990
rect 255451 373556 255517 373557
rect 255451 373492 255452 373556
rect 255516 373492 255517 373556
rect 255451 373491 255517 373492
rect 256739 373556 256805 373557
rect 256739 373492 256740 373556
rect 256804 373492 256805 373556
rect 256739 373491 256805 373492
rect 257846 373149 257906 374990
rect 253979 373148 254045 373149
rect 253979 373084 253980 373148
rect 254044 373084 254045 373148
rect 253979 373083 254045 373084
rect 257843 373148 257909 373149
rect 257843 373084 257844 373148
rect 257908 373084 257909 373148
rect 257843 373083 257909 373084
rect 247907 371380 247973 371381
rect 247907 371316 247908 371380
rect 247972 371316 247973 371380
rect 247907 371315 247973 371316
rect 253611 371380 253677 371381
rect 253611 371316 253612 371380
rect 253676 371316 253677 371380
rect 253611 371315 253677 371316
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 355308 247574 356058
rect 253794 363454 254414 373000
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 355308 254414 362898
rect 257514 367174 258134 373000
rect 258398 371381 258458 374990
rect 259502 372605 259562 374990
rect 260054 374990 260702 375050
rect 260974 374990 261110 375050
rect 261342 374990 261790 375050
rect 262262 374990 262878 375050
rect 260054 373421 260114 374990
rect 260051 373420 260117 373421
rect 260051 373356 260052 373420
rect 260116 373356 260117 373420
rect 260051 373355 260117 373356
rect 259499 372604 259565 372605
rect 259499 372540 259500 372604
rect 259564 372540 259565 372604
rect 259499 372539 259565 372540
rect 260974 371381 261034 374990
rect 261342 373149 261402 374990
rect 261339 373148 261405 373149
rect 261339 373084 261340 373148
rect 261404 373084 261405 373148
rect 261339 373083 261405 373084
rect 258395 371380 258461 371381
rect 258395 371316 258396 371380
rect 258460 371316 258461 371380
rect 258395 371315 258461 371316
rect 260971 371380 261037 371381
rect 260971 371316 260972 371380
rect 261036 371316 261037 371380
rect 260971 371315 261037 371316
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 355308 258134 366618
rect 261234 370894 261854 373000
rect 262262 372605 262322 374990
rect 262259 372604 262325 372605
rect 262259 372540 262260 372604
rect 262324 372540 262325 372604
rect 262259 372539 262325 372540
rect 263550 371381 263610 375050
rect 263734 374990 263966 375050
rect 265022 374990 265326 375050
rect 265758 374990 266006 375050
rect 266310 374990 266414 375050
rect 267046 374990 267638 375050
rect 267782 374990 268318 375050
rect 268518 374990 268726 375050
rect 269254 374990 269814 375050
rect 270910 374990 271038 375050
rect 263734 374373 263794 374990
rect 263731 374372 263797 374373
rect 263731 374308 263732 374372
rect 263796 374308 263797 374372
rect 263731 374307 263797 374308
rect 265022 373149 265082 374990
rect 265019 373148 265085 373149
rect 265019 373084 265020 373148
rect 265084 373084 265085 373148
rect 265019 373083 265085 373084
rect 263547 371380 263613 371381
rect 263547 371316 263548 371380
rect 263612 371316 263613 371380
rect 263547 371315 263613 371316
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 355308 261854 370338
rect 264954 357554 265574 373000
rect 265758 371381 265818 374990
rect 266310 372605 266370 374990
rect 266307 372604 266373 372605
rect 266307 372540 266308 372604
rect 266372 372540 266373 372604
rect 266307 372539 266373 372540
rect 267046 371381 267106 374990
rect 267782 371381 267842 374990
rect 268518 373829 268578 374990
rect 268515 373828 268581 373829
rect 268515 373764 268516 373828
rect 268580 373764 268581 373828
rect 268515 373763 268581 373764
rect 269254 373421 269314 374990
rect 269251 373420 269317 373421
rect 269251 373356 269252 373420
rect 269316 373356 269317 373420
rect 269251 373355 269317 373356
rect 270910 371381 270970 374990
rect 271144 374509 271204 375020
rect 272262 374990 272626 375050
rect 271141 374508 271207 374509
rect 271141 374444 271142 374508
rect 271206 374444 271207 374508
rect 271141 374443 271207 374444
rect 265755 371380 265821 371381
rect 265755 371316 265756 371380
rect 265820 371316 265821 371380
rect 265755 371315 265821 371316
rect 267043 371380 267109 371381
rect 267043 371316 267044 371380
rect 267108 371316 267109 371380
rect 267043 371315 267109 371316
rect 267779 371380 267845 371381
rect 267779 371316 267780 371380
rect 267844 371316 267845 371380
rect 267779 371315 267845 371316
rect 270907 371380 270973 371381
rect 270907 371316 270908 371380
rect 270972 371316 270973 371380
rect 270907 371315 270973 371316
rect 264954 357318 264986 357554
rect 265222 357318 265306 357554
rect 265542 357318 265574 357554
rect 264954 357234 265574 357318
rect 264954 356998 264986 357234
rect 265222 356998 265306 357234
rect 265542 356998 265574 357234
rect 264954 355308 265574 356998
rect 271794 364394 272414 373000
rect 272566 372605 272626 374990
rect 272563 372604 272629 372605
rect 272563 372540 272564 372604
rect 272628 372540 272629 372604
rect 272563 372539 272629 372540
rect 273302 372061 273362 375050
rect 273622 374990 273730 375050
rect 273299 372060 273365 372061
rect 273299 371996 273300 372060
rect 273364 371996 273365 372060
rect 273299 371995 273365 371996
rect 273670 371789 273730 374990
rect 273854 374990 274438 375050
rect 275142 374990 275798 375050
rect 276070 374990 276306 375050
rect 273667 371788 273733 371789
rect 273667 371724 273668 371788
rect 273732 371724 273733 371788
rect 273667 371723 273733 371724
rect 273854 371381 273914 374990
rect 275142 374101 275202 374990
rect 275139 374100 275205 374101
rect 275139 374036 275140 374100
rect 275204 374036 275205 374100
rect 275139 374035 275205 374036
rect 273851 371380 273917 371381
rect 273851 371316 273852 371380
rect 273916 371316 273917 371380
rect 273851 371315 273917 371316
rect 271794 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 272414 364394
rect 271794 364074 272414 364158
rect 271794 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 272414 364074
rect 271794 355308 272414 363838
rect 275514 366234 276134 373000
rect 276246 371381 276306 374990
rect 276982 372333 277042 375050
rect 277534 374990 278110 375050
rect 278270 374990 278518 375050
rect 278822 374990 279198 375050
rect 280294 374990 280966 375050
rect 283550 374990 283850 375050
rect 277534 372469 277594 374990
rect 277531 372468 277597 372469
rect 277531 372404 277532 372468
rect 277596 372404 277597 372468
rect 277531 372403 277597 372404
rect 276979 372332 277045 372333
rect 276979 372268 276980 372332
rect 277044 372268 277045 372332
rect 276979 372267 277045 372268
rect 278270 371517 278330 374990
rect 278822 373285 278882 374990
rect 278819 373284 278885 373285
rect 278819 373220 278820 373284
rect 278884 373220 278885 373284
rect 278819 373219 278885 373220
rect 278267 371516 278333 371517
rect 278267 371452 278268 371516
rect 278332 371452 278333 371516
rect 278267 371451 278333 371452
rect 276243 371380 276309 371381
rect 276243 371316 276244 371380
rect 276308 371316 276309 371380
rect 276243 371315 276309 371316
rect 275514 365998 275546 366234
rect 275782 365998 275866 366234
rect 276102 365998 276134 366234
rect 275514 365914 276134 365998
rect 275514 365678 275546 365914
rect 275782 365678 275866 365914
rect 276102 365678 276134 365914
rect 275514 355308 276134 365678
rect 279234 369954 279854 373000
rect 280294 371381 280354 374990
rect 280291 371380 280357 371381
rect 280291 371316 280292 371380
rect 280356 371316 280357 371380
rect 280291 371315 280357 371316
rect 279234 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 279854 369954
rect 279234 369634 279854 369718
rect 279234 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 279854 369634
rect 279234 355308 279854 369398
rect 282954 356614 283574 373000
rect 283790 371381 283850 374990
rect 285814 374990 285998 375050
rect 287654 374990 288310 375050
rect 290598 374990 291030 375050
rect 292806 374990 293478 375050
rect 295382 374990 295926 375050
rect 298142 374990 298510 375050
rect 285814 371381 285874 374990
rect 287654 371381 287714 374990
rect 283787 371380 283853 371381
rect 283787 371316 283788 371380
rect 283852 371316 283853 371380
rect 283787 371315 283853 371316
rect 285811 371380 285877 371381
rect 285811 371316 285812 371380
rect 285876 371316 285877 371380
rect 285811 371315 285877 371316
rect 287651 371380 287717 371381
rect 287651 371316 287652 371380
rect 287716 371316 287717 371380
rect 287651 371315 287717 371316
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 355308 283574 356058
rect 289794 363454 290414 373000
rect 290598 371381 290658 374990
rect 292806 371381 292866 374990
rect 290595 371380 290661 371381
rect 290595 371316 290596 371380
rect 290660 371316 290661 371380
rect 290595 371315 290661 371316
rect 292803 371380 292869 371381
rect 292803 371316 292804 371380
rect 292868 371316 292869 371380
rect 292803 371315 292869 371316
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 355308 290414 362898
rect 293514 367174 294134 373000
rect 295382 371381 295442 374990
rect 295379 371380 295445 371381
rect 295379 371316 295380 371380
rect 295444 371316 295445 371380
rect 295379 371315 295445 371316
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 355308 294134 366618
rect 297234 370894 297854 373000
rect 298142 371381 298202 374990
rect 300902 373149 300962 375050
rect 302926 374990 303542 375050
rect 305318 374990 305990 375050
rect 308574 374990 308690 375050
rect 300899 373148 300965 373149
rect 300899 373084 300900 373148
rect 300964 373084 300965 373148
rect 300899 373083 300965 373084
rect 298139 371380 298205 371381
rect 298139 371316 298140 371380
rect 298204 371316 298205 371380
rect 298139 371315 298205 371316
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 355308 297854 370338
rect 300954 357554 301574 373000
rect 302926 371381 302986 374990
rect 305318 372333 305378 374990
rect 305315 372332 305381 372333
rect 305315 372268 305316 372332
rect 305380 372268 305381 372332
rect 305315 372267 305381 372268
rect 302923 371380 302989 371381
rect 302923 371316 302924 371380
rect 302988 371316 302989 371380
rect 302923 371315 302989 371316
rect 300954 357318 300986 357554
rect 301222 357318 301306 357554
rect 301542 357318 301574 357554
rect 300954 357234 301574 357318
rect 300954 356998 300986 357234
rect 301222 356998 301306 357234
rect 301542 356998 301574 357234
rect 300954 355308 301574 356998
rect 307794 364394 308414 373000
rect 308630 371381 308690 374990
rect 310654 374990 311022 375050
rect 310654 372605 310714 374990
rect 310651 372604 310717 372605
rect 310651 372540 310652 372604
rect 310716 372540 310717 372604
rect 310651 372539 310717 372540
rect 308627 371380 308693 371381
rect 308627 371316 308628 371380
rect 308692 371316 308693 371380
rect 308627 371315 308693 371316
rect 307794 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 308414 364394
rect 307794 364074 308414 364158
rect 307794 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 308414 364074
rect 307794 355308 308414 363838
rect 311514 366234 312134 373000
rect 313414 372469 313474 375050
rect 315070 374990 315918 375050
rect 317830 374990 318502 375050
rect 315070 372605 315130 374990
rect 315067 372604 315133 372605
rect 315067 372540 315068 372604
rect 315132 372540 315133 372604
rect 315067 372539 315133 372540
rect 313411 372468 313477 372469
rect 313411 372404 313412 372468
rect 313476 372404 313477 372468
rect 313411 372403 313477 372404
rect 311514 365998 311546 366234
rect 311782 365998 311866 366234
rect 312102 365998 312134 366234
rect 311514 365914 312134 365998
rect 311514 365678 311546 365914
rect 311782 365678 311866 365914
rect 312102 365678 312134 365914
rect 311514 355308 312134 365678
rect 315234 369954 315854 373000
rect 317830 371789 317890 374990
rect 320920 374509 320980 375020
rect 322982 374990 323398 375050
rect 325982 374990 326722 375050
rect 320917 374508 320983 374509
rect 320917 374444 320918 374508
rect 320982 374444 320983 374508
rect 320917 374443 320983 374444
rect 317827 371788 317893 371789
rect 317827 371724 317828 371788
rect 317892 371724 317893 371788
rect 317827 371723 317893 371724
rect 315234 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 315854 369954
rect 315234 369634 315854 369718
rect 315234 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 315854 369634
rect 315234 355308 315854 369398
rect 318954 356614 319574 373000
rect 322982 372605 323042 374990
rect 322979 372604 323045 372605
rect 322979 372540 322980 372604
rect 323044 372540 323045 372604
rect 322979 372539 323045 372540
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 355308 319574 356058
rect 325794 363454 326414 373000
rect 326662 371381 326722 374990
rect 343038 374990 343254 375050
rect 343390 374990 343466 375050
rect 326659 371380 326725 371381
rect 326659 371316 326660 371380
rect 326724 371316 326725 371380
rect 326659 371315 326725 371316
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 355308 326414 362898
rect 329514 367174 330134 373000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 355308 330134 366618
rect 333234 370894 333854 373000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 355308 333854 370338
rect 336954 357554 337574 373000
rect 343038 371381 343098 374990
rect 343406 371381 343466 374990
rect 343035 371380 343101 371381
rect 343035 371316 343036 371380
rect 343100 371316 343101 371380
rect 343035 371315 343101 371316
rect 343403 371380 343469 371381
rect 343403 371316 343404 371380
rect 343468 371316 343469 371380
rect 343403 371315 343469 371316
rect 336954 357318 336986 357554
rect 337222 357318 337306 357554
rect 337542 357318 337574 357554
rect 336954 357234 337574 357318
rect 336954 356998 336986 357234
rect 337222 356998 337306 357234
rect 337542 356998 337574 357234
rect 336954 355308 337574 356998
rect 343794 364394 344414 373000
rect 343794 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 344414 364394
rect 343794 364074 344414 364158
rect 343794 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 344414 364074
rect 343794 355308 344414 363838
rect 347514 366234 348134 373000
rect 347514 365998 347546 366234
rect 347782 365998 347866 366234
rect 348102 365998 348134 366234
rect 347514 365914 348134 365998
rect 347514 365678 347546 365914
rect 347782 365678 347866 365914
rect 348102 365678 348134 365914
rect 347514 355308 348134 365678
rect 351234 369954 351854 373000
rect 351234 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 351854 369954
rect 351234 369634 351854 369718
rect 351234 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 351854 369634
rect 351234 355308 351854 369398
rect 354954 356614 355574 373000
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 355308 355574 356058
rect 338435 355060 338501 355061
rect 338435 354996 338436 355060
rect 338500 354996 338501 355060
rect 338435 354995 338501 354996
rect 350947 355060 351013 355061
rect 350947 354996 350948 355060
rect 351012 354996 351013 355060
rect 350947 354995 351013 354996
rect 338438 353970 338498 354995
rect 339723 354788 339789 354789
rect 339723 354724 339724 354788
rect 339788 354724 339789 354788
rect 339723 354723 339789 354724
rect 339726 353970 339786 354723
rect 350950 353970 351010 354995
rect 338438 353910 338524 353970
rect 338464 353260 338524 353910
rect 339688 353910 339786 353970
rect 350840 353910 351010 353970
rect 339688 353260 339748 353910
rect 350840 353260 350900 353910
rect 220272 345454 220620 345486
rect 220272 345218 220328 345454
rect 220564 345218 220620 345454
rect 220272 345134 220620 345218
rect 220272 344898 220328 345134
rect 220564 344898 220620 345134
rect 220272 344866 220620 344898
rect 356000 345454 356348 345486
rect 356000 345218 356056 345454
rect 356292 345218 356348 345454
rect 356000 345134 356348 345218
rect 356000 344898 356056 345134
rect 356292 344898 356348 345134
rect 356000 344866 356348 344898
rect 220952 327454 221300 327486
rect 220952 327218 221008 327454
rect 221244 327218 221300 327454
rect 220952 327134 221300 327218
rect 220952 326898 221008 327134
rect 221244 326898 221300 327134
rect 220952 326866 221300 326898
rect 355320 327454 355668 327486
rect 355320 327218 355376 327454
rect 355612 327218 355668 327454
rect 355320 327134 355668 327218
rect 355320 326898 355376 327134
rect 355612 326898 355668 327134
rect 355320 326866 355668 326898
rect 220272 309454 220620 309486
rect 220272 309218 220328 309454
rect 220564 309218 220620 309454
rect 220272 309134 220620 309218
rect 220272 308898 220328 309134
rect 220564 308898 220620 309134
rect 220272 308866 220620 308898
rect 356000 309454 356348 309486
rect 356000 309218 356056 309454
rect 356292 309218 356348 309454
rect 356000 309134 356348 309218
rect 356000 308898 356056 309134
rect 356292 308898 356348 309134
rect 356000 308866 356348 308898
rect 220952 291454 221300 291486
rect 220952 291218 221008 291454
rect 221244 291218 221300 291454
rect 220952 291134 221300 291218
rect 220952 290898 221008 291134
rect 221244 290898 221300 291134
rect 220952 290866 221300 290898
rect 355320 291454 355668 291486
rect 355320 291218 355376 291454
rect 355612 291218 355668 291454
rect 355320 291134 355668 291218
rect 355320 290898 355376 291134
rect 355612 290898 355668 291134
rect 355320 290866 355668 290898
rect 220272 273454 220620 273486
rect 220272 273218 220328 273454
rect 220564 273218 220620 273454
rect 220272 273134 220620 273218
rect 220272 272898 220328 273134
rect 220564 272898 220620 273134
rect 220272 272866 220620 272898
rect 356000 273454 356348 273486
rect 356000 273218 356056 273454
rect 356292 273218 356348 273454
rect 356000 273134 356348 273218
rect 356000 272898 356056 273134
rect 356292 272898 356348 273134
rect 356000 272866 356348 272898
rect 236056 269650 236116 270106
rect 237144 269650 237204 270106
rect 238232 269650 238292 270106
rect 239592 269650 239652 270106
rect 236056 269590 236562 269650
rect 221514 259174 222134 268000
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 250308 222134 258618
rect 225234 262894 225854 268000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 250308 225854 262338
rect 228954 266614 229574 268000
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 250308 229574 266058
rect 235794 256394 236414 268000
rect 236502 267069 236562 269590
rect 237054 269590 237204 269650
rect 238158 269590 238292 269650
rect 239262 269590 239652 269650
rect 240544 269650 240604 270106
rect 241768 269650 241828 270106
rect 243128 269650 243188 270106
rect 240544 269590 240610 269650
rect 236499 267068 236565 267069
rect 236499 267004 236500 267068
rect 236564 267004 236565 267068
rect 236499 267003 236565 267004
rect 237054 266933 237114 269590
rect 238158 267205 238218 269590
rect 238155 267204 238221 267205
rect 238155 267140 238156 267204
rect 238220 267140 238221 267204
rect 238155 267139 238221 267140
rect 237051 266932 237117 266933
rect 237051 266868 237052 266932
rect 237116 266868 237117 266932
rect 237051 266867 237117 266868
rect 239262 266253 239322 269590
rect 239259 266252 239325 266253
rect 239259 266188 239260 266252
rect 239324 266188 239325 266252
rect 239259 266187 239325 266188
rect 235794 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 236414 256394
rect 235794 256074 236414 256158
rect 235794 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 236414 256074
rect 235794 250308 236414 255838
rect 239514 260114 240134 268000
rect 240550 265709 240610 269590
rect 241654 269590 241828 269650
rect 243126 269590 243188 269650
rect 244216 269650 244276 270106
rect 245440 269650 245500 270106
rect 246528 269650 246588 270106
rect 244216 269590 244290 269650
rect 240547 265708 240613 265709
rect 240547 265644 240548 265708
rect 240612 265644 240613 265708
rect 240547 265643 240613 265644
rect 241654 265573 241714 269590
rect 243126 268837 243186 269590
rect 243123 268836 243189 268837
rect 243123 268772 243124 268836
rect 243188 268772 243189 268836
rect 243123 268771 243189 268772
rect 241651 265572 241717 265573
rect 241651 265508 241652 265572
rect 241716 265508 241717 265572
rect 241651 265507 241717 265508
rect 239514 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 240134 260114
rect 239514 259794 240134 259878
rect 239514 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 240134 259794
rect 239514 250308 240134 259558
rect 243234 261954 243854 268000
rect 244230 266525 244290 269590
rect 245334 269590 245500 269650
rect 246438 269590 246588 269650
rect 247616 269650 247676 270106
rect 248296 269650 248356 270106
rect 248704 269650 248764 270106
rect 247616 269590 247786 269650
rect 244227 266524 244293 266525
rect 244227 266460 244228 266524
rect 244292 266460 244293 266524
rect 244227 266459 244293 266460
rect 245334 266389 245394 269590
rect 246438 266389 246498 269590
rect 245331 266388 245397 266389
rect 245331 266324 245332 266388
rect 245396 266324 245397 266388
rect 245331 266323 245397 266324
rect 246435 266388 246501 266389
rect 246435 266324 246436 266388
rect 246500 266324 246501 266388
rect 246435 266323 246501 266324
rect 243234 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 243854 261954
rect 243234 261634 243854 261718
rect 243234 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 243854 261634
rect 243234 250308 243854 261398
rect 246954 265674 247574 268000
rect 247726 266389 247786 269590
rect 248278 269590 248356 269650
rect 248646 269590 248764 269650
rect 250064 269650 250124 270106
rect 250744 269925 250804 270106
rect 250741 269924 250807 269925
rect 250741 269860 250742 269924
rect 250806 269860 250807 269924
rect 250741 269859 250807 269860
rect 251288 269650 251348 270106
rect 252376 269650 252436 270106
rect 253464 269650 253524 270106
rect 250064 269590 250178 269650
rect 248278 266933 248338 269590
rect 248275 266932 248341 266933
rect 248275 266868 248276 266932
rect 248340 266868 248341 266932
rect 248275 266867 248341 266868
rect 248646 266389 248706 269590
rect 250118 266389 250178 269590
rect 251222 269590 251348 269650
rect 252326 269590 252436 269650
rect 253430 269590 253524 269650
rect 253600 269650 253660 270106
rect 254552 269650 254612 270106
rect 255912 269650 255972 270106
rect 253600 269590 253674 269650
rect 251222 266389 251282 269590
rect 252326 266525 252386 269590
rect 252323 266524 252389 266525
rect 252323 266460 252324 266524
rect 252388 266460 252389 266524
rect 252323 266459 252389 266460
rect 253430 266389 253490 269590
rect 253614 266933 253674 269590
rect 254534 269590 254612 269650
rect 255822 269590 255972 269650
rect 256048 269650 256108 270106
rect 257000 269650 257060 270106
rect 258088 269650 258148 270106
rect 258496 269650 258556 270106
rect 256048 269590 256250 269650
rect 253611 266932 253677 266933
rect 253611 266868 253612 266932
rect 253676 266868 253677 266932
rect 253611 266867 253677 266868
rect 247723 266388 247789 266389
rect 247723 266324 247724 266388
rect 247788 266324 247789 266388
rect 247723 266323 247789 266324
rect 248643 266388 248709 266389
rect 248643 266324 248644 266388
rect 248708 266324 248709 266388
rect 248643 266323 248709 266324
rect 250115 266388 250181 266389
rect 250115 266324 250116 266388
rect 250180 266324 250181 266388
rect 250115 266323 250181 266324
rect 251219 266388 251285 266389
rect 251219 266324 251220 266388
rect 251284 266324 251285 266388
rect 251219 266323 251285 266324
rect 253427 266388 253493 266389
rect 253427 266324 253428 266388
rect 253492 266324 253493 266388
rect 253427 266323 253493 266324
rect 246954 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 247574 265674
rect 246954 265354 247574 265438
rect 246954 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 247574 265354
rect 246954 250308 247574 265118
rect 253794 255454 254414 268000
rect 254534 266389 254594 269590
rect 255822 267749 255882 269590
rect 255819 267748 255885 267749
rect 255819 267684 255820 267748
rect 255884 267684 255885 267748
rect 255819 267683 255885 267684
rect 256190 267069 256250 269590
rect 256926 269590 257060 269650
rect 257846 269590 258148 269650
rect 258398 269590 258556 269650
rect 259448 269650 259508 270106
rect 260672 269650 260732 270106
rect 261080 269650 261140 270106
rect 261760 269650 261820 270106
rect 262848 269650 262908 270106
rect 259448 269590 259562 269650
rect 256187 267068 256253 267069
rect 256187 267004 256188 267068
rect 256252 267004 256253 267068
rect 256187 267003 256253 267004
rect 256926 266389 256986 269590
rect 257846 268837 257906 269590
rect 257843 268836 257909 268837
rect 257843 268772 257844 268836
rect 257908 268772 257909 268836
rect 257843 268771 257909 268772
rect 254531 266388 254597 266389
rect 254531 266324 254532 266388
rect 254596 266324 254597 266388
rect 254531 266323 254597 266324
rect 256923 266388 256989 266389
rect 256923 266324 256924 266388
rect 256988 266324 256989 266388
rect 256923 266323 256989 266324
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 250308 254414 254898
rect 257514 259174 258134 268000
rect 258398 267205 258458 269590
rect 258395 267204 258461 267205
rect 258395 267140 258396 267204
rect 258460 267140 258461 267204
rect 258395 267139 258461 267140
rect 259502 266389 259562 269590
rect 260606 269590 260732 269650
rect 260974 269590 261140 269650
rect 261710 269590 261820 269650
rect 262814 269590 262908 269650
rect 263528 269650 263588 270106
rect 263936 269650 263996 270106
rect 265296 269650 265356 270106
rect 265976 269650 266036 270106
rect 266384 269925 266444 270106
rect 266381 269924 266447 269925
rect 266381 269860 266382 269924
rect 266446 269860 266447 269924
rect 266381 269859 266447 269860
rect 267608 269650 267668 270106
rect 263528 269590 263794 269650
rect 260606 266525 260666 269590
rect 260974 267749 261034 269590
rect 261710 268837 261770 269590
rect 261707 268836 261773 268837
rect 261707 268772 261708 268836
rect 261772 268772 261773 268836
rect 261707 268771 261773 268772
rect 260971 267748 261037 267749
rect 260971 267684 260972 267748
rect 261036 267684 261037 267748
rect 260971 267683 261037 267684
rect 260603 266524 260669 266525
rect 260603 266460 260604 266524
rect 260668 266460 260669 266524
rect 260603 266459 260669 266460
rect 259499 266388 259565 266389
rect 259499 266324 259500 266388
rect 259564 266324 259565 266388
rect 259499 266323 259565 266324
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 250308 258134 258618
rect 261234 262894 261854 268000
rect 262814 266389 262874 269590
rect 263734 267749 263794 269590
rect 263918 269590 263996 269650
rect 265206 269590 265356 269650
rect 265942 269590 266036 269650
rect 267598 269590 267668 269650
rect 268288 269650 268348 270106
rect 268696 269650 268756 270106
rect 269784 269650 269844 270106
rect 271008 269650 271068 270106
rect 268288 269590 268394 269650
rect 268696 269590 268762 269650
rect 269784 269590 269866 269650
rect 263731 267748 263797 267749
rect 263731 267684 263732 267748
rect 263796 267684 263797 267748
rect 263731 267683 263797 267684
rect 263918 266933 263978 269590
rect 265206 268157 265266 269590
rect 265203 268156 265269 268157
rect 265203 268092 265204 268156
rect 265268 268092 265269 268156
rect 265203 268091 265269 268092
rect 263915 266932 263981 266933
rect 263915 266868 263916 266932
rect 263980 266868 263981 266932
rect 263915 266867 263981 266868
rect 264954 266614 265574 268000
rect 265942 267749 266002 269590
rect 267598 267749 267658 269590
rect 268334 267749 268394 269590
rect 265939 267748 266005 267749
rect 265939 267684 265940 267748
rect 266004 267684 266005 267748
rect 265939 267683 266005 267684
rect 267595 267748 267661 267749
rect 267595 267684 267596 267748
rect 267660 267684 267661 267748
rect 267595 267683 267661 267684
rect 268331 267748 268397 267749
rect 268331 267684 268332 267748
rect 268396 267684 268397 267748
rect 268331 267683 268397 267684
rect 268702 266933 268762 269590
rect 269806 267205 269866 269590
rect 270910 269590 271068 269650
rect 271144 269650 271204 270106
rect 272232 269650 272292 270106
rect 273320 269650 273380 270106
rect 273592 269650 273652 270106
rect 274408 269789 274468 270106
rect 275768 269789 275828 270106
rect 274405 269788 274471 269789
rect 274405 269724 274406 269788
rect 274470 269724 274471 269788
rect 274405 269723 274471 269724
rect 275765 269788 275831 269789
rect 275765 269724 275766 269788
rect 275830 269724 275831 269788
rect 275765 269723 275831 269724
rect 271144 269590 271338 269650
rect 270910 267749 270970 269590
rect 270907 267748 270973 267749
rect 270907 267684 270908 267748
rect 270972 267684 270973 267748
rect 270907 267683 270973 267684
rect 271278 267205 271338 269590
rect 272198 269590 272292 269650
rect 273302 269590 273380 269650
rect 273486 269590 273652 269650
rect 276040 269650 276100 270106
rect 276992 269650 277052 270106
rect 276040 269590 276306 269650
rect 272198 268157 272258 269590
rect 272195 268156 272261 268157
rect 272195 268092 272196 268156
rect 272260 268092 272261 268156
rect 272195 268091 272261 268092
rect 269803 267204 269869 267205
rect 269803 267140 269804 267204
rect 269868 267140 269869 267204
rect 269803 267139 269869 267140
rect 271275 267204 271341 267205
rect 271275 267140 271276 267204
rect 271340 267140 271341 267204
rect 271275 267139 271341 267140
rect 268699 266932 268765 266933
rect 268699 266868 268700 266932
rect 268764 266868 268765 266932
rect 268699 266867 268765 266868
rect 262811 266388 262877 266389
rect 262811 266324 262812 266388
rect 262876 266324 262877 266388
rect 262811 266323 262877 266324
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 250308 261854 262338
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 250308 265574 266058
rect 271794 256394 272414 268000
rect 273302 267069 273362 269590
rect 273486 267749 273546 269590
rect 273483 267748 273549 267749
rect 273483 267684 273484 267748
rect 273548 267684 273549 267748
rect 273483 267683 273549 267684
rect 273299 267068 273365 267069
rect 273299 267004 273300 267068
rect 273364 267004 273365 267068
rect 273299 267003 273365 267004
rect 271794 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 272414 256394
rect 271794 256074 272414 256158
rect 271794 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 272414 256074
rect 271794 250308 272414 255838
rect 275514 260114 276134 268000
rect 276246 267749 276306 269590
rect 276982 269590 277052 269650
rect 278080 269650 278140 270106
rect 278488 269650 278548 270106
rect 279168 269653 279228 270106
rect 280936 269789 280996 270106
rect 280933 269788 280999 269789
rect 280933 269724 280934 269788
rect 280998 269724 280999 269788
rect 280933 269723 280999 269724
rect 283520 269653 283580 270106
rect 285968 269653 286028 270106
rect 288280 269653 288340 270106
rect 279165 269652 279231 269653
rect 279165 269650 279166 269652
rect 278080 269590 278146 269650
rect 276243 267748 276309 267749
rect 276243 267684 276244 267748
rect 276308 267684 276309 267748
rect 276243 267683 276309 267684
rect 276982 267205 277042 269590
rect 278086 267205 278146 269590
rect 278454 269590 278548 269650
rect 279006 269590 279166 269650
rect 278454 268973 278514 269590
rect 278451 268972 278517 268973
rect 278451 268908 278452 268972
rect 278516 268908 278517 268972
rect 278451 268907 278517 268908
rect 276979 267204 277045 267205
rect 276979 267140 276980 267204
rect 277044 267140 277045 267204
rect 276979 267139 277045 267140
rect 278083 267204 278149 267205
rect 278083 267140 278084 267204
rect 278148 267140 278149 267204
rect 278083 267139 278149 267140
rect 279006 266389 279066 269590
rect 279165 269588 279166 269590
rect 279230 269588 279231 269652
rect 279165 269587 279231 269588
rect 283517 269652 283583 269653
rect 283517 269588 283518 269652
rect 283582 269588 283583 269652
rect 283517 269587 283583 269588
rect 285965 269652 286031 269653
rect 285965 269588 285966 269652
rect 286030 269588 286031 269652
rect 285965 269587 286031 269588
rect 288277 269652 288343 269653
rect 288277 269588 288278 269652
rect 288342 269588 288343 269652
rect 291000 269650 291060 270106
rect 293448 269653 293508 270106
rect 288277 269587 288343 269588
rect 290966 269590 291060 269650
rect 293445 269652 293511 269653
rect 290966 268973 291026 269590
rect 293445 269588 293446 269652
rect 293510 269588 293511 269652
rect 295896 269650 295956 270106
rect 298480 269650 298540 270106
rect 300928 269650 300988 270106
rect 303512 269650 303572 270106
rect 305960 269650 306020 270106
rect 308544 269653 308604 270106
rect 295896 269590 295994 269650
rect 298480 269590 298570 269650
rect 293445 269587 293511 269588
rect 295934 268973 295994 269590
rect 298510 269109 298570 269590
rect 300902 269590 300988 269650
rect 303478 269590 303572 269650
rect 305870 269590 306020 269650
rect 308541 269652 308607 269653
rect 300902 269109 300962 269590
rect 298507 269108 298573 269109
rect 298507 269044 298508 269108
rect 298572 269044 298573 269108
rect 298507 269043 298573 269044
rect 300899 269108 300965 269109
rect 300899 269044 300900 269108
rect 300964 269044 300965 269108
rect 300899 269043 300965 269044
rect 290963 268972 291029 268973
rect 290963 268908 290964 268972
rect 291028 268908 291029 268972
rect 290963 268907 291029 268908
rect 295931 268972 295997 268973
rect 295931 268908 295932 268972
rect 295996 268908 295997 268972
rect 295931 268907 295997 268908
rect 279003 266388 279069 266389
rect 279003 266324 279004 266388
rect 279068 266324 279069 266388
rect 279003 266323 279069 266324
rect 275514 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 276134 260114
rect 275514 259794 276134 259878
rect 275514 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 276134 259794
rect 275514 250308 276134 259558
rect 279234 261954 279854 268000
rect 279234 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 279854 261954
rect 279234 261634 279854 261718
rect 279234 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 279854 261634
rect 279234 250308 279854 261398
rect 282954 265674 283574 268000
rect 282954 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 283574 265674
rect 282954 265354 283574 265438
rect 282954 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 283574 265354
rect 282954 250308 283574 265118
rect 289794 255454 290414 268000
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 250308 290414 254898
rect 293514 259174 294134 268000
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 250308 294134 258618
rect 297234 262894 297854 268000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 250308 297854 262338
rect 300954 266614 301574 268000
rect 303478 267749 303538 269590
rect 305870 268973 305930 269590
rect 308541 269588 308542 269652
rect 308606 269588 308607 269652
rect 310992 269650 311052 270106
rect 313440 269650 313500 270106
rect 315888 269789 315948 270106
rect 315885 269788 315951 269789
rect 315885 269724 315886 269788
rect 315950 269724 315951 269788
rect 315885 269723 315951 269724
rect 318472 269653 318532 270106
rect 310992 269590 311082 269650
rect 308541 269587 308607 269588
rect 305867 268972 305933 268973
rect 305867 268908 305868 268972
rect 305932 268908 305933 268972
rect 305867 268907 305933 268908
rect 303475 267748 303541 267749
rect 303475 267684 303476 267748
rect 303540 267684 303541 267748
rect 303475 267683 303541 267684
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 250308 301574 266058
rect 307794 256394 308414 268000
rect 311022 266933 311082 269590
rect 313414 269590 313500 269650
rect 318469 269652 318535 269653
rect 311019 266932 311085 266933
rect 311019 266868 311020 266932
rect 311084 266868 311085 266932
rect 311019 266867 311085 266868
rect 307794 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 308414 256394
rect 307794 256074 308414 256158
rect 307794 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 308414 256074
rect 307794 250308 308414 255838
rect 311514 260114 312134 268000
rect 313414 267341 313474 269590
rect 318469 269588 318470 269652
rect 318534 269588 318535 269652
rect 320920 269650 320980 270106
rect 323368 269650 323428 270106
rect 320920 269590 321018 269650
rect 318469 269587 318535 269588
rect 313411 267340 313477 267341
rect 313411 267276 313412 267340
rect 313476 267276 313477 267340
rect 313411 267275 313477 267276
rect 311514 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 312134 260114
rect 311514 259794 312134 259878
rect 311514 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 312134 259794
rect 311514 250308 312134 259558
rect 315234 261954 315854 268000
rect 315234 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 315854 261954
rect 315234 261634 315854 261718
rect 315234 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 315854 261634
rect 315234 250308 315854 261398
rect 318954 265674 319574 268000
rect 320958 267477 321018 269590
rect 323350 269590 323428 269650
rect 325952 269650 326012 270106
rect 343224 269650 343284 270106
rect 325952 269590 326722 269650
rect 323350 267613 323410 269590
rect 323347 267612 323413 267613
rect 323347 267548 323348 267612
rect 323412 267548 323413 267612
rect 323347 267547 323413 267548
rect 320955 267476 321021 267477
rect 320955 267412 320956 267476
rect 321020 267412 321021 267476
rect 320955 267411 321021 267412
rect 318954 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 319574 265674
rect 318954 265354 319574 265438
rect 318954 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 319574 265354
rect 318954 250308 319574 265118
rect 325794 255454 326414 268000
rect 326662 266797 326722 269590
rect 343222 269590 343284 269650
rect 343360 269650 343420 270106
rect 343360 269590 343466 269650
rect 326659 266796 326725 266797
rect 326659 266732 326660 266796
rect 326724 266732 326725 266796
rect 326659 266731 326725 266732
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 250308 326414 254898
rect 329514 259174 330134 268000
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 250308 330134 258618
rect 333234 262894 333854 268000
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 250308 333854 262338
rect 336954 266614 337574 268000
rect 343222 267341 343282 269590
rect 343406 267477 343466 269590
rect 343403 267476 343469 267477
rect 343403 267412 343404 267476
rect 343468 267412 343469 267476
rect 343403 267411 343469 267412
rect 343219 267340 343285 267341
rect 343219 267276 343220 267340
rect 343284 267276 343285 267340
rect 343219 267275 343285 267276
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 250308 337574 266058
rect 343794 256394 344414 268000
rect 343794 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 344414 256394
rect 343794 256074 344414 256158
rect 343794 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 344414 256074
rect 343794 250308 344414 255838
rect 347514 260114 348134 268000
rect 347514 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 348134 260114
rect 347514 259794 348134 259878
rect 347514 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 348134 259794
rect 347514 250308 348134 259558
rect 351234 261954 351854 268000
rect 351234 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 351854 261954
rect 351234 261634 351854 261718
rect 351234 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 351854 261634
rect 351234 250308 351854 261398
rect 354954 265674 355574 268000
rect 354954 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 355574 265674
rect 354954 265354 355574 265438
rect 354954 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 355574 265354
rect 354954 250308 355574 265118
rect 338435 249932 338501 249933
rect 338435 249868 338436 249932
rect 338500 249868 338501 249932
rect 338435 249867 338501 249868
rect 339723 249932 339789 249933
rect 339723 249868 339724 249932
rect 339788 249868 339789 249932
rect 339723 249867 339789 249868
rect 350947 249932 351013 249933
rect 350947 249868 350948 249932
rect 351012 249868 351013 249932
rect 350947 249867 351013 249868
rect 338438 248430 338498 249867
rect 339726 248430 339786 249867
rect 350950 248430 351010 249867
rect 338438 248370 338524 248430
rect 338464 248202 338524 248370
rect 339688 248370 339786 248430
rect 350840 248370 351010 248430
rect 339688 248202 339748 248370
rect 350840 248202 350900 248370
rect 220272 237454 220620 237486
rect 220272 237218 220328 237454
rect 220564 237218 220620 237454
rect 220272 237134 220620 237218
rect 220272 236898 220328 237134
rect 220564 236898 220620 237134
rect 220272 236866 220620 236898
rect 356000 237454 356348 237486
rect 356000 237218 356056 237454
rect 356292 237218 356348 237454
rect 356000 237134 356348 237218
rect 356000 236898 356056 237134
rect 356292 236898 356348 237134
rect 356000 236866 356348 236898
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 201454 220620 201486
rect 220272 201218 220328 201454
rect 220564 201218 220620 201454
rect 220272 201134 220620 201218
rect 220272 200898 220328 201134
rect 220564 200898 220620 201134
rect 220272 200866 220620 200898
rect 356000 201454 356348 201486
rect 356000 201218 356056 201454
rect 356292 201218 356348 201454
rect 356000 201134 356348 201218
rect 356000 200898 356056 201134
rect 356292 200898 356348 201134
rect 356000 200866 356348 200898
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 164930 236116 165106
rect 237144 164930 237204 165106
rect 238232 164930 238292 165106
rect 235950 164870 236116 164930
rect 237054 164870 237204 164930
rect 238158 164870 238292 164930
rect 235950 163165 236010 164870
rect 235947 163164 236013 163165
rect 235947 163100 235948 163164
rect 236012 163100 236013 163164
rect 235947 163099 236013 163100
rect 221514 151174 222134 163000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 145308 222134 150618
rect 225234 154894 225854 163000
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 145308 225854 154338
rect 228954 158614 229574 163000
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 145308 229574 158058
rect 235794 148394 236414 163000
rect 237054 162757 237114 164870
rect 238158 162757 238218 164870
rect 239592 164658 239652 165106
rect 239446 164598 239652 164658
rect 240544 164658 240604 165106
rect 241768 164930 241828 165106
rect 241654 164870 241828 164930
rect 240544 164598 240610 164658
rect 239446 164250 239506 164598
rect 238526 164190 239506 164250
rect 237051 162756 237117 162757
rect 237051 162692 237052 162756
rect 237116 162692 237117 162756
rect 237051 162691 237117 162692
rect 238155 162756 238221 162757
rect 238155 162692 238156 162756
rect 238220 162692 238221 162756
rect 238155 162691 238221 162692
rect 238526 161530 238586 164190
rect 238707 161532 238773 161533
rect 238707 161530 238708 161532
rect 238526 161470 238708 161530
rect 238707 161468 238708 161470
rect 238772 161468 238773 161532
rect 238707 161467 238773 161468
rect 235794 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 236414 148394
rect 235794 148074 236414 148158
rect 235794 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 236414 148074
rect 235794 145308 236414 147838
rect 239514 152114 240134 163000
rect 240550 162757 240610 164598
rect 241654 162757 241714 164870
rect 243128 164658 243188 165106
rect 244216 164930 244276 165106
rect 245440 164930 245500 165106
rect 246528 164930 246588 165106
rect 244216 164870 244290 164930
rect 242942 164598 243188 164658
rect 242942 162757 243002 164598
rect 240547 162756 240613 162757
rect 240547 162692 240548 162756
rect 240612 162692 240613 162756
rect 240547 162691 240613 162692
rect 241651 162756 241717 162757
rect 241651 162692 241652 162756
rect 241716 162692 241717 162756
rect 241651 162691 241717 162692
rect 242939 162756 243005 162757
rect 242939 162692 242940 162756
rect 243004 162692 243005 162756
rect 242939 162691 243005 162692
rect 239514 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 240134 152114
rect 239514 151794 240134 151878
rect 239514 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 240134 151794
rect 239514 145308 240134 151558
rect 243234 153954 243854 163000
rect 244230 162757 244290 164870
rect 245334 164870 245500 164930
rect 246438 164870 246588 164930
rect 247616 164930 247676 165106
rect 247616 164870 247786 164930
rect 244227 162756 244293 162757
rect 244227 162692 244228 162756
rect 244292 162692 244293 162756
rect 244227 162691 244293 162692
rect 245334 162213 245394 164870
rect 246438 162757 246498 164870
rect 246435 162756 246501 162757
rect 246435 162692 246436 162756
rect 246500 162692 246501 162756
rect 246435 162691 246501 162692
rect 245331 162212 245397 162213
rect 245331 162148 245332 162212
rect 245396 162148 245397 162212
rect 245331 162147 245397 162148
rect 243234 153718 243266 153954
rect 243502 153718 243586 153954
rect 243822 153718 243854 153954
rect 243234 153634 243854 153718
rect 243234 153398 243266 153634
rect 243502 153398 243586 153634
rect 243822 153398 243854 153634
rect 243234 145308 243854 153398
rect 246954 157674 247574 163000
rect 247726 162757 247786 164870
rect 248296 164658 248356 165106
rect 248704 164658 248764 165106
rect 248278 164598 248356 164658
rect 248646 164598 248764 164658
rect 250064 164658 250124 165106
rect 250744 164930 250804 165106
rect 251288 164930 251348 165106
rect 250670 164870 250804 164930
rect 251222 164870 251348 164930
rect 250064 164598 250178 164658
rect 248278 162757 248338 164598
rect 248646 162757 248706 164598
rect 250118 162757 250178 164598
rect 247723 162756 247789 162757
rect 247723 162692 247724 162756
rect 247788 162692 247789 162756
rect 247723 162691 247789 162692
rect 248275 162756 248341 162757
rect 248275 162692 248276 162756
rect 248340 162692 248341 162756
rect 248275 162691 248341 162692
rect 248643 162756 248709 162757
rect 248643 162692 248644 162756
rect 248708 162692 248709 162756
rect 248643 162691 248709 162692
rect 250115 162756 250181 162757
rect 250115 162692 250116 162756
rect 250180 162692 250181 162756
rect 250115 162691 250181 162692
rect 250670 162349 250730 164870
rect 251222 162757 251282 164870
rect 252376 164658 252436 165106
rect 253464 164658 253524 165106
rect 252326 164598 252436 164658
rect 253430 164598 253524 164658
rect 253600 164658 253660 165106
rect 254552 164658 254612 165106
rect 255912 164930 255972 165106
rect 253600 164598 253674 164658
rect 251219 162756 251285 162757
rect 251219 162692 251220 162756
rect 251284 162692 251285 162756
rect 251219 162691 251285 162692
rect 252326 162485 252386 164598
rect 253430 162757 253490 164598
rect 253427 162756 253493 162757
rect 253427 162692 253428 162756
rect 253492 162692 253493 162756
rect 253427 162691 253493 162692
rect 252323 162484 252389 162485
rect 252323 162420 252324 162484
rect 252388 162420 252389 162484
rect 252323 162419 252389 162420
rect 253614 162349 253674 164598
rect 254534 164598 254612 164658
rect 255822 164870 255972 164930
rect 250667 162348 250733 162349
rect 250667 162284 250668 162348
rect 250732 162284 250733 162348
rect 250667 162283 250733 162284
rect 253611 162348 253677 162349
rect 253611 162284 253612 162348
rect 253676 162284 253677 162348
rect 253611 162283 253677 162284
rect 246954 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 247574 157674
rect 246954 157354 247574 157438
rect 246954 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 247574 157354
rect 246954 145308 247574 157118
rect 253794 147454 254414 163000
rect 254534 162757 254594 164598
rect 255822 162757 255882 164870
rect 256048 164658 256108 165106
rect 257000 164930 257060 165106
rect 256006 164598 256108 164658
rect 256926 164870 257060 164930
rect 258088 164930 258148 165106
rect 258088 164870 258274 164930
rect 256006 162757 256066 164598
rect 256926 162757 256986 164870
rect 254531 162756 254597 162757
rect 254531 162692 254532 162756
rect 254596 162692 254597 162756
rect 254531 162691 254597 162692
rect 255819 162756 255885 162757
rect 255819 162692 255820 162756
rect 255884 162692 255885 162756
rect 255819 162691 255885 162692
rect 256003 162756 256069 162757
rect 256003 162692 256004 162756
rect 256068 162692 256069 162756
rect 256003 162691 256069 162692
rect 256923 162756 256989 162757
rect 256923 162692 256924 162756
rect 256988 162692 256989 162756
rect 256923 162691 256989 162692
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 145308 254414 146898
rect 257514 151174 258134 163000
rect 258214 162210 258274 164870
rect 258496 164797 258556 165106
rect 259448 164930 259508 165106
rect 260672 164930 260732 165106
rect 259448 164870 259562 164930
rect 258493 164796 258559 164797
rect 258493 164732 258494 164796
rect 258558 164732 258559 164796
rect 258493 164731 258559 164732
rect 259502 162757 259562 164870
rect 260606 164870 260732 164930
rect 259499 162756 259565 162757
rect 259499 162692 259500 162756
rect 259564 162692 259565 162756
rect 259499 162691 259565 162692
rect 260606 162621 260666 164870
rect 261080 164661 261140 165106
rect 261760 164930 261820 165106
rect 262848 164930 262908 165106
rect 261710 164870 261820 164930
rect 262814 164870 262908 164930
rect 263528 164930 263588 165106
rect 263936 164930 263996 165106
rect 265296 164930 265356 165106
rect 265976 164930 266036 165106
rect 266384 164930 266444 165106
rect 267608 164930 267668 165106
rect 263528 164870 263610 164930
rect 261077 164660 261143 164661
rect 261077 164596 261078 164660
rect 261142 164596 261143 164660
rect 261077 164595 261143 164596
rect 261710 163165 261770 164870
rect 261707 163164 261773 163165
rect 261707 163100 261708 163164
rect 261772 163100 261773 163164
rect 261707 163099 261773 163100
rect 260603 162620 260669 162621
rect 260603 162556 260604 162620
rect 260668 162556 260669 162620
rect 260603 162555 260669 162556
rect 258395 162212 258461 162213
rect 258395 162210 258396 162212
rect 258214 162150 258396 162210
rect 258395 162148 258396 162150
rect 258460 162148 258461 162212
rect 258395 162147 258461 162148
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 145308 258134 150618
rect 261234 154894 261854 163000
rect 262814 162757 262874 164870
rect 262811 162756 262877 162757
rect 262811 162692 262812 162756
rect 262876 162692 262877 162756
rect 262811 162691 262877 162692
rect 263550 162621 263610 164870
rect 263918 164870 263996 164930
rect 265206 164870 265356 164930
rect 265942 164870 266036 164930
rect 266310 164870 266444 164930
rect 267598 164870 267668 164930
rect 263918 162757 263978 164870
rect 265206 163165 265266 164870
rect 265203 163164 265269 163165
rect 265203 163100 265204 163164
rect 265268 163100 265269 163164
rect 265203 163099 265269 163100
rect 263915 162756 263981 162757
rect 263915 162692 263916 162756
rect 263980 162692 263981 162756
rect 263915 162691 263981 162692
rect 263547 162620 263613 162621
rect 263547 162556 263548 162620
rect 263612 162556 263613 162620
rect 263547 162555 263613 162556
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 145308 261854 154338
rect 264954 158614 265574 163000
rect 265942 162757 266002 164870
rect 266310 162757 266370 164870
rect 267598 162757 267658 164870
rect 268288 164658 268348 165106
rect 268696 164658 268756 165106
rect 269784 164658 269844 165106
rect 271008 164930 271068 165106
rect 270910 164870 271068 164930
rect 268288 164598 268394 164658
rect 268696 164598 268762 164658
rect 269784 164598 269866 164658
rect 265939 162756 266005 162757
rect 265939 162692 265940 162756
rect 266004 162692 266005 162756
rect 265939 162691 266005 162692
rect 266307 162756 266373 162757
rect 266307 162692 266308 162756
rect 266372 162692 266373 162756
rect 266307 162691 266373 162692
rect 267595 162756 267661 162757
rect 267595 162692 267596 162756
rect 267660 162692 267661 162756
rect 267595 162691 267661 162692
rect 268334 162621 268394 164598
rect 268702 162757 268762 164598
rect 269806 162757 269866 164598
rect 270910 163437 270970 164870
rect 271144 164658 271204 165106
rect 272232 164658 272292 165106
rect 273320 164658 273380 165106
rect 273592 164930 273652 165106
rect 271094 164598 271204 164658
rect 272198 164598 272292 164658
rect 273302 164598 273380 164658
rect 273486 164870 273652 164930
rect 270907 163436 270973 163437
rect 270907 163372 270908 163436
rect 270972 163372 270973 163436
rect 270907 163371 270973 163372
rect 271094 162757 271154 164598
rect 272198 163165 272258 164598
rect 272195 163164 272261 163165
rect 272195 163100 272196 163164
rect 272260 163100 272261 163164
rect 272195 163099 272261 163100
rect 268699 162756 268765 162757
rect 268699 162692 268700 162756
rect 268764 162692 268765 162756
rect 268699 162691 268765 162692
rect 269803 162756 269869 162757
rect 269803 162692 269804 162756
rect 269868 162692 269869 162756
rect 269803 162691 269869 162692
rect 271091 162756 271157 162757
rect 271091 162692 271092 162756
rect 271156 162692 271157 162756
rect 271091 162691 271157 162692
rect 268331 162620 268397 162621
rect 268331 162556 268332 162620
rect 268396 162556 268397 162620
rect 268331 162555 268397 162556
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 145308 265574 158058
rect 271794 148394 272414 163000
rect 273302 162621 273362 164598
rect 273299 162620 273365 162621
rect 273299 162556 273300 162620
rect 273364 162556 273365 162620
rect 273299 162555 273365 162556
rect 273486 162349 273546 164870
rect 274408 164658 274468 165106
rect 275768 164661 275828 165106
rect 274406 164598 274468 164658
rect 275765 164660 275831 164661
rect 274406 162757 274466 164598
rect 275765 164596 275766 164660
rect 275830 164596 275831 164660
rect 276040 164658 276100 165106
rect 276992 164658 277052 165106
rect 278080 164930 278140 165106
rect 276040 164598 276306 164658
rect 275765 164595 275831 164596
rect 274403 162756 274469 162757
rect 274403 162692 274404 162756
rect 274468 162692 274469 162756
rect 274403 162691 274469 162692
rect 273483 162348 273549 162349
rect 273483 162284 273484 162348
rect 273548 162284 273549 162348
rect 273483 162283 273549 162284
rect 271794 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 272414 148394
rect 271794 148074 272414 148158
rect 271794 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 272414 148074
rect 271794 145308 272414 147838
rect 275514 152114 276134 163000
rect 276246 162485 276306 164598
rect 276982 164598 277052 164658
rect 277166 164870 278140 164930
rect 276982 162757 277042 164598
rect 276979 162756 277045 162757
rect 276979 162692 276980 162756
rect 277044 162692 277045 162756
rect 276979 162691 277045 162692
rect 276243 162484 276309 162485
rect 276243 162420 276244 162484
rect 276308 162420 276309 162484
rect 276243 162419 276309 162420
rect 277166 161530 277226 164870
rect 278488 164658 278548 165106
rect 279168 164658 279228 165106
rect 280936 164930 280996 165106
rect 278454 164598 278548 164658
rect 279006 164598 279228 164658
rect 280846 164870 280996 164930
rect 278454 162757 278514 164598
rect 279006 162757 279066 164598
rect 278451 162756 278517 162757
rect 278451 162692 278452 162756
rect 278516 162692 278517 162756
rect 278451 162691 278517 162692
rect 279003 162756 279069 162757
rect 279003 162692 279004 162756
rect 279068 162692 279069 162756
rect 279003 162691 279069 162692
rect 277347 161532 277413 161533
rect 277347 161530 277348 161532
rect 277166 161470 277348 161530
rect 277347 161468 277348 161470
rect 277412 161468 277413 161532
rect 277347 161467 277413 161468
rect 275514 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 276134 152114
rect 275514 151794 276134 151878
rect 275514 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 276134 151794
rect 275514 145308 276134 151558
rect 279234 153954 279854 163000
rect 280846 162757 280906 164870
rect 283520 164658 283580 165106
rect 285968 164658 286028 165106
rect 288280 164661 288340 165106
rect 291000 164930 291060 165106
rect 293448 164930 293508 165106
rect 290966 164870 291060 164930
rect 293358 164870 293508 164930
rect 288277 164660 288343 164661
rect 283520 164598 283850 164658
rect 285968 164598 286058 164658
rect 280843 162756 280909 162757
rect 280843 162692 280844 162756
rect 280908 162692 280909 162756
rect 280843 162691 280909 162692
rect 279234 153718 279266 153954
rect 279502 153718 279586 153954
rect 279822 153718 279854 153954
rect 279234 153634 279854 153718
rect 279234 153398 279266 153634
rect 279502 153398 279586 153634
rect 279822 153398 279854 153634
rect 279234 145308 279854 153398
rect 282954 157674 283574 163000
rect 283790 162757 283850 164598
rect 285998 162757 286058 164598
rect 288277 164596 288278 164660
rect 288342 164596 288343 164660
rect 288277 164595 288343 164596
rect 290966 163573 291026 164870
rect 290963 163572 291029 163573
rect 290963 163508 290964 163572
rect 291028 163508 291029 163572
rect 290963 163507 291029 163508
rect 283787 162756 283853 162757
rect 283787 162692 283788 162756
rect 283852 162692 283853 162756
rect 283787 162691 283853 162692
rect 285995 162756 286061 162757
rect 285995 162692 285996 162756
rect 286060 162692 286061 162756
rect 285995 162691 286061 162692
rect 282954 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 283574 157674
rect 282954 157354 283574 157438
rect 282954 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 283574 157354
rect 282954 145308 283574 157118
rect 289794 147454 290414 163000
rect 293358 162757 293418 164870
rect 295896 164797 295956 165106
rect 298480 164930 298540 165106
rect 300928 164930 300988 165106
rect 303512 164930 303572 165106
rect 298480 164870 298570 164930
rect 295893 164796 295959 164797
rect 295893 164732 295894 164796
rect 295958 164732 295959 164796
rect 295893 164731 295959 164732
rect 298510 164253 298570 164870
rect 300902 164870 300988 164930
rect 303478 164870 303572 164930
rect 300902 164253 300962 164870
rect 298507 164252 298573 164253
rect 298507 164188 298508 164252
rect 298572 164188 298573 164252
rect 298507 164187 298573 164188
rect 300899 164252 300965 164253
rect 300899 164188 300900 164252
rect 300964 164188 300965 164252
rect 300899 164187 300965 164188
rect 293355 162756 293421 162757
rect 293355 162692 293356 162756
rect 293420 162692 293421 162756
rect 293355 162691 293421 162692
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 145308 290414 146898
rect 293514 151174 294134 163000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 145308 294134 150618
rect 297234 154894 297854 163000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 145308 297854 154338
rect 300954 158614 301574 163000
rect 303478 162757 303538 164870
rect 305960 164661 306020 165106
rect 308544 164930 308604 165106
rect 310992 164930 311052 165106
rect 313440 164930 313500 165106
rect 315888 164930 315948 165106
rect 308544 164870 308690 164930
rect 310992 164870 311082 164930
rect 305957 164660 306023 164661
rect 305957 164596 305958 164660
rect 306022 164596 306023 164660
rect 305957 164595 306023 164596
rect 303475 162756 303541 162757
rect 303475 162692 303476 162756
rect 303540 162692 303541 162756
rect 303475 162691 303541 162692
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 145308 301574 158058
rect 307794 148394 308414 163000
rect 308630 162757 308690 164870
rect 311022 163981 311082 164870
rect 313414 164870 313500 164930
rect 315806 164870 315948 164930
rect 311019 163980 311085 163981
rect 311019 163916 311020 163980
rect 311084 163916 311085 163980
rect 311019 163915 311085 163916
rect 313414 163845 313474 164870
rect 313411 163844 313477 163845
rect 313411 163780 313412 163844
rect 313476 163780 313477 163844
rect 313411 163779 313477 163780
rect 315806 163709 315866 164870
rect 318472 164661 318532 165106
rect 320920 164930 320980 165106
rect 323368 164930 323428 165106
rect 325952 164930 326012 165106
rect 343224 164930 343284 165106
rect 320920 164870 321018 164930
rect 318469 164660 318535 164661
rect 318469 164596 318470 164660
rect 318534 164596 318535 164660
rect 318469 164595 318535 164596
rect 315803 163708 315869 163709
rect 315803 163644 315804 163708
rect 315868 163644 315869 163708
rect 315803 163643 315869 163644
rect 308627 162756 308693 162757
rect 308627 162692 308628 162756
rect 308692 162692 308693 162756
rect 308627 162691 308693 162692
rect 307794 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 308414 148394
rect 307794 148074 308414 148158
rect 307794 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 308414 148074
rect 307794 145308 308414 147838
rect 311514 152114 312134 163000
rect 311514 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 312134 152114
rect 311514 151794 312134 151878
rect 311514 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 312134 151794
rect 311514 145308 312134 151558
rect 315234 153954 315854 163000
rect 315234 153718 315266 153954
rect 315502 153718 315586 153954
rect 315822 153718 315854 153954
rect 315234 153634 315854 153718
rect 315234 153398 315266 153634
rect 315502 153398 315586 153634
rect 315822 153398 315854 153634
rect 315234 145308 315854 153398
rect 318954 157674 319574 163000
rect 320958 162621 321018 164870
rect 323350 164870 323428 164930
rect 325926 164870 326012 164930
rect 343222 164870 343284 164930
rect 343360 164930 343420 165106
rect 343360 164870 343466 164930
rect 323350 164117 323410 164870
rect 323347 164116 323413 164117
rect 323347 164052 323348 164116
rect 323412 164052 323413 164116
rect 323347 164051 323413 164052
rect 325926 163165 325986 164870
rect 325923 163164 325989 163165
rect 325923 163100 325924 163164
rect 325988 163100 325989 163164
rect 325923 163099 325989 163100
rect 320955 162620 321021 162621
rect 320955 162556 320956 162620
rect 321020 162556 321021 162620
rect 320955 162555 321021 162556
rect 318954 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 319574 157674
rect 318954 157354 319574 157438
rect 318954 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 319574 157354
rect 318954 145308 319574 157118
rect 325794 147454 326414 163000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 145308 326414 146898
rect 329514 151174 330134 163000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 145308 330134 150618
rect 333234 154894 333854 163000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 145308 333854 154338
rect 336954 158614 337574 163000
rect 343222 162621 343282 164870
rect 343406 162757 343466 164870
rect 343403 162756 343469 162757
rect 343403 162692 343404 162756
rect 343468 162692 343469 162756
rect 343403 162691 343469 162692
rect 343219 162620 343285 162621
rect 343219 162556 343220 162620
rect 343284 162556 343285 162620
rect 343219 162555 343285 162556
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 145308 337574 158058
rect 343794 148394 344414 163000
rect 343794 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 344414 148394
rect 343794 148074 344414 148158
rect 343794 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 344414 148074
rect 343794 145308 344414 147838
rect 347514 152114 348134 163000
rect 347514 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 348134 152114
rect 347514 151794 348134 151878
rect 347514 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 348134 151794
rect 347514 145308 348134 151558
rect 351234 153954 351854 163000
rect 351234 153718 351266 153954
rect 351502 153718 351586 153954
rect 351822 153718 351854 153954
rect 351234 153634 351854 153718
rect 351234 153398 351266 153634
rect 351502 153398 351586 153634
rect 351822 153398 351854 153634
rect 351234 145308 351854 153398
rect 354954 157674 355574 163000
rect 354954 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 355574 157674
rect 354954 157354 355574 157438
rect 354954 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 355574 157354
rect 354954 145308 355574 157118
rect 338435 144940 338501 144941
rect 338435 144876 338436 144940
rect 338500 144876 338501 144940
rect 338435 144875 338501 144876
rect 339723 144940 339789 144941
rect 339723 144876 339724 144940
rect 339788 144876 339789 144940
rect 339723 144875 339789 144876
rect 350947 144940 351013 144941
rect 350947 144876 350948 144940
rect 351012 144876 351013 144940
rect 350947 144875 351013 144876
rect 338438 143850 338498 144875
rect 339726 143850 339786 144875
rect 350950 143850 351010 144875
rect 338438 143790 338524 143850
rect 338464 143202 338524 143790
rect 339688 143790 339786 143850
rect 350840 143790 351010 143850
rect 339688 143202 339748 143790
rect 350840 143202 350900 143790
rect 220272 129454 220620 129486
rect 220272 129218 220328 129454
rect 220564 129218 220620 129454
rect 220272 129134 220620 129218
rect 220272 128898 220328 129134
rect 220564 128898 220620 129134
rect 220272 128866 220620 128898
rect 356000 129454 356348 129486
rect 356000 129218 356056 129454
rect 356292 129218 356348 129454
rect 356000 129134 356348 129218
rect 356000 128898 356056 129134
rect 356292 128898 356348 129134
rect 356000 128866 356348 128898
rect 220952 111454 221300 111486
rect 220952 111218 221008 111454
rect 221244 111218 221300 111454
rect 220952 111134 221300 111218
rect 220952 110898 221008 111134
rect 221244 110898 221300 111134
rect 220952 110866 221300 110898
rect 355320 111454 355668 111486
rect 355320 111218 355376 111454
rect 355612 111218 355668 111454
rect 355320 111134 355668 111218
rect 355320 110898 355376 111134
rect 355612 110898 355668 111134
rect 355320 110866 355668 110898
rect 220272 93454 220620 93486
rect 220272 93218 220328 93454
rect 220564 93218 220620 93454
rect 220272 93134 220620 93218
rect 220272 92898 220328 93134
rect 220564 92898 220620 93134
rect 220272 92866 220620 92898
rect 356000 93454 356348 93486
rect 356000 93218 356056 93454
rect 356292 93218 356348 93454
rect 356000 93134 356348 93218
rect 356000 92898 356056 93134
rect 356292 92898 356348 93134
rect 356000 92866 356348 92898
rect 220952 75454 221300 75486
rect 220952 75218 221008 75454
rect 221244 75218 221300 75454
rect 220952 75134 221300 75218
rect 220952 74898 221008 75134
rect 221244 74898 221300 75134
rect 220952 74866 221300 74898
rect 355320 75454 355668 75486
rect 355320 75218 355376 75454
rect 355612 75218 355668 75454
rect 355320 75134 355668 75218
rect 355320 74898 355376 75134
rect 355612 74898 355668 75134
rect 355320 74866 355668 74898
rect 236056 59530 236116 60106
rect 237144 59805 237204 60106
rect 237141 59804 237207 59805
rect 237141 59740 237142 59804
rect 237206 59740 237207 59804
rect 237141 59739 237207 59740
rect 238232 59530 238292 60106
rect 239592 59530 239652 60106
rect 235950 59470 236116 59530
rect 238158 59470 238292 59530
rect 239262 59470 239652 59530
rect 240544 59530 240604 60106
rect 241768 59530 241828 60106
rect 243128 59530 243188 60106
rect 240544 59470 240610 59530
rect 235950 58173 236010 59470
rect 235947 58172 236013 58173
rect 235947 58108 235948 58172
rect 236012 58108 236013 58172
rect 235947 58107 236013 58108
rect 219939 56540 220005 56541
rect 219939 56476 219940 56540
rect 220004 56476 220005 56540
rect 219939 56475 220005 56476
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 238158 57901 238218 59470
rect 239262 57901 239322 59470
rect 238155 57900 238221 57901
rect 238155 57836 238156 57900
rect 238220 57836 238221 57900
rect 238155 57835 238221 57836
rect 239259 57900 239325 57901
rect 239259 57836 239260 57900
rect 239324 57836 239325 57900
rect 239259 57835 239325 57836
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 240550 57493 240610 59470
rect 241654 59470 241828 59530
rect 242942 59470 243188 59530
rect 244216 59530 244276 60106
rect 245440 59530 245500 60106
rect 246528 59530 246588 60106
rect 244216 59470 244290 59530
rect 241654 57493 241714 59470
rect 242942 57901 243002 59470
rect 242939 57900 243005 57901
rect 242939 57836 242940 57900
rect 243004 57836 243005 57900
rect 242939 57835 243005 57836
rect 240547 57492 240613 57493
rect 240547 57428 240548 57492
rect 240612 57428 240613 57492
rect 240547 57427 240613 57428
rect 241651 57492 241717 57493
rect 241651 57428 241652 57492
rect 241716 57428 241717 57492
rect 241651 57427 241717 57428
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 244230 57493 244290 59470
rect 245334 59470 245500 59530
rect 246438 59470 246588 59530
rect 247616 59530 247676 60106
rect 248296 59530 248356 60106
rect 248704 59530 248764 60106
rect 247616 59470 247786 59530
rect 245334 57901 245394 59470
rect 246438 57901 246498 59470
rect 245331 57900 245397 57901
rect 245331 57836 245332 57900
rect 245396 57836 245397 57900
rect 245331 57835 245397 57836
rect 246435 57900 246501 57901
rect 246435 57836 246436 57900
rect 246500 57836 246501 57900
rect 246435 57835 246501 57836
rect 244227 57492 244293 57493
rect 244227 57428 244228 57492
rect 244292 57428 244293 57492
rect 244227 57427 244293 57428
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 247726 57493 247786 59470
rect 248278 59470 248356 59530
rect 248646 59470 248764 59530
rect 250064 59530 250124 60106
rect 250744 59530 250804 60106
rect 251288 59530 251348 60106
rect 252376 59530 252436 60106
rect 253464 59530 253524 60106
rect 250064 59470 250178 59530
rect 247723 57492 247789 57493
rect 247723 57428 247724 57492
rect 247788 57428 247789 57492
rect 247723 57427 247789 57428
rect 248278 56949 248338 59470
rect 248646 57901 248706 59470
rect 248643 57900 248709 57901
rect 248643 57836 248644 57900
rect 248708 57836 248709 57900
rect 248643 57835 248709 57836
rect 250118 57493 250178 59470
rect 250670 59470 250804 59530
rect 251222 59470 251348 59530
rect 252326 59470 252436 59530
rect 253430 59470 253524 59530
rect 253600 59530 253660 60106
rect 254552 59530 254612 60106
rect 255912 59805 255972 60106
rect 255909 59804 255975 59805
rect 255909 59740 255910 59804
rect 255974 59740 255975 59804
rect 255909 59739 255975 59740
rect 256048 59530 256108 60106
rect 257000 59669 257060 60106
rect 258088 59669 258148 60106
rect 256997 59668 257063 59669
rect 256997 59604 256998 59668
rect 257062 59604 257063 59668
rect 256997 59603 257063 59604
rect 258085 59668 258151 59669
rect 258085 59604 258086 59668
rect 258150 59604 258151 59668
rect 258085 59603 258151 59604
rect 258496 59530 258556 60106
rect 259448 59805 259508 60106
rect 260672 59805 260732 60106
rect 259445 59804 259511 59805
rect 259445 59740 259446 59804
rect 259510 59740 259511 59804
rect 259445 59739 259511 59740
rect 260669 59804 260735 59805
rect 260669 59740 260670 59804
rect 260734 59740 260735 59804
rect 260669 59739 260735 59740
rect 261080 59530 261140 60106
rect 261760 59805 261820 60106
rect 261757 59804 261823 59805
rect 261757 59740 261758 59804
rect 261822 59740 261823 59804
rect 261757 59739 261823 59740
rect 262848 59533 262908 60106
rect 253600 59470 253674 59530
rect 250115 57492 250181 57493
rect 250115 57428 250116 57492
rect 250180 57428 250181 57492
rect 250115 57427 250181 57428
rect 250670 57085 250730 59470
rect 251222 57901 251282 59470
rect 251219 57900 251285 57901
rect 251219 57836 251220 57900
rect 251284 57836 251285 57900
rect 251219 57835 251285 57836
rect 252326 57493 252386 59470
rect 253430 57901 253490 59470
rect 253427 57900 253493 57901
rect 253427 57836 253428 57900
rect 253492 57836 253493 57900
rect 253427 57835 253493 57836
rect 252323 57492 252389 57493
rect 252323 57428 252324 57492
rect 252388 57428 252389 57492
rect 252323 57427 252389 57428
rect 253614 57221 253674 59470
rect 254534 59470 254612 59530
rect 256006 59470 256108 59530
rect 258398 59470 258556 59530
rect 260974 59470 261140 59530
rect 262811 59532 262908 59533
rect 253611 57220 253677 57221
rect 253611 57156 253612 57220
rect 253676 57156 253677 57220
rect 253611 57155 253677 57156
rect 250667 57084 250733 57085
rect 250667 57020 250668 57084
rect 250732 57020 250733 57084
rect 250667 57019 250733 57020
rect 248275 56948 248341 56949
rect 248275 56884 248276 56948
rect 248340 56884 248341 56948
rect 248275 56883 248341 56884
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 254534 57493 254594 59470
rect 256006 58445 256066 59470
rect 256003 58444 256069 58445
rect 256003 58380 256004 58444
rect 256068 58380 256069 58444
rect 256003 58379 256069 58380
rect 254531 57492 254597 57493
rect 254531 57428 254532 57492
rect 254596 57428 254597 57492
rect 254531 57427 254597 57428
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 258398 57357 258458 59470
rect 260974 57629 261034 59470
rect 262811 59468 262812 59532
rect 262876 59470 262908 59532
rect 263528 59530 263588 60106
rect 263936 59805 263996 60106
rect 263933 59804 263999 59805
rect 263933 59740 263934 59804
rect 263998 59740 263999 59804
rect 263933 59739 263999 59740
rect 265296 59669 265356 60106
rect 265293 59668 265359 59669
rect 265293 59604 265294 59668
rect 265358 59604 265359 59668
rect 265293 59603 265359 59604
rect 265976 59530 266036 60106
rect 266384 59530 266444 60106
rect 267608 59530 267668 60106
rect 263528 59470 263610 59530
rect 262876 59468 262877 59470
rect 262811 59467 262877 59468
rect 263550 59397 263610 59470
rect 265942 59470 266036 59530
rect 266310 59470 266444 59530
rect 267598 59470 267668 59530
rect 268288 59530 268348 60106
rect 268696 59530 268756 60106
rect 269784 59530 269844 60106
rect 271008 59666 271068 60106
rect 270910 59606 271068 59666
rect 268288 59470 268394 59530
rect 268696 59470 268762 59530
rect 269784 59470 269866 59530
rect 263547 59396 263613 59397
rect 263547 59332 263548 59396
rect 263612 59332 263613 59396
rect 263547 59331 263613 59332
rect 260971 57628 261037 57629
rect 260971 57564 260972 57628
rect 261036 57564 261037 57628
rect 260971 57563 261037 57564
rect 258395 57356 258461 57357
rect 258395 57292 258396 57356
rect 258460 57292 258461 57356
rect 258395 57291 258461 57292
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 265942 57901 266002 59470
rect 266310 57901 266370 59470
rect 267598 57901 267658 59470
rect 268334 58581 268394 59470
rect 268331 58580 268397 58581
rect 268331 58516 268332 58580
rect 268396 58516 268397 58580
rect 268331 58515 268397 58516
rect 265939 57900 266005 57901
rect 265939 57836 265940 57900
rect 266004 57836 266005 57900
rect 265939 57835 266005 57836
rect 266307 57900 266373 57901
rect 266307 57836 266308 57900
rect 266372 57836 266373 57900
rect 266307 57835 266373 57836
rect 267595 57900 267661 57901
rect 267595 57836 267596 57900
rect 267660 57836 267661 57900
rect 267595 57835 267661 57836
rect 268702 57629 268762 59470
rect 269806 57901 269866 59470
rect 269803 57900 269869 57901
rect 269803 57836 269804 57900
rect 269868 57836 269869 57900
rect 269803 57835 269869 57836
rect 270910 57765 270970 59606
rect 271144 59530 271204 60106
rect 272232 59530 272292 60106
rect 273320 59530 273380 60106
rect 273592 59666 273652 60106
rect 271094 59470 271204 59530
rect 272198 59470 272292 59530
rect 273302 59470 273380 59530
rect 273486 59606 273652 59666
rect 270907 57764 270973 57765
rect 270907 57700 270908 57764
rect 270972 57700 270973 57764
rect 270907 57699 270973 57700
rect 271094 57629 271154 59470
rect 272198 58173 272258 59470
rect 272195 58172 272261 58173
rect 272195 58108 272196 58172
rect 272260 58108 272261 58172
rect 272195 58107 272261 58108
rect 268699 57628 268765 57629
rect 268699 57564 268700 57628
rect 268764 57564 268765 57628
rect 268699 57563 268765 57564
rect 271091 57628 271157 57629
rect 271091 57564 271092 57628
rect 271156 57564 271157 57628
rect 271091 57563 271157 57564
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 58000
rect 273302 57629 273362 59470
rect 273486 58853 273546 59606
rect 274408 59530 274468 60106
rect 275768 59666 275828 60106
rect 274406 59470 274468 59530
rect 275694 59606 275828 59666
rect 273483 58852 273549 58853
rect 273483 58788 273484 58852
rect 273548 58788 273549 58852
rect 273483 58787 273549 58788
rect 274406 57901 274466 59470
rect 275694 58173 275754 59606
rect 276040 59530 276100 60106
rect 276992 59530 277052 60106
rect 276040 59470 276122 59530
rect 276062 58717 276122 59470
rect 276982 59470 277052 59530
rect 278080 59530 278140 60106
rect 278488 59530 278548 60106
rect 279168 59530 279228 60106
rect 280936 59530 280996 60106
rect 278080 59470 278146 59530
rect 276059 58716 276125 58717
rect 276059 58652 276060 58716
rect 276124 58652 276125 58716
rect 276059 58651 276125 58652
rect 275691 58172 275757 58173
rect 275691 58108 275692 58172
rect 275756 58108 275757 58172
rect 275691 58107 275757 58108
rect 274403 57900 274469 57901
rect 274403 57836 274404 57900
rect 274468 57836 274469 57900
rect 274403 57835 274469 57836
rect 273299 57628 273365 57629
rect 273299 57564 273300 57628
rect 273364 57564 273365 57628
rect 273299 57563 273365 57564
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 276982 56405 277042 59470
rect 278086 57629 278146 59470
rect 278454 59470 278548 59530
rect 279006 59470 279228 59530
rect 280846 59470 280996 59530
rect 283520 59530 283580 60106
rect 285968 59530 286028 60106
rect 288280 59530 288340 60106
rect 291000 59530 291060 60106
rect 293448 59530 293508 60106
rect 283520 59470 283850 59530
rect 285968 59470 286058 59530
rect 278083 57628 278149 57629
rect 278083 57564 278084 57628
rect 278148 57564 278149 57628
rect 278083 57563 278149 57564
rect 278454 56813 278514 59470
rect 279006 57901 279066 59470
rect 280846 59125 280906 59470
rect 280843 59124 280909 59125
rect 280843 59060 280844 59124
rect 280908 59060 280909 59124
rect 280843 59059 280909 59060
rect 279003 57900 279069 57901
rect 279003 57836 279004 57900
rect 279068 57836 279069 57900
rect 279003 57835 279069 57836
rect 278451 56812 278517 56813
rect 278451 56748 278452 56812
rect 278516 56748 278517 56812
rect 278451 56747 278517 56748
rect 276979 56404 277045 56405
rect 276979 56340 276980 56404
rect 277044 56340 277045 56404
rect 276979 56339 277045 56340
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 283790 57901 283850 59470
rect 285998 59261 286058 59470
rect 288206 59470 288340 59530
rect 290966 59470 291060 59530
rect 293358 59470 293508 59530
rect 295896 59530 295956 60106
rect 298480 59530 298540 60106
rect 300928 59530 300988 60106
rect 303512 59530 303572 60106
rect 305960 59530 306020 60106
rect 295896 59470 295994 59530
rect 298480 59470 298570 59530
rect 285995 59260 286061 59261
rect 285995 59196 285996 59260
rect 286060 59196 286061 59260
rect 285995 59195 286061 59196
rect 288206 57901 288266 59470
rect 290966 58989 291026 59470
rect 290963 58988 291029 58989
rect 290963 58924 290964 58988
rect 291028 58924 291029 58988
rect 290963 58923 291029 58924
rect 283787 57900 283853 57901
rect 283787 57836 283788 57900
rect 283852 57836 283853 57900
rect 283787 57835 283853 57836
rect 288203 57900 288269 57901
rect 288203 57836 288204 57900
rect 288268 57836 288269 57900
rect 288203 57835 288269 57836
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 293358 57901 293418 59470
rect 295934 59261 295994 59470
rect 298510 59261 298570 59470
rect 300902 59470 300988 59530
rect 303478 59470 303572 59530
rect 305870 59470 306020 59530
rect 308544 59530 308604 60106
rect 310992 59530 311052 60106
rect 313440 59530 313500 60106
rect 315888 59669 315948 60106
rect 315885 59668 315951 59669
rect 315885 59604 315886 59668
rect 315950 59604 315951 59668
rect 318472 59666 318532 60106
rect 315885 59603 315951 59604
rect 318382 59606 318532 59666
rect 308544 59470 308690 59530
rect 310992 59470 311082 59530
rect 295931 59260 295997 59261
rect 295931 59196 295932 59260
rect 295996 59196 295997 59260
rect 295931 59195 295997 59196
rect 298507 59260 298573 59261
rect 298507 59196 298508 59260
rect 298572 59196 298573 59260
rect 298507 59195 298573 59196
rect 300902 58173 300962 59470
rect 303478 59261 303538 59470
rect 303475 59260 303541 59261
rect 303475 59196 303476 59260
rect 303540 59196 303541 59260
rect 303475 59195 303541 59196
rect 300899 58172 300965 58173
rect 300899 58108 300900 58172
rect 300964 58108 300965 58172
rect 300899 58107 300965 58108
rect 293355 57900 293421 57901
rect 293355 57836 293356 57900
rect 293420 57836 293421 57900
rect 293355 57835 293421 57836
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 305870 57901 305930 59470
rect 305867 57900 305933 57901
rect 305867 57836 305868 57900
rect 305932 57836 305933 57900
rect 305867 57835 305933 57836
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 308630 57629 308690 59470
rect 311022 57901 311082 59470
rect 313414 59470 313500 59530
rect 311019 57900 311085 57901
rect 311019 57836 311020 57900
rect 311084 57836 311085 57900
rect 311019 57835 311085 57836
rect 308627 57628 308693 57629
rect 308627 57564 308628 57628
rect 308692 57564 308693 57628
rect 308627 57563 308693 57564
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 313414 57901 313474 59470
rect 313411 57900 313477 57901
rect 313411 57836 313412 57900
rect 313476 57836 313477 57900
rect 313411 57835 313477 57836
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 318382 57901 318442 59606
rect 320920 59530 320980 60106
rect 323368 59530 323428 60106
rect 325952 59530 326012 60106
rect 343224 59530 343284 60106
rect 320920 59470 321018 59530
rect 318379 57900 318445 57901
rect 318379 57836 318380 57900
rect 318444 57836 318445 57900
rect 318379 57835 318445 57836
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 320958 57901 321018 59470
rect 323350 59470 323428 59530
rect 325926 59470 326012 59530
rect 343222 59470 343284 59530
rect 343360 59530 343420 60106
rect 343360 59470 343466 59530
rect 323350 59261 323410 59470
rect 323347 59260 323413 59261
rect 323347 59196 323348 59260
rect 323412 59196 323413 59260
rect 323347 59195 323413 59196
rect 325926 58173 325986 59470
rect 325923 58172 325989 58173
rect 325923 58108 325924 58172
rect 325988 58108 325989 58172
rect 325923 58107 325989 58108
rect 320955 57900 321021 57901
rect 320955 57836 320956 57900
rect 321020 57836 321021 57900
rect 320955 57835 321021 57836
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 343222 57901 343282 59470
rect 343406 57901 343466 59470
rect 357942 59261 358002 478755
rect 360147 478684 360213 478685
rect 360147 478620 360148 478684
rect 360212 478620 360213 478684
rect 360147 478619 360213 478620
rect 358123 472836 358189 472837
rect 358123 472772 358124 472836
rect 358188 472772 358189 472836
rect 358123 472771 358189 472772
rect 357939 59260 358005 59261
rect 357939 59196 357940 59260
rect 358004 59196 358005 59260
rect 357939 59195 358005 59196
rect 343219 57900 343285 57901
rect 343219 57836 343220 57900
rect 343284 57836 343285 57900
rect 343219 57835 343285 57836
rect 343403 57900 343469 57901
rect 343403 57836 343404 57900
rect 343468 57836 343469 57900
rect 343403 57835 343469 57836
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 358126 57765 358186 472771
rect 359595 471340 359661 471341
rect 359595 471276 359596 471340
rect 359660 471276 359661 471340
rect 359595 471275 359661 471276
rect 359411 468756 359477 468757
rect 359411 468692 359412 468756
rect 359476 468692 359477 468756
rect 359411 468691 359477 468692
rect 359414 269245 359474 468691
rect 359598 373693 359658 471275
rect 359963 465900 360029 465901
rect 359963 465836 359964 465900
rect 360028 465836 360029 465900
rect 359963 465835 360029 465836
rect 359779 463044 359845 463045
rect 359779 462980 359780 463044
rect 359844 462980 359845 463044
rect 359779 462979 359845 462980
rect 359595 373692 359661 373693
rect 359595 373628 359596 373692
rect 359660 373628 359661 373692
rect 359595 373627 359661 373628
rect 359782 371245 359842 462979
rect 359966 373285 360026 465835
rect 360150 408645 360210 478619
rect 360147 408644 360213 408645
rect 360147 408580 360148 408644
rect 360212 408580 360213 408644
rect 360147 408579 360213 408580
rect 359963 373284 360029 373285
rect 359963 373220 359964 373284
rect 360028 373220 360029 373284
rect 359963 373219 360029 373220
rect 359779 371244 359845 371245
rect 359779 371180 359780 371244
rect 359844 371180 359845 371244
rect 359779 371179 359845 371180
rect 359411 269244 359477 269245
rect 359411 269180 359412 269244
rect 359476 269180 359477 269244
rect 359411 269179 359477 269180
rect 360702 149157 360762 485011
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 365514 511174 366134 518000
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 369234 514894 369854 518000
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 367691 478548 367757 478549
rect 367691 478484 367692 478548
rect 367756 478484 367757 478548
rect 367691 478483 367757 478484
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 362907 468484 362973 468485
rect 362907 468420 362908 468484
rect 362972 468420 362973 468484
rect 362907 468419 362973 468420
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 362910 372741 362970 468419
rect 364931 465764 364997 465765
rect 364931 465700 364932 465764
rect 364996 465700 364997 465764
rect 364931 465699 364997 465700
rect 362907 372740 362973 372741
rect 362907 372676 362908 372740
rect 362972 372676 362973 372740
rect 362907 372675 362973 372676
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 360699 149156 360765 149157
rect 360699 149092 360700 149156
rect 360764 149092 360765 149156
rect 360699 149091 360765 149092
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 358123 57764 358189 57765
rect 358123 57700 358124 57764
rect 358188 57700 358189 57764
rect 358123 57699 358189 57700
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 74898
rect 364934 57493 364994 465699
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 364931 57492 364997 57493
rect 364931 57428 364932 57492
rect 364996 57428 364997 57492
rect 364931 57427 364997 57428
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 78618
rect 367694 59125 367754 478483
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 372954 482614 373574 518000
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 371739 478412 371805 478413
rect 371739 478348 371740 478412
rect 371804 478348 371805 478412
rect 371739 478347 371805 478348
rect 369234 442894 369854 478338
rect 370451 472700 370517 472701
rect 370451 472636 370452 472700
rect 370516 472636 370517 472700
rect 370451 472635 370517 472636
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 367691 59124 367757 59125
rect 367691 59060 367692 59124
rect 367756 59060 367757 59124
rect 367691 59059 367757 59060
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 82338
rect 370454 56677 370514 472635
rect 371742 58717 371802 478347
rect 372954 446614 373574 482058
rect 379794 489454 380414 518000
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 374499 478276 374565 478277
rect 374499 478212 374500 478276
rect 374564 478212 374565 478276
rect 374499 478211 374565 478212
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 357554 373574 374058
rect 372954 357318 372986 357554
rect 373222 357318 373306 357554
rect 373542 357318 373574 357554
rect 372954 357234 373574 357318
rect 372954 356998 372986 357234
rect 373222 356998 373306 357234
rect 373542 356998 373574 357234
rect 372954 338614 373574 356998
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 371739 58716 371805 58717
rect 371739 58652 371740 58716
rect 371804 58652 371805 58716
rect 371739 58651 371805 58652
rect 370451 56676 370517 56677
rect 370451 56612 370452 56676
rect 370516 56612 370517 56676
rect 370451 56611 370517 56612
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 86058
rect 374502 58989 374562 478211
rect 375971 478140 376037 478141
rect 375971 478076 375972 478140
rect 376036 478076 376037 478140
rect 375971 478075 376037 478076
rect 374499 58988 374565 58989
rect 374499 58924 374500 58988
rect 374564 58924 374565 58988
rect 374499 58923 374565 58924
rect 375974 58853 376034 478075
rect 377259 476780 377325 476781
rect 377259 476716 377260 476780
rect 377324 476716 377325 476780
rect 377259 476715 377325 476716
rect 376155 472564 376221 472565
rect 376155 472500 376156 472564
rect 376220 472500 376221 472564
rect 376155 472499 376221 472500
rect 375971 58852 376037 58853
rect 375971 58788 375972 58852
rect 376036 58788 376037 58852
rect 375971 58787 376037 58788
rect 376158 57629 376218 472499
rect 376891 464404 376957 464405
rect 376891 464340 376892 464404
rect 376956 464340 376957 464404
rect 376891 464339 376957 464340
rect 376894 372741 376954 464339
rect 376891 372740 376957 372741
rect 376891 372676 376892 372740
rect 376956 372676 376957 372740
rect 376891 372675 376957 372676
rect 376894 372469 376954 372675
rect 376891 372468 376957 372469
rect 376891 372404 376892 372468
rect 376956 372404 376957 372468
rect 376891 372403 376957 372404
rect 376891 368524 376957 368525
rect 376891 368460 376892 368524
rect 376956 368460 376957 368524
rect 376891 368459 376957 368460
rect 376894 269381 376954 368459
rect 376891 269380 376957 269381
rect 376891 269316 376892 269380
rect 376956 269316 376957 269380
rect 376891 269315 376957 269316
rect 377262 268973 377322 476715
rect 378731 475420 378797 475421
rect 378731 475356 378732 475420
rect 378796 475356 378797 475420
rect 378731 475355 378797 475356
rect 378179 474060 378245 474061
rect 378179 473996 378180 474060
rect 378244 473996 378245 474060
rect 378179 473995 378245 473996
rect 377443 469980 377509 469981
rect 377443 469916 377444 469980
rect 377508 469916 377509 469980
rect 377443 469915 377509 469916
rect 377446 373965 377506 469915
rect 377627 462908 377693 462909
rect 377627 462844 377628 462908
rect 377692 462844 377693 462908
rect 377627 462843 377693 462844
rect 377443 373964 377509 373965
rect 377443 373900 377444 373964
rect 377508 373900 377509 373964
rect 377443 373899 377509 373900
rect 377630 373829 377690 462843
rect 377627 373828 377693 373829
rect 377627 373764 377628 373828
rect 377692 373764 377693 373828
rect 377627 373763 377693 373764
rect 377811 371924 377877 371925
rect 377811 371860 377812 371924
rect 377876 371860 377877 371924
rect 377811 371859 377877 371860
rect 377627 269380 377693 269381
rect 377627 269316 377628 269380
rect 377692 269316 377693 269380
rect 377627 269315 377693 269316
rect 377259 268972 377325 268973
rect 377259 268908 377260 268972
rect 377324 268908 377325 268972
rect 377259 268907 377325 268908
rect 377630 268837 377690 269315
rect 377627 268836 377693 268837
rect 377627 268772 377628 268836
rect 377692 268772 377693 268836
rect 377627 268771 377693 268772
rect 377814 263533 377874 371859
rect 378182 270469 378242 473995
rect 378179 270468 378245 270469
rect 378179 270404 378180 270468
rect 378244 270404 378245 270468
rect 378179 270403 378245 270404
rect 377995 270332 378061 270333
rect 377995 270268 377996 270332
rect 378060 270268 378061 270332
rect 377995 270267 378061 270268
rect 377811 263532 377877 263533
rect 377811 263468 377812 263532
rect 377876 263468 377877 263532
rect 377811 263467 377877 263468
rect 377814 164253 377874 263467
rect 377811 164252 377877 164253
rect 377811 164188 377812 164252
rect 377876 164188 377877 164252
rect 377811 164187 377877 164188
rect 377259 158812 377325 158813
rect 377259 158748 377260 158812
rect 377324 158748 377325 158812
rect 377259 158747 377325 158748
rect 377262 58445 377322 158747
rect 377998 146301 378058 270267
rect 377995 146300 378061 146301
rect 377995 146236 377996 146300
rect 378060 146236 378061 146300
rect 377995 146235 378061 146236
rect 377443 143716 377509 143717
rect 377443 143652 377444 143716
rect 377508 143652 377509 143716
rect 377443 143651 377509 143652
rect 377259 58444 377325 58445
rect 377259 58380 377260 58444
rect 377324 58380 377325 58444
rect 377259 58379 377325 58380
rect 376155 57628 376221 57629
rect 376155 57564 376156 57628
rect 376220 57564 376221 57628
rect 376155 57563 376221 57564
rect 377446 55181 377506 143651
rect 377998 58581 378058 146235
rect 377995 58580 378061 58581
rect 377995 58516 377996 58580
rect 378060 58516 378061 58580
rect 377995 58515 378061 58516
rect 378734 57085 378794 475355
rect 378915 471204 378981 471205
rect 378915 471140 378916 471204
rect 378980 471140 378981 471204
rect 378915 471139 378981 471140
rect 378918 57357 378978 471139
rect 379099 469844 379165 469845
rect 379099 469780 379100 469844
rect 379164 469780 379165 469844
rect 379099 469779 379165 469780
rect 378915 57356 378981 57357
rect 378915 57292 378916 57356
rect 378980 57292 378981 57356
rect 378915 57291 378981 57292
rect 379102 57221 379162 469779
rect 379467 468620 379533 468621
rect 379467 468556 379468 468620
rect 379532 468556 379533 468620
rect 379467 468555 379533 468556
rect 379470 460950 379530 468555
rect 379470 460890 379714 460950
rect 379654 267750 379714 460890
rect 379794 460308 380414 488898
rect 383514 493174 384134 518000
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 460308 384134 492618
rect 387234 496894 387854 518000
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460308 387854 496338
rect 390954 500614 391574 518000
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 460308 391574 464058
rect 397794 507454 398414 518000
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 460308 398414 470898
rect 401514 511174 402134 518000
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 460308 402134 474618
rect 405234 514894 405854 518000
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 460308 405854 478338
rect 408954 482614 409574 518000
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 460308 409574 482058
rect 415794 489454 416414 518000
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 460308 416414 488898
rect 419514 493174 420134 518000
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 460308 420134 492618
rect 423234 496894 423854 518000
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460308 423854 496338
rect 426954 500614 427574 518000
rect 430806 517309 430866 592179
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 430803 517308 430869 517309
rect 430803 517244 430804 517308
rect 430868 517244 430869 517308
rect 430803 517243 430869 517244
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 460308 427574 464058
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 460308 434414 470898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 460308 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 460308 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 460308 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 460308 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 622000 459854 640338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 622000 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 622000 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 622000 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 622000 477854 622338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 622000 481574 626058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 622000 488414 632898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 622000 492134 636618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 622000 495854 640338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 622000 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 622000 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 622000 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 479568 597454 479888 597486
rect 479568 597218 479610 597454
rect 479846 597218 479888 597454
rect 479568 597134 479888 597218
rect 479568 596898 479610 597134
rect 479846 596898 479888 597134
rect 479568 596866 479888 596898
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 464208 579454 464528 579486
rect 464208 579218 464250 579454
rect 464486 579218 464528 579454
rect 464208 579134 464528 579218
rect 464208 578898 464250 579134
rect 464486 578898 464528 579134
rect 464208 578866 464528 578898
rect 494928 579454 495248 579486
rect 494928 579218 494970 579454
rect 495206 579218 495248 579454
rect 494928 579134 495248 579218
rect 494928 578898 494970 579134
rect 495206 578898 495248 579134
rect 494928 578866 495248 578898
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 460308 456134 492618
rect 459234 532894 459854 568000
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460308 459854 496338
rect 462954 536614 463574 568000
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 460308 463574 464058
rect 469794 543454 470414 568000
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 460308 470414 470898
rect 473514 547174 474134 568000
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 460308 474134 474618
rect 477234 550894 477854 568000
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 460308 477854 478338
rect 480954 554614 481574 568000
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 460308 481574 482058
rect 487794 561454 488414 568000
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 460308 488414 488898
rect 491514 565174 492134 568000
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 460308 492134 492618
rect 495234 532894 495854 568000
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460308 495854 496338
rect 498954 536614 499574 568000
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498515 461004 498581 461005
rect 498515 460940 498516 461004
rect 498580 460940 498581 461004
rect 498515 460939 498581 460940
rect 498518 458690 498578 460939
rect 498954 460308 499574 464058
rect 505794 543454 506414 568000
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 499803 461004 499869 461005
rect 499803 460940 499804 461004
rect 499868 460940 499869 461004
rect 499803 460939 499869 460940
rect 499806 458690 499866 460939
rect 505794 460308 506414 470898
rect 509514 547174 510134 568000
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 460308 510134 474618
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 510843 462228 510909 462229
rect 510843 462164 510844 462228
rect 510908 462164 510909 462228
rect 510843 462163 510909 462164
rect 510846 458690 510906 462163
rect 513234 460308 513854 478338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 460308 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 498464 458630 498578 458690
rect 499688 458630 499866 458690
rect 510840 458630 510906 458690
rect 498464 458202 498524 458630
rect 499688 458202 499748 458630
rect 510840 458202 510900 458630
rect 380272 453454 380620 453486
rect 380272 453218 380328 453454
rect 380564 453218 380620 453454
rect 380272 453134 380620 453218
rect 380272 452898 380328 453134
rect 380564 452898 380620 453134
rect 380272 452866 380620 452898
rect 516000 453454 516348 453486
rect 516000 453218 516056 453454
rect 516292 453218 516348 453454
rect 516000 453134 516348 453218
rect 516000 452898 516056 453134
rect 516292 452898 516348 453134
rect 516000 452866 516348 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 380952 435454 381300 435486
rect 380952 435218 381008 435454
rect 381244 435218 381300 435454
rect 380952 435134 381300 435218
rect 380952 434898 381008 435134
rect 381244 434898 381300 435134
rect 380952 434866 381300 434898
rect 515320 435454 515668 435486
rect 515320 435218 515376 435454
rect 515612 435218 515668 435454
rect 515320 435134 515668 435218
rect 515320 434898 515376 435134
rect 515612 434898 515668 435134
rect 515320 434866 515668 434898
rect 380272 417454 380620 417486
rect 380272 417218 380328 417454
rect 380564 417218 380620 417454
rect 380272 417134 380620 417218
rect 380272 416898 380328 417134
rect 380564 416898 380620 417134
rect 380272 416866 380620 416898
rect 516000 417454 516348 417486
rect 516000 417218 516056 417454
rect 516292 417218 516348 417454
rect 516000 417134 516348 417218
rect 516000 416898 516056 417134
rect 516292 416898 516348 417134
rect 516000 416866 516348 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 380952 399454 381300 399486
rect 380952 399218 381008 399454
rect 381244 399218 381300 399454
rect 380952 399134 381300 399218
rect 380952 398898 381008 399134
rect 381244 398898 381300 399134
rect 380952 398866 381300 398898
rect 515320 399454 515668 399486
rect 515320 399218 515376 399454
rect 515612 399218 515668 399454
rect 515320 399134 515668 399218
rect 515320 398898 515376 399134
rect 515612 398898 515668 399134
rect 515320 398866 515668 398898
rect 380272 381454 380620 381486
rect 380272 381218 380328 381454
rect 380564 381218 380620 381454
rect 380272 381134 380620 381218
rect 380272 380898 380328 381134
rect 380564 380898 380620 381134
rect 380272 380866 380620 380898
rect 516000 381454 516348 381486
rect 516000 381218 516056 381454
rect 516292 381218 516348 381454
rect 516000 381134 516348 381218
rect 516000 380898 516056 381134
rect 516292 380898 516348 381134
rect 516000 380866 516348 380898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 405963 375052 406029 375053
rect 396086 374990 396274 375050
rect 379794 364394 380414 373000
rect 379794 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 380414 364394
rect 379794 364074 380414 364158
rect 379794 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 380414 364074
rect 379794 355308 380414 363838
rect 383514 366234 384134 373000
rect 383514 365998 383546 366234
rect 383782 365998 383866 366234
rect 384102 365998 384134 366234
rect 383514 365914 384134 365998
rect 383514 365678 383546 365914
rect 383782 365678 383866 365914
rect 384102 365678 384134 365914
rect 383514 355308 384134 365678
rect 387234 369954 387854 373000
rect 387234 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 387854 369954
rect 387234 369634 387854 369718
rect 387234 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 387854 369634
rect 387234 355308 387854 369398
rect 390954 356614 391574 373000
rect 396214 372197 396274 374990
rect 396582 374990 397174 375050
rect 397502 374990 398262 375050
rect 398974 374990 399622 375050
rect 400262 374990 400574 375050
rect 401798 374990 402346 375050
rect 396211 372196 396277 372197
rect 396211 372132 396212 372196
rect 396276 372132 396277 372196
rect 396211 372131 396277 372132
rect 396582 371381 396642 374990
rect 397502 372061 397562 374990
rect 397499 372060 397565 372061
rect 397499 371996 397500 372060
rect 397564 371996 397565 372060
rect 397499 371995 397565 371996
rect 396579 371380 396645 371381
rect 396579 371316 396580 371380
rect 396644 371316 396645 371380
rect 396579 371315 396645 371316
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 355308 391574 356058
rect 397794 363454 398414 373000
rect 398974 371653 399034 374990
rect 400262 372605 400322 374990
rect 400259 372604 400325 372605
rect 400259 372540 400260 372604
rect 400324 372540 400325 372604
rect 400259 372539 400325 372540
rect 398971 371652 399037 371653
rect 398971 371588 398972 371652
rect 399036 371588 399037 371652
rect 398971 371587 399037 371588
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 355308 398414 362898
rect 401514 367174 402134 373000
rect 402286 371789 402346 374990
rect 403022 374990 403158 375050
rect 403574 374990 404246 375050
rect 404862 374990 405470 375050
rect 402283 371788 402349 371789
rect 402283 371724 402284 371788
rect 402348 371724 402349 371788
rect 402283 371723 402349 371724
rect 403022 371381 403082 374990
rect 403574 372605 403634 374990
rect 403571 372604 403637 372605
rect 403571 372540 403572 372604
rect 403636 372540 403637 372604
rect 403571 372539 403637 372540
rect 404862 372061 404922 374990
rect 405963 374988 405964 375052
rect 406028 375050 406029 375052
rect 407803 375052 407869 375053
rect 406028 374990 406558 375050
rect 407254 374990 407646 375050
rect 406028 374988 406029 374990
rect 405963 374987 406029 374988
rect 404859 372060 404925 372061
rect 404859 371996 404860 372060
rect 404924 371996 404925 372060
rect 404859 371995 404925 371996
rect 403019 371380 403085 371381
rect 403019 371316 403020 371380
rect 403084 371316 403085 371380
rect 403019 371315 403085 371316
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 355308 402134 366618
rect 405234 370894 405854 373000
rect 407254 372061 407314 374990
rect 407803 374988 407804 375052
rect 407868 375050 407869 375052
rect 425099 375052 425165 375053
rect 407868 374990 408326 375050
rect 408542 374990 408734 375050
rect 410014 374990 410094 375050
rect 407868 374988 407869 374990
rect 407803 374987 407869 374988
rect 408542 373285 408602 374990
rect 408539 373284 408605 373285
rect 408539 373220 408540 373284
rect 408604 373220 408605 373284
rect 408539 373219 408605 373220
rect 407251 372060 407317 372061
rect 407251 371996 407252 372060
rect 407316 371996 407317 372060
rect 407251 371995 407317 371996
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 355308 405854 370338
rect 408954 357554 409574 373000
rect 410014 371789 410074 374990
rect 410744 374645 410804 375020
rect 410741 374644 410807 374645
rect 410741 374580 410742 374644
rect 410806 374580 410807 374644
rect 410741 374579 410807 374580
rect 410011 371788 410077 371789
rect 410011 371724 410012 371788
rect 410076 371724 410077 371788
rect 410011 371723 410077 371724
rect 411302 371653 411362 375050
rect 411854 374990 412406 375050
rect 412774 374990 413494 375050
rect 413630 374990 413754 375050
rect 411299 371652 411365 371653
rect 411299 371588 411300 371652
rect 411364 371588 411365 371652
rect 411299 371587 411365 371588
rect 411854 371517 411914 374990
rect 411851 371516 411917 371517
rect 411851 371452 411852 371516
rect 411916 371452 411917 371516
rect 411851 371451 411917 371452
rect 412774 371381 412834 374990
rect 413694 371381 413754 374990
rect 414062 374990 414582 375050
rect 415534 374990 415942 375050
rect 416078 374990 416146 375050
rect 414062 371381 414122 374990
rect 415534 371381 415594 374990
rect 416086 374101 416146 374990
rect 416822 374990 417030 375050
rect 416083 374100 416149 374101
rect 416083 374036 416084 374100
rect 416148 374036 416149 374100
rect 416083 374035 416149 374036
rect 412771 371380 412837 371381
rect 412771 371316 412772 371380
rect 412836 371316 412837 371380
rect 412771 371315 412837 371316
rect 413691 371380 413757 371381
rect 413691 371316 413692 371380
rect 413756 371316 413757 371380
rect 413691 371315 413757 371316
rect 414059 371380 414125 371381
rect 414059 371316 414060 371380
rect 414124 371316 414125 371380
rect 414059 371315 414125 371316
rect 415531 371380 415597 371381
rect 415531 371316 415532 371380
rect 415596 371316 415597 371380
rect 415531 371315 415597 371316
rect 408954 357318 408986 357554
rect 409222 357318 409306 357554
rect 409542 357318 409574 357554
rect 408954 357234 409574 357318
rect 408954 356998 408986 357234
rect 409222 356998 409306 357234
rect 409542 356998 409574 357234
rect 408954 355308 409574 356998
rect 415794 364394 416414 373000
rect 416822 371381 416882 374990
rect 418110 371381 418170 375050
rect 418294 374990 418526 375050
rect 418846 374990 419478 375050
rect 420318 374990 420702 375050
rect 418294 373693 418354 374990
rect 418291 373692 418357 373693
rect 418291 373628 418292 373692
rect 418356 373628 418357 373692
rect 418291 373627 418357 373628
rect 418846 371517 418906 374990
rect 418843 371516 418909 371517
rect 418843 371452 418844 371516
rect 418908 371452 418909 371516
rect 418843 371451 418909 371452
rect 416819 371380 416885 371381
rect 416819 371316 416820 371380
rect 416884 371316 416885 371380
rect 416819 371315 416885 371316
rect 418107 371380 418173 371381
rect 418107 371316 418108 371380
rect 418172 371316 418173 371380
rect 418107 371315 418173 371316
rect 415794 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 416414 364394
rect 415794 364074 416414 364158
rect 415794 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 416414 364074
rect 415794 355308 416414 363838
rect 419514 366234 420134 373000
rect 420318 371381 420378 374990
rect 421054 371381 421114 375050
rect 421238 374990 421790 375050
rect 422342 374990 422878 375050
rect 423078 374990 423558 375050
rect 423966 374990 424058 375050
rect 421238 371517 421298 374990
rect 422342 372061 422402 374990
rect 423078 373693 423138 374990
rect 423075 373692 423141 373693
rect 423075 373628 423076 373692
rect 423140 373628 423141 373692
rect 423075 373627 423141 373628
rect 422339 372060 422405 372061
rect 422339 371996 422340 372060
rect 422404 371996 422405 372060
rect 422339 371995 422405 371996
rect 421235 371516 421301 371517
rect 421235 371452 421236 371516
rect 421300 371452 421301 371516
rect 421235 371451 421301 371452
rect 420315 371380 420381 371381
rect 420315 371316 420316 371380
rect 420380 371316 420381 371380
rect 420315 371315 420381 371316
rect 421051 371380 421117 371381
rect 421051 371316 421052 371380
rect 421116 371316 421117 371380
rect 421051 371315 421117 371316
rect 419514 365998 419546 366234
rect 419782 365998 419866 366234
rect 420102 365998 420134 366234
rect 419514 365914 420134 365998
rect 419514 365678 419546 365914
rect 419782 365678 419866 365914
rect 420102 365678 420134 365914
rect 419514 355308 420134 365678
rect 423234 369954 423854 373000
rect 423998 371517 424058 374990
rect 425099 374988 425100 375052
rect 425164 375050 425165 375052
rect 440371 375052 440437 375053
rect 425164 374990 425326 375050
rect 425654 374990 426006 375050
rect 425164 374988 425165 374990
rect 425099 374987 425165 374988
rect 423995 371516 424061 371517
rect 423995 371452 423996 371516
rect 424060 371452 424061 371516
rect 423995 371451 424061 371452
rect 425654 371381 425714 374990
rect 426390 371517 426450 375050
rect 426942 374990 427638 375050
rect 427862 374990 428318 375050
rect 428598 374990 428726 375050
rect 429334 374990 429814 375050
rect 430622 374990 431038 375050
rect 426942 373693 427002 374990
rect 426939 373692 427005 373693
rect 426939 373628 426940 373692
rect 427004 373628 427005 373692
rect 426939 373627 427005 373628
rect 427862 373557 427922 374990
rect 427859 373556 427925 373557
rect 427859 373492 427860 373556
rect 427924 373492 427925 373556
rect 427859 373491 427925 373492
rect 426387 371516 426453 371517
rect 426387 371452 426388 371516
rect 426452 371452 426453 371516
rect 426387 371451 426453 371452
rect 425651 371380 425717 371381
rect 425651 371316 425652 371380
rect 425716 371316 425717 371380
rect 425651 371315 425717 371316
rect 423234 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 423854 369954
rect 423234 369634 423854 369718
rect 423234 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 423854 369634
rect 423234 355308 423854 369398
rect 426954 356614 427574 373000
rect 428598 371381 428658 374990
rect 429334 371381 429394 374990
rect 430622 371381 430682 374990
rect 431174 371517 431234 375050
rect 432094 374990 432262 375050
rect 431171 371516 431237 371517
rect 431171 371452 431172 371516
rect 431236 371452 431237 371516
rect 431171 371451 431237 371452
rect 432094 371381 432154 374990
rect 433320 374370 433380 375020
rect 433592 374509 433652 375020
rect 433750 374990 434438 375050
rect 434854 374990 435798 375050
rect 433589 374508 433655 374509
rect 433589 374444 433590 374508
rect 433654 374444 433655 374508
rect 433589 374443 433655 374444
rect 433320 374310 433442 374370
rect 433382 371381 433442 374310
rect 433750 374010 433810 374990
rect 433566 373950 433810 374010
rect 433566 372469 433626 373950
rect 433563 372468 433629 372469
rect 433563 372404 433564 372468
rect 433628 372404 433629 372468
rect 433563 372403 433629 372404
rect 428595 371380 428661 371381
rect 428595 371316 428596 371380
rect 428660 371316 428661 371380
rect 428595 371315 428661 371316
rect 429331 371380 429397 371381
rect 429331 371316 429332 371380
rect 429396 371316 429397 371380
rect 429331 371315 429397 371316
rect 430619 371380 430685 371381
rect 430619 371316 430620 371380
rect 430684 371316 430685 371380
rect 430619 371315 430685 371316
rect 432091 371380 432157 371381
rect 432091 371316 432092 371380
rect 432156 371316 432157 371380
rect 432091 371315 432157 371316
rect 433379 371380 433445 371381
rect 433379 371316 433380 371380
rect 433444 371316 433445 371380
rect 433379 371315 433445 371316
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 355308 427574 356058
rect 433794 363454 434414 373000
rect 434854 371381 434914 374990
rect 436040 374509 436100 375020
rect 436326 374990 437022 375050
rect 438110 374990 438410 375050
rect 436037 374508 436103 374509
rect 436037 374444 436038 374508
rect 436102 374444 436103 374508
rect 436037 374443 436103 374444
rect 436326 371381 436386 374990
rect 434851 371380 434917 371381
rect 434851 371316 434852 371380
rect 434916 371316 434917 371380
rect 434851 371315 434917 371316
rect 436323 371380 436389 371381
rect 436323 371316 436324 371380
rect 436388 371316 436389 371380
rect 436323 371315 436389 371316
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 355308 434414 362898
rect 437514 367174 438134 373000
rect 438350 371925 438410 374990
rect 438488 374509 438548 375020
rect 438902 374990 439198 375050
rect 438485 374508 438551 374509
rect 438485 374444 438486 374508
rect 438550 374444 438551 374508
rect 438485 374443 438551 374444
rect 438902 372333 438962 374990
rect 440371 374988 440372 375052
rect 440436 375050 440437 375052
rect 443131 375052 443197 375053
rect 440436 374990 440966 375050
rect 440436 374988 440437 374990
rect 440371 374987 440437 374988
rect 443131 374988 443132 375052
rect 443196 375050 443197 375052
rect 452883 375052 452949 375053
rect 443196 374990 443550 375050
rect 445894 374990 445998 375050
rect 447734 374990 448310 375050
rect 450310 374990 451030 375050
rect 443196 374988 443197 374990
rect 443131 374987 443197 374988
rect 445894 373693 445954 374990
rect 445891 373692 445957 373693
rect 445891 373628 445892 373692
rect 445956 373628 445957 373692
rect 445891 373627 445957 373628
rect 447734 373421 447794 374990
rect 450310 373557 450370 374990
rect 452883 374988 452884 375052
rect 452948 375050 452949 375052
rect 452948 374990 453478 375050
rect 455462 374990 455926 375050
rect 458222 374990 458510 375050
rect 460958 374990 461042 375050
rect 452948 374988 452949 374990
rect 452883 374987 452949 374988
rect 455462 373557 455522 374990
rect 450307 373556 450373 373557
rect 450307 373492 450308 373556
rect 450372 373492 450373 373556
rect 450307 373491 450373 373492
rect 455459 373556 455525 373557
rect 455459 373492 455460 373556
rect 455524 373492 455525 373556
rect 455459 373491 455525 373492
rect 447731 373420 447797 373421
rect 447731 373356 447732 373420
rect 447796 373356 447797 373420
rect 447731 373355 447797 373356
rect 438899 372332 438965 372333
rect 438899 372268 438900 372332
rect 438964 372268 438965 372332
rect 438899 372267 438965 372268
rect 438347 371924 438413 371925
rect 438347 371860 438348 371924
rect 438412 371860 438413 371924
rect 438347 371859 438413 371860
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 355308 438134 366618
rect 441234 370894 441854 373000
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 355308 441854 370338
rect 444954 357554 445574 373000
rect 444954 357318 444986 357554
rect 445222 357318 445306 357554
rect 445542 357318 445574 357554
rect 444954 357234 445574 357318
rect 444954 356998 444986 357234
rect 445222 356998 445306 357234
rect 445542 356998 445574 357234
rect 444954 355308 445574 356998
rect 451794 364394 452414 373000
rect 451794 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 452414 364394
rect 451794 364074 452414 364158
rect 451794 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 452414 364074
rect 451794 355308 452414 363838
rect 455514 366234 456134 373000
rect 458222 371381 458282 374990
rect 460982 373829 461042 374990
rect 462822 374990 463542 375050
rect 465398 374990 465990 375050
rect 467974 374990 468574 375050
rect 470734 374990 471022 375050
rect 473310 374990 473470 375050
rect 475334 374990 475918 375050
rect 478094 374990 478502 375050
rect 480302 374990 480950 375050
rect 483246 374990 483398 375050
rect 485822 374990 485982 375050
rect 503118 374990 503254 375050
rect 503390 374990 503546 375050
rect 460979 373828 461045 373829
rect 460979 373764 460980 373828
rect 461044 373764 461045 373828
rect 460979 373763 461045 373764
rect 462822 373421 462882 374990
rect 462819 373420 462885 373421
rect 462819 373356 462820 373420
rect 462884 373356 462885 373420
rect 462819 373355 462885 373356
rect 458219 371380 458285 371381
rect 458219 371316 458220 371380
rect 458284 371316 458285 371380
rect 458219 371315 458285 371316
rect 455514 365998 455546 366234
rect 455782 365998 455866 366234
rect 456102 365998 456134 366234
rect 455514 365914 456134 365998
rect 455514 365678 455546 365914
rect 455782 365678 455866 365914
rect 456102 365678 456134 365914
rect 455514 355308 456134 365678
rect 459234 369954 459854 373000
rect 459234 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 459854 369954
rect 459234 369634 459854 369718
rect 459234 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 459854 369634
rect 459234 355308 459854 369398
rect 462954 356614 463574 373000
rect 465398 371653 465458 374990
rect 465395 371652 465461 371653
rect 465395 371588 465396 371652
rect 465460 371588 465461 371652
rect 465395 371587 465461 371588
rect 467974 371245 468034 374990
rect 467971 371244 468037 371245
rect 467971 371180 467972 371244
rect 468036 371180 468037 371244
rect 467971 371179 468037 371180
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 355308 463574 356058
rect 469794 363454 470414 373000
rect 470734 372333 470794 374990
rect 470731 372332 470797 372333
rect 470731 372268 470732 372332
rect 470796 372268 470797 372332
rect 470731 372267 470797 372268
rect 473310 371381 473370 374990
rect 473307 371380 473373 371381
rect 473307 371316 473308 371380
rect 473372 371316 473373 371380
rect 473307 371315 473373 371316
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 355308 470414 362898
rect 473514 367174 474134 373000
rect 475334 371381 475394 374990
rect 475331 371380 475397 371381
rect 475331 371316 475332 371380
rect 475396 371316 475397 371380
rect 475331 371315 475397 371316
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 355308 474134 366618
rect 477234 370894 477854 373000
rect 478094 371381 478154 374990
rect 480302 371381 480362 374990
rect 478091 371380 478157 371381
rect 478091 371316 478092 371380
rect 478156 371316 478157 371380
rect 478091 371315 478157 371316
rect 480299 371380 480365 371381
rect 480299 371316 480300 371380
rect 480364 371316 480365 371380
rect 480299 371315 480365 371316
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 355308 477854 370338
rect 480954 357554 481574 373000
rect 483246 371925 483306 374990
rect 485822 373965 485882 374990
rect 485819 373964 485885 373965
rect 485819 373900 485820 373964
rect 485884 373900 485885 373964
rect 485819 373899 485885 373900
rect 483243 371924 483309 371925
rect 483243 371860 483244 371924
rect 483308 371860 483309 371924
rect 483243 371859 483309 371860
rect 480954 357318 480986 357554
rect 481222 357318 481306 357554
rect 481542 357318 481574 357554
rect 480954 357234 481574 357318
rect 480954 356998 480986 357234
rect 481222 356998 481306 357234
rect 481542 356998 481574 357234
rect 480954 355308 481574 356998
rect 487794 364394 488414 373000
rect 487794 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 487794 364074 488414 364158
rect 487794 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 487794 355308 488414 363838
rect 491514 366234 492134 373000
rect 491514 365998 491546 366234
rect 491782 365998 491866 366234
rect 492102 365998 492134 366234
rect 491514 365914 492134 365998
rect 491514 365678 491546 365914
rect 491782 365678 491866 365914
rect 492102 365678 492134 365914
rect 491514 355308 492134 365678
rect 495234 369954 495854 373000
rect 495234 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 495234 369634 495854 369718
rect 495234 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 495234 355308 495854 369398
rect 498954 356614 499574 373000
rect 503118 372197 503178 374990
rect 503486 372197 503546 374990
rect 503115 372196 503181 372197
rect 503115 372132 503116 372196
rect 503180 372132 503181 372196
rect 503115 372131 503181 372132
rect 503483 372196 503549 372197
rect 503483 372132 503484 372196
rect 503548 372132 503549 372196
rect 503483 372131 503549 372132
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 355308 499574 356058
rect 505794 363454 506414 373000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 355308 506414 362898
rect 509514 367174 510134 373000
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 355308 510134 366618
rect 513234 370894 513854 373000
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 355308 513854 370338
rect 516954 357554 517574 373000
rect 516954 357318 516986 357554
rect 517222 357318 517306 357554
rect 517542 357318 517574 357554
rect 516954 357234 517574 357318
rect 516954 356998 516986 357234
rect 517222 356998 517306 357234
rect 517542 356998 517574 357234
rect 516954 355308 517574 356998
rect 498515 355060 498581 355061
rect 498515 354996 498516 355060
rect 498580 354996 498581 355060
rect 498515 354995 498581 354996
rect 498518 353970 498578 354995
rect 499803 354924 499869 354925
rect 499803 354860 499804 354924
rect 499868 354860 499869 354924
rect 499803 354859 499869 354860
rect 499806 353970 499866 354859
rect 510843 354788 510909 354789
rect 510843 354724 510844 354788
rect 510908 354724 510909 354788
rect 510843 354723 510909 354724
rect 510846 353970 510906 354723
rect 498464 353910 498578 353970
rect 499688 353910 499866 353970
rect 510840 353910 510906 353970
rect 498464 353260 498524 353910
rect 499688 353260 499748 353910
rect 510840 353260 510900 353910
rect 380272 345454 380620 345486
rect 380272 345218 380328 345454
rect 380564 345218 380620 345454
rect 380272 345134 380620 345218
rect 380272 344898 380328 345134
rect 380564 344898 380620 345134
rect 380272 344866 380620 344898
rect 516000 345454 516348 345486
rect 516000 345218 516056 345454
rect 516292 345218 516348 345454
rect 516000 345134 516348 345218
rect 516000 344898 516056 345134
rect 516292 344898 516348 345134
rect 516000 344866 516348 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 380952 327454 381300 327486
rect 380952 327218 381008 327454
rect 381244 327218 381300 327454
rect 380952 327134 381300 327218
rect 380952 326898 381008 327134
rect 381244 326898 381300 327134
rect 380952 326866 381300 326898
rect 515320 327454 515668 327486
rect 515320 327218 515376 327454
rect 515612 327218 515668 327454
rect 515320 327134 515668 327218
rect 515320 326898 515376 327134
rect 515612 326898 515668 327134
rect 515320 326866 515668 326898
rect 380272 309454 380620 309486
rect 380272 309218 380328 309454
rect 380564 309218 380620 309454
rect 380272 309134 380620 309218
rect 380272 308898 380328 309134
rect 380564 308898 380620 309134
rect 380272 308866 380620 308898
rect 516000 309454 516348 309486
rect 516000 309218 516056 309454
rect 516292 309218 516348 309454
rect 516000 309134 516348 309218
rect 516000 308898 516056 309134
rect 516292 308898 516348 309134
rect 516000 308866 516348 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 380952 291454 381300 291486
rect 380952 291218 381008 291454
rect 381244 291218 381300 291454
rect 380952 291134 381300 291218
rect 380952 290898 381008 291134
rect 381244 290898 381300 291134
rect 380952 290866 381300 290898
rect 515320 291454 515668 291486
rect 515320 291218 515376 291454
rect 515612 291218 515668 291454
rect 515320 291134 515668 291218
rect 515320 290898 515376 291134
rect 515612 290898 515668 291134
rect 515320 290866 515668 290898
rect 380272 273454 380620 273486
rect 380272 273218 380328 273454
rect 380564 273218 380620 273454
rect 380272 273134 380620 273218
rect 380272 272898 380328 273134
rect 380564 272898 380620 273134
rect 380272 272866 380620 272898
rect 516000 273454 516348 273486
rect 516000 273218 516056 273454
rect 516292 273218 516348 273454
rect 516000 273134 516348 273218
rect 516000 272898 516056 273134
rect 516292 272898 516348 273134
rect 516000 272866 516348 272898
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 396056 269650 396116 270106
rect 397144 269650 397204 270106
rect 396056 269590 396274 269650
rect 379470 267690 379714 267750
rect 379470 267341 379530 267690
rect 379467 267340 379533 267341
rect 379467 267276 379468 267340
rect 379532 267276 379533 267340
rect 379467 267275 379533 267276
rect 379794 256394 380414 268000
rect 379794 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 380414 256394
rect 379794 256074 380414 256158
rect 379794 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 380414 256074
rect 379794 250308 380414 255838
rect 383514 260114 384134 268000
rect 383514 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 384134 260114
rect 383514 259794 384134 259878
rect 383514 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 384134 259794
rect 383514 250308 384134 259558
rect 387234 261954 387854 268000
rect 387234 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 387854 261954
rect 387234 261634 387854 261718
rect 387234 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 387854 261634
rect 387234 250308 387854 261398
rect 390954 265674 391574 268000
rect 396214 267069 396274 269590
rect 397134 269590 397204 269650
rect 398232 269650 398292 270106
rect 399592 269650 399652 270106
rect 400544 269650 400604 270106
rect 401768 269650 401828 270106
rect 403128 269650 403188 270106
rect 404216 269650 404276 270106
rect 405440 269650 405500 270106
rect 406528 269650 406588 270106
rect 398232 269590 398298 269650
rect 397134 267205 397194 269590
rect 398238 268157 398298 269590
rect 399526 269590 399652 269650
rect 400446 269590 400604 269650
rect 401734 269590 401828 269650
rect 403022 269590 403188 269650
rect 404126 269590 404276 269650
rect 405046 269590 405500 269650
rect 406518 269590 406588 269650
rect 407616 269650 407676 270106
rect 408296 269650 408356 270106
rect 407616 269590 407682 269650
rect 398235 268156 398301 268157
rect 398235 268092 398236 268156
rect 398300 268092 398301 268156
rect 398235 268091 398301 268092
rect 397131 267204 397197 267205
rect 397131 267140 397132 267204
rect 397196 267140 397197 267204
rect 397131 267139 397197 267140
rect 396211 267068 396277 267069
rect 396211 267004 396212 267068
rect 396276 267004 396277 267068
rect 396211 267003 396277 267004
rect 390954 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 391574 265674
rect 390954 265354 391574 265438
rect 390954 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 391574 265354
rect 390954 250308 391574 265118
rect 397794 255454 398414 268000
rect 399526 266389 399586 269590
rect 400446 266389 400506 269590
rect 401734 268157 401794 269590
rect 401731 268156 401797 268157
rect 401731 268092 401732 268156
rect 401796 268092 401797 268156
rect 401731 268091 401797 268092
rect 399523 266388 399589 266389
rect 399523 266324 399524 266388
rect 399588 266324 399589 266388
rect 399523 266323 399589 266324
rect 400443 266388 400509 266389
rect 400443 266324 400444 266388
rect 400508 266324 400509 266388
rect 400443 266323 400509 266324
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 250308 398414 254898
rect 401514 259174 402134 268000
rect 403022 267749 403082 269590
rect 403019 267748 403085 267749
rect 403019 267684 403020 267748
rect 403084 267684 403085 267748
rect 403019 267683 403085 267684
rect 404126 266389 404186 269590
rect 405046 266389 405106 269590
rect 404123 266388 404189 266389
rect 404123 266324 404124 266388
rect 404188 266324 404189 266388
rect 404123 266323 404189 266324
rect 405043 266388 405109 266389
rect 405043 266324 405044 266388
rect 405108 266324 405109 266388
rect 405043 266323 405109 266324
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 250308 402134 258618
rect 405234 262894 405854 268000
rect 406518 266389 406578 269590
rect 407622 266389 407682 269590
rect 408174 269590 408356 269650
rect 408704 269650 408764 270106
rect 410064 269650 410124 270106
rect 408704 269590 408786 269650
rect 408174 267069 408234 269590
rect 408171 267068 408237 267069
rect 408171 267004 408172 267068
rect 408236 267004 408237 267068
rect 408171 267003 408237 267004
rect 408726 266389 408786 269590
rect 410014 269590 410124 269650
rect 410744 269650 410804 270106
rect 411288 269650 411348 270106
rect 412376 269650 412436 270106
rect 413464 269650 413524 270106
rect 410744 269590 410810 269650
rect 411288 269590 411362 269650
rect 412376 269590 412466 269650
rect 408954 266614 409574 268000
rect 406515 266388 406581 266389
rect 406515 266324 406516 266388
rect 406580 266324 406581 266388
rect 406515 266323 406581 266324
rect 407619 266388 407685 266389
rect 407619 266324 407620 266388
rect 407684 266324 407685 266388
rect 407619 266323 407685 266324
rect 408723 266388 408789 266389
rect 408723 266324 408724 266388
rect 408788 266324 408789 266388
rect 408723 266323 408789 266324
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 410014 266389 410074 269590
rect 410750 267069 410810 269590
rect 410747 267068 410813 267069
rect 410747 267004 410748 267068
rect 410812 267004 410813 267068
rect 410747 267003 410813 267004
rect 411302 266389 411362 269590
rect 412406 266525 412466 269590
rect 413326 269590 413524 269650
rect 413600 269650 413660 270106
rect 414552 269650 414612 270106
rect 415912 269650 415972 270106
rect 413600 269590 413754 269650
rect 412403 266524 412469 266525
rect 412403 266460 412404 266524
rect 412468 266460 412469 266524
rect 412403 266459 412469 266460
rect 413326 266389 413386 269590
rect 413694 267069 413754 269590
rect 414430 269590 414612 269650
rect 415902 269590 415972 269650
rect 416048 269650 416108 270106
rect 417000 269650 417060 270106
rect 418088 269650 418148 270106
rect 418496 269789 418556 270106
rect 418493 269788 418559 269789
rect 418493 269724 418494 269788
rect 418558 269724 418559 269788
rect 418493 269723 418559 269724
rect 419448 269650 419508 270106
rect 416048 269590 416146 269650
rect 417000 269590 417066 269650
rect 418088 269590 418170 269650
rect 414430 267749 414490 269590
rect 415902 268837 415962 269590
rect 415899 268836 415965 268837
rect 415899 268772 415900 268836
rect 415964 268772 415965 268836
rect 415899 268771 415965 268772
rect 416086 268157 416146 269590
rect 416083 268156 416149 268157
rect 416083 268092 416084 268156
rect 416148 268092 416149 268156
rect 416083 268091 416149 268092
rect 414427 267748 414493 267749
rect 414427 267684 414428 267748
rect 414492 267684 414493 267748
rect 414427 267683 414493 267684
rect 413691 267068 413757 267069
rect 413691 267004 413692 267068
rect 413756 267004 413757 267068
rect 413691 267003 413757 267004
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 250308 405854 262338
rect 408954 266294 409574 266378
rect 410011 266388 410077 266389
rect 410011 266324 410012 266388
rect 410076 266324 410077 266388
rect 410011 266323 410077 266324
rect 411299 266388 411365 266389
rect 411299 266324 411300 266388
rect 411364 266324 411365 266388
rect 411299 266323 411365 266324
rect 413323 266388 413389 266389
rect 413323 266324 413324 266388
rect 413388 266324 413389 266388
rect 413323 266323 413389 266324
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 250308 409574 266058
rect 415794 256394 416414 268000
rect 417006 266389 417066 269590
rect 418110 266389 418170 269590
rect 419214 269590 419508 269650
rect 420672 269650 420732 270106
rect 421080 269650 421140 270106
rect 420672 269590 420746 269650
rect 419214 266525 419274 269590
rect 419211 266524 419277 266525
rect 419211 266460 419212 266524
rect 419276 266460 419277 266524
rect 419211 266459 419277 266460
rect 417003 266388 417069 266389
rect 417003 266324 417004 266388
rect 417068 266324 417069 266388
rect 417003 266323 417069 266324
rect 418107 266388 418173 266389
rect 418107 266324 418108 266388
rect 418172 266324 418173 266388
rect 418107 266323 418173 266324
rect 415794 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 416414 256394
rect 415794 256074 416414 256158
rect 415794 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 416414 256074
rect 415794 250308 416414 255838
rect 419514 260114 420134 268000
rect 420686 266389 420746 269590
rect 421054 269590 421140 269650
rect 421760 269650 421820 270106
rect 422848 269650 422908 270106
rect 423528 269653 423588 270106
rect 423525 269652 423591 269653
rect 421760 269590 421850 269650
rect 422848 269590 422954 269650
rect 421054 268837 421114 269590
rect 421051 268836 421117 268837
rect 421051 268772 421052 268836
rect 421116 268772 421117 268836
rect 421051 268771 421117 268772
rect 421790 266389 421850 269590
rect 422894 267069 422954 269590
rect 423525 269588 423526 269652
rect 423590 269588 423591 269652
rect 423936 269650 423996 270106
rect 425296 269789 425356 270106
rect 425293 269788 425359 269789
rect 425293 269724 425294 269788
rect 425358 269724 425359 269788
rect 425293 269723 425359 269724
rect 425976 269650 426036 270106
rect 426384 269653 426444 270106
rect 426384 269652 426453 269653
rect 423936 269590 424058 269650
rect 425976 269590 426082 269650
rect 426384 269590 426388 269652
rect 423525 269587 423591 269588
rect 423998 268701 424058 269590
rect 426022 268973 426082 269590
rect 426387 269588 426388 269590
rect 426452 269588 426453 269652
rect 427608 269650 427668 270106
rect 428288 269650 428348 270106
rect 427608 269590 427738 269650
rect 426387 269587 426453 269588
rect 426019 268972 426085 268973
rect 426019 268908 426020 268972
rect 426084 268908 426085 268972
rect 426019 268907 426085 268908
rect 423995 268700 424061 268701
rect 423995 268636 423996 268700
rect 424060 268636 424061 268700
rect 423995 268635 424061 268636
rect 422891 267068 422957 267069
rect 422891 267004 422892 267068
rect 422956 267004 422957 267068
rect 422891 267003 422957 267004
rect 420683 266388 420749 266389
rect 420683 266324 420684 266388
rect 420748 266324 420749 266388
rect 420683 266323 420749 266324
rect 421787 266388 421853 266389
rect 421787 266324 421788 266388
rect 421852 266324 421853 266388
rect 421787 266323 421853 266324
rect 419514 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 420134 260114
rect 419514 259794 420134 259878
rect 419514 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 420134 259794
rect 419514 250308 420134 259558
rect 423234 261954 423854 268000
rect 423234 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 423854 261954
rect 423234 261634 423854 261718
rect 423234 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 423854 261634
rect 423234 250308 423854 261398
rect 426954 265674 427574 268000
rect 426954 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 427574 265674
rect 427678 265573 427738 269590
rect 428230 269590 428348 269650
rect 428696 269650 428756 270106
rect 429784 269650 429844 270106
rect 431008 269650 431068 270106
rect 428696 269590 428842 269650
rect 429784 269590 429946 269650
rect 428230 267341 428290 269590
rect 428227 267340 428293 267341
rect 428227 267276 428228 267340
rect 428292 267276 428293 267340
rect 428227 267275 428293 267276
rect 428782 266389 428842 269590
rect 429886 266389 429946 269590
rect 430990 269590 431068 269650
rect 431144 269650 431204 270106
rect 432232 269650 432292 270106
rect 433320 269650 433380 270106
rect 433592 269653 433652 270106
rect 433589 269652 433655 269653
rect 431144 269590 431234 269650
rect 432232 269590 432338 269650
rect 433320 269590 433442 269650
rect 430990 268973 431050 269590
rect 430987 268972 431053 268973
rect 430987 268908 430988 268972
rect 431052 268908 431053 268972
rect 430987 268907 431053 268908
rect 431174 266389 431234 269590
rect 432278 267749 432338 269590
rect 433382 268973 433442 269590
rect 433589 269588 433590 269652
rect 433654 269588 433655 269652
rect 434408 269650 434468 270106
rect 433589 269587 433655 269588
rect 434302 269590 434468 269650
rect 435768 269650 435828 270106
rect 436040 269650 436100 270106
rect 436992 269650 437052 270106
rect 435768 269590 435834 269650
rect 433379 268972 433445 268973
rect 433379 268908 433380 268972
rect 433444 268908 433445 268972
rect 433379 268907 433445 268908
rect 434302 268157 434362 269590
rect 434299 268156 434365 268157
rect 434299 268092 434300 268156
rect 434364 268092 434365 268156
rect 434299 268091 434365 268092
rect 432275 267748 432341 267749
rect 432275 267684 432276 267748
rect 432340 267684 432341 267748
rect 432275 267683 432341 267684
rect 428779 266388 428845 266389
rect 428779 266324 428780 266388
rect 428844 266324 428845 266388
rect 428779 266323 428845 266324
rect 429883 266388 429949 266389
rect 429883 266324 429884 266388
rect 429948 266324 429949 266388
rect 429883 266323 429949 266324
rect 431171 266388 431237 266389
rect 431171 266324 431172 266388
rect 431236 266324 431237 266388
rect 431171 266323 431237 266324
rect 427675 265572 427741 265573
rect 427675 265508 427676 265572
rect 427740 265508 427741 265572
rect 427675 265507 427741 265508
rect 426954 265354 427574 265438
rect 426954 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 427574 265354
rect 426954 250308 427574 265118
rect 433794 255454 434414 268000
rect 435774 267749 435834 269590
rect 435958 269590 436100 269650
rect 436878 269590 437052 269650
rect 438080 269650 438140 270106
rect 438488 269650 438548 270106
rect 439168 269650 439228 270106
rect 440936 269650 440996 270106
rect 443520 269650 443580 270106
rect 445968 269650 446028 270106
rect 438080 269590 438410 269650
rect 438488 269590 438594 269650
rect 435958 267749 436018 269590
rect 435771 267748 435837 267749
rect 435771 267684 435772 267748
rect 435836 267684 435837 267748
rect 435771 267683 435837 267684
rect 435955 267748 436021 267749
rect 435955 267684 435956 267748
rect 436020 267684 436021 267748
rect 435955 267683 436021 267684
rect 436878 266389 436938 269590
rect 436875 266388 436941 266389
rect 436875 266324 436876 266388
rect 436940 266324 436941 266388
rect 436875 266323 436941 266324
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 250308 434414 254898
rect 437514 259174 438134 268000
rect 438350 266389 438410 269590
rect 438534 267341 438594 269590
rect 439086 269590 439228 269650
rect 440926 269590 440996 269650
rect 443502 269590 443580 269650
rect 445894 269590 446028 269650
rect 448280 269650 448340 270106
rect 451000 269650 451060 270106
rect 453448 269653 453508 270106
rect 453445 269652 453511 269653
rect 448280 269590 448346 269650
rect 451000 269590 451106 269650
rect 438531 267340 438597 267341
rect 438531 267276 438532 267340
rect 438596 267276 438597 267340
rect 438531 267275 438597 267276
rect 439086 266389 439146 269590
rect 440926 267205 440986 269590
rect 440923 267204 440989 267205
rect 440923 267140 440924 267204
rect 440988 267140 440989 267204
rect 440923 267139 440989 267140
rect 438347 266388 438413 266389
rect 438347 266324 438348 266388
rect 438412 266324 438413 266388
rect 438347 266323 438413 266324
rect 439083 266388 439149 266389
rect 439083 266324 439084 266388
rect 439148 266324 439149 266388
rect 439083 266323 439149 266324
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 250308 438134 258618
rect 441234 262894 441854 268000
rect 443502 267341 443562 269590
rect 443499 267340 443565 267341
rect 443499 267276 443500 267340
rect 443564 267276 443565 267340
rect 443499 267275 443565 267276
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 250308 441854 262338
rect 444954 266614 445574 268000
rect 445894 267749 445954 269590
rect 448286 267749 448346 269590
rect 451046 267749 451106 269590
rect 453445 269588 453446 269652
rect 453510 269588 453511 269652
rect 455896 269650 455956 270106
rect 458480 269650 458540 270106
rect 453445 269587 453511 269588
rect 455830 269590 455956 269650
rect 458406 269590 458540 269650
rect 460928 269650 460988 270106
rect 463512 269650 463572 270106
rect 465960 269650 466020 270106
rect 468544 269653 468604 270106
rect 460928 269590 461042 269650
rect 455830 268157 455890 269590
rect 455827 268156 455893 268157
rect 455827 268092 455828 268156
rect 455892 268092 455893 268156
rect 455827 268091 455893 268092
rect 445891 267748 445957 267749
rect 445891 267684 445892 267748
rect 445956 267684 445957 267748
rect 445891 267683 445957 267684
rect 448283 267748 448349 267749
rect 448283 267684 448284 267748
rect 448348 267684 448349 267748
rect 448283 267683 448349 267684
rect 451043 267748 451109 267749
rect 451043 267684 451044 267748
rect 451108 267684 451109 267748
rect 451043 267683 451109 267684
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 250308 445574 266058
rect 451794 256394 452414 268000
rect 451794 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 452414 256394
rect 451794 256074 452414 256158
rect 451794 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 452414 256074
rect 451794 250308 452414 255838
rect 455514 260114 456134 268000
rect 458406 267749 458466 269590
rect 458403 267748 458469 267749
rect 458403 267684 458404 267748
rect 458468 267684 458469 267748
rect 458403 267683 458469 267684
rect 455514 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 456134 260114
rect 455514 259794 456134 259878
rect 455514 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 456134 259794
rect 455514 250308 456134 259558
rect 459234 261954 459854 268000
rect 460982 267477 461042 269590
rect 462638 269590 463572 269650
rect 465950 269590 466020 269650
rect 468541 269652 468607 269653
rect 460979 267476 461045 267477
rect 460979 267412 460980 267476
rect 461044 267412 461045 267476
rect 460979 267411 461045 267412
rect 462638 266933 462698 269590
rect 462635 266932 462701 266933
rect 462635 266868 462636 266932
rect 462700 266868 462701 266932
rect 462635 266867 462701 266868
rect 459234 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 459854 261954
rect 459234 261634 459854 261718
rect 459234 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 459854 261634
rect 459234 250308 459854 261398
rect 462954 265674 463574 268000
rect 465950 267613 466010 269590
rect 468541 269588 468542 269652
rect 468606 269588 468607 269652
rect 470992 269650 471052 270106
rect 473440 269650 473500 270106
rect 475888 269650 475948 270106
rect 478472 269650 478532 270106
rect 480920 269653 480980 270106
rect 468541 269587 468607 269588
rect 470918 269590 471052 269650
rect 473310 269590 473500 269650
rect 475886 269590 475948 269650
rect 478462 269590 478532 269650
rect 480917 269652 480983 269653
rect 470918 269245 470978 269590
rect 470915 269244 470981 269245
rect 470915 269180 470916 269244
rect 470980 269180 470981 269244
rect 470915 269179 470981 269180
rect 465947 267612 466013 267613
rect 465947 267548 465948 267612
rect 466012 267548 466013 267612
rect 465947 267547 466013 267548
rect 462954 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 463574 265674
rect 462954 265354 463574 265438
rect 462954 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 463574 265354
rect 462954 250308 463574 265118
rect 469794 255454 470414 268000
rect 473310 267749 473370 269590
rect 475886 268973 475946 269590
rect 478462 268973 478522 269590
rect 480917 269588 480918 269652
rect 480982 269588 480983 269652
rect 483368 269650 483428 270106
rect 485952 269650 486012 270106
rect 503224 269650 503284 270106
rect 483368 269590 483490 269650
rect 485952 269590 486066 269650
rect 480917 269587 480983 269588
rect 483430 268973 483490 269590
rect 486006 269109 486066 269590
rect 503118 269590 503284 269650
rect 503360 269650 503420 270106
rect 503360 269590 503546 269650
rect 486003 269108 486069 269109
rect 486003 269044 486004 269108
rect 486068 269044 486069 269108
rect 486003 269043 486069 269044
rect 475883 268972 475949 268973
rect 475883 268908 475884 268972
rect 475948 268908 475949 268972
rect 475883 268907 475949 268908
rect 478459 268972 478525 268973
rect 478459 268908 478460 268972
rect 478524 268908 478525 268972
rect 478459 268907 478525 268908
rect 483427 268972 483493 268973
rect 483427 268908 483428 268972
rect 483492 268908 483493 268972
rect 483427 268907 483493 268908
rect 473307 267748 473373 267749
rect 473307 267684 473308 267748
rect 473372 267684 473373 267748
rect 473307 267683 473373 267684
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 250308 470414 254898
rect 473514 259174 474134 268000
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 250308 474134 258618
rect 477234 262894 477854 268000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 250308 477854 262338
rect 480954 266614 481574 268000
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 250308 481574 266058
rect 487794 256394 488414 268000
rect 487794 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 487794 256074 488414 256158
rect 487794 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 487794 250308 488414 255838
rect 491514 260114 492134 268000
rect 491514 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 491514 259794 492134 259878
rect 491514 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 491514 250308 492134 259558
rect 495234 261954 495854 268000
rect 495234 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 495234 261634 495854 261718
rect 495234 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 495234 250308 495854 261398
rect 498954 265674 499574 268000
rect 503118 267341 503178 269590
rect 503486 267477 503546 269590
rect 503483 267476 503549 267477
rect 503483 267412 503484 267476
rect 503548 267412 503549 267476
rect 503483 267411 503549 267412
rect 503115 267340 503181 267341
rect 503115 267276 503116 267340
rect 503180 267276 503181 267340
rect 503115 267275 503181 267276
rect 498954 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 498954 265354 499574 265438
rect 498954 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 498954 250308 499574 265118
rect 505794 255454 506414 268000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 250308 506414 254898
rect 509514 259174 510134 268000
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 250308 510134 258618
rect 513234 262894 513854 268000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 250308 513854 262338
rect 516954 266614 517574 268000
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 250308 517574 266058
rect 498515 249932 498581 249933
rect 498515 249868 498516 249932
rect 498580 249868 498581 249932
rect 498515 249867 498581 249868
rect 499803 249932 499869 249933
rect 499803 249868 499804 249932
rect 499868 249868 499869 249932
rect 499803 249867 499869 249868
rect 510843 249932 510909 249933
rect 510843 249868 510844 249932
rect 510908 249868 510909 249932
rect 510843 249867 510909 249868
rect 498518 248430 498578 249867
rect 499806 248430 499866 249867
rect 510846 248430 510906 249867
rect 498464 248370 498578 248430
rect 499688 248370 499866 248430
rect 510840 248370 510906 248430
rect 498464 248202 498524 248370
rect 499688 248202 499748 248370
rect 510840 248202 510900 248370
rect 380272 237454 380620 237486
rect 380272 237218 380328 237454
rect 380564 237218 380620 237454
rect 380272 237134 380620 237218
rect 380272 236898 380328 237134
rect 380564 236898 380620 237134
rect 380272 236866 380620 236898
rect 516000 237454 516348 237486
rect 516000 237218 516056 237454
rect 516292 237218 516348 237454
rect 516000 237134 516348 237218
rect 516000 236898 516056 237134
rect 516292 236898 516348 237134
rect 516000 236866 516348 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 380952 219454 381300 219486
rect 380952 219218 381008 219454
rect 381244 219218 381300 219454
rect 380952 219134 381300 219218
rect 380952 218898 381008 219134
rect 381244 218898 381300 219134
rect 380952 218866 381300 218898
rect 515320 219454 515668 219486
rect 515320 219218 515376 219454
rect 515612 219218 515668 219454
rect 515320 219134 515668 219218
rect 515320 218898 515376 219134
rect 515612 218898 515668 219134
rect 515320 218866 515668 218898
rect 380272 201454 380620 201486
rect 380272 201218 380328 201454
rect 380564 201218 380620 201454
rect 380272 201134 380620 201218
rect 380272 200898 380328 201134
rect 380564 200898 380620 201134
rect 380272 200866 380620 200898
rect 516000 201454 516348 201486
rect 516000 201218 516056 201454
rect 516292 201218 516348 201454
rect 516000 201134 516348 201218
rect 516000 200898 516056 201134
rect 516292 200898 516348 201134
rect 516000 200866 516348 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 380952 183454 381300 183486
rect 380952 183218 381008 183454
rect 381244 183218 381300 183454
rect 380952 183134 381300 183218
rect 380952 182898 381008 183134
rect 381244 182898 381300 183134
rect 380952 182866 381300 182898
rect 515320 183454 515668 183486
rect 515320 183218 515376 183454
rect 515612 183218 515668 183454
rect 515320 183134 515668 183218
rect 515320 182898 515376 183134
rect 515612 182898 515668 183134
rect 515320 182866 515668 182898
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 396056 164930 396116 165106
rect 397144 164930 397204 165106
rect 396030 164870 396116 164930
rect 397134 164870 397204 164930
rect 398232 164930 398292 165106
rect 399592 164930 399652 165106
rect 400544 164930 400604 165106
rect 401768 164930 401828 165106
rect 403128 164930 403188 165106
rect 404216 164930 404276 165106
rect 405440 164930 405500 165106
rect 406528 164930 406588 165106
rect 398232 164870 398298 164930
rect 379794 148394 380414 163000
rect 379794 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 380414 148394
rect 379794 148074 380414 148158
rect 379794 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 380414 148074
rect 379794 145308 380414 147838
rect 383514 152114 384134 163000
rect 383514 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 384134 152114
rect 383514 151794 384134 151878
rect 383514 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 384134 151794
rect 383514 145308 384134 151558
rect 387234 153954 387854 163000
rect 387234 153718 387266 153954
rect 387502 153718 387586 153954
rect 387822 153718 387854 153954
rect 387234 153634 387854 153718
rect 387234 153398 387266 153634
rect 387502 153398 387586 153634
rect 387822 153398 387854 153634
rect 387234 145308 387854 153398
rect 390954 157674 391574 163000
rect 396030 162757 396090 164870
rect 396027 162756 396093 162757
rect 396027 162692 396028 162756
rect 396092 162692 396093 162756
rect 396027 162691 396093 162692
rect 397134 162213 397194 164870
rect 398238 163165 398298 164870
rect 399526 164870 399652 164930
rect 400446 164870 400604 164930
rect 401734 164870 401828 164930
rect 403022 164870 403188 164930
rect 404126 164870 404276 164930
rect 405046 164870 405500 164930
rect 406518 164870 406588 164930
rect 407616 164930 407676 165106
rect 408296 164930 408356 165106
rect 408704 164930 408764 165106
rect 410064 164930 410124 165106
rect 407616 164870 407682 164930
rect 408296 164870 408418 164930
rect 408704 164870 408786 164930
rect 398235 163164 398301 163165
rect 398235 163100 398236 163164
rect 398300 163100 398301 163164
rect 398235 163099 398301 163100
rect 397131 162212 397197 162213
rect 397131 162148 397132 162212
rect 397196 162148 397197 162212
rect 397131 162147 397197 162148
rect 390954 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 391574 157674
rect 390954 157354 391574 157438
rect 390954 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 391574 157354
rect 390954 145308 391574 157118
rect 397794 147454 398414 163000
rect 399526 162757 399586 164870
rect 400446 162757 400506 164870
rect 401734 163165 401794 164870
rect 401731 163164 401797 163165
rect 401731 163100 401732 163164
rect 401796 163100 401797 163164
rect 401731 163099 401797 163100
rect 399523 162756 399589 162757
rect 399523 162692 399524 162756
rect 399588 162692 399589 162756
rect 399523 162691 399589 162692
rect 400443 162756 400509 162757
rect 400443 162692 400444 162756
rect 400508 162692 400509 162756
rect 400443 162691 400509 162692
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 145308 398414 146898
rect 401514 151174 402134 163000
rect 403022 162757 403082 164870
rect 403019 162756 403085 162757
rect 403019 162692 403020 162756
rect 403084 162692 403085 162756
rect 403019 162691 403085 162692
rect 404126 162213 404186 164870
rect 405046 162757 405106 164870
rect 405043 162756 405109 162757
rect 405043 162692 405044 162756
rect 405108 162692 405109 162756
rect 405043 162691 405109 162692
rect 404123 162212 404189 162213
rect 404123 162148 404124 162212
rect 404188 162148 404189 162212
rect 404123 162147 404189 162148
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 145308 402134 150618
rect 405234 154894 405854 163000
rect 406518 162757 406578 164870
rect 407622 162757 407682 164870
rect 408358 162757 408418 164870
rect 408726 162757 408786 164870
rect 410014 164870 410124 164930
rect 410744 164930 410804 165106
rect 411288 164930 411348 165106
rect 412376 164930 412436 165106
rect 410744 164870 410810 164930
rect 411288 164870 411362 164930
rect 412376 164870 412466 164930
rect 406515 162756 406581 162757
rect 406515 162692 406516 162756
rect 406580 162692 406581 162756
rect 406515 162691 406581 162692
rect 407619 162756 407685 162757
rect 407619 162692 407620 162756
rect 407684 162692 407685 162756
rect 407619 162691 407685 162692
rect 408355 162756 408421 162757
rect 408355 162692 408356 162756
rect 408420 162692 408421 162756
rect 408355 162691 408421 162692
rect 408723 162756 408789 162757
rect 408723 162692 408724 162756
rect 408788 162692 408789 162756
rect 408723 162691 408789 162692
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 145308 405854 154338
rect 408954 158614 409574 163000
rect 410014 162757 410074 164870
rect 410750 162757 410810 164870
rect 411302 162757 411362 164870
rect 410011 162756 410077 162757
rect 410011 162692 410012 162756
rect 410076 162692 410077 162756
rect 410011 162691 410077 162692
rect 410747 162756 410813 162757
rect 410747 162692 410748 162756
rect 410812 162692 410813 162756
rect 410747 162691 410813 162692
rect 411299 162756 411365 162757
rect 411299 162692 411300 162756
rect 411364 162692 411365 162756
rect 411299 162691 411365 162692
rect 412406 162213 412466 164870
rect 413464 164250 413524 165106
rect 413600 164930 413660 165106
rect 414552 164930 414612 165106
rect 415912 164930 415972 165106
rect 413600 164870 413754 164930
rect 414552 164870 414674 164930
rect 413464 164190 413570 164250
rect 413510 162757 413570 164190
rect 413694 162757 413754 164870
rect 414614 162757 414674 164870
rect 415534 164870 415972 164930
rect 416048 164930 416108 165106
rect 417000 164930 417060 165106
rect 418088 164930 418148 165106
rect 418496 164930 418556 165106
rect 419448 164930 419508 165106
rect 416048 164870 416146 164930
rect 417000 164870 417066 164930
rect 418088 164870 418170 164930
rect 415534 162757 415594 164870
rect 416086 164253 416146 164870
rect 416083 164252 416149 164253
rect 416083 164188 416084 164252
rect 416148 164188 416149 164252
rect 416083 164187 416149 164188
rect 413507 162756 413573 162757
rect 413507 162692 413508 162756
rect 413572 162692 413573 162756
rect 413507 162691 413573 162692
rect 413691 162756 413757 162757
rect 413691 162692 413692 162756
rect 413756 162692 413757 162756
rect 413691 162691 413757 162692
rect 414611 162756 414677 162757
rect 414611 162692 414612 162756
rect 414676 162692 414677 162756
rect 414611 162691 414677 162692
rect 415531 162756 415597 162757
rect 415531 162692 415532 162756
rect 415596 162692 415597 162756
rect 415531 162691 415597 162692
rect 412403 162212 412469 162213
rect 412403 162148 412404 162212
rect 412468 162148 412469 162212
rect 412403 162147 412469 162148
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 145308 409574 158058
rect 415794 148394 416414 163000
rect 417006 162757 417066 164870
rect 418110 162893 418170 164870
rect 418478 164870 418556 164930
rect 419214 164870 419508 164930
rect 420672 164930 420732 165106
rect 421080 164930 421140 165106
rect 420672 164870 420746 164930
rect 418107 162892 418173 162893
rect 418107 162828 418108 162892
rect 418172 162828 418173 162892
rect 418107 162827 418173 162828
rect 417003 162756 417069 162757
rect 417003 162692 417004 162756
rect 417068 162692 417069 162756
rect 417003 162691 417069 162692
rect 418478 162213 418538 164870
rect 419214 162757 419274 164870
rect 419211 162756 419277 162757
rect 419211 162692 419212 162756
rect 419276 162692 419277 162756
rect 419211 162691 419277 162692
rect 418475 162212 418541 162213
rect 418475 162148 418476 162212
rect 418540 162148 418541 162212
rect 418475 162147 418541 162148
rect 415794 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 416414 148394
rect 415794 148074 416414 148158
rect 415794 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 416414 148074
rect 415794 145308 416414 147838
rect 419514 152114 420134 163000
rect 420686 162757 420746 164870
rect 421054 164870 421140 164930
rect 421760 164930 421820 165106
rect 422848 164930 422908 165106
rect 421760 164870 421850 164930
rect 422848 164870 422954 164930
rect 421054 164253 421114 164870
rect 421051 164252 421117 164253
rect 421051 164188 421052 164252
rect 421116 164188 421117 164252
rect 421051 164187 421117 164188
rect 421790 162757 421850 164870
rect 422894 162757 422954 164870
rect 423528 164661 423588 165106
rect 423936 164930 423996 165106
rect 425296 164930 425356 165106
rect 423936 164870 424058 164930
rect 423525 164660 423591 164661
rect 423525 164596 423526 164660
rect 423590 164596 423591 164660
rect 423525 164595 423591 164596
rect 420683 162756 420749 162757
rect 420683 162692 420684 162756
rect 420748 162692 420749 162756
rect 420683 162691 420749 162692
rect 421787 162756 421853 162757
rect 421787 162692 421788 162756
rect 421852 162692 421853 162756
rect 421787 162691 421853 162692
rect 422891 162756 422957 162757
rect 422891 162692 422892 162756
rect 422956 162692 422957 162756
rect 422891 162691 422957 162692
rect 419514 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 420134 152114
rect 419514 151794 420134 151878
rect 419514 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 420134 151794
rect 419514 145308 420134 151558
rect 423234 153954 423854 163000
rect 423998 162757 424058 164870
rect 425286 164870 425356 164930
rect 425286 162757 425346 164870
rect 425976 164797 426036 165106
rect 426384 164930 426444 165106
rect 427608 164930 427668 165106
rect 428288 164930 428348 165106
rect 426384 164870 426450 164930
rect 427608 164870 427738 164930
rect 425973 164796 426039 164797
rect 425973 164732 425974 164796
rect 426038 164732 426039 164796
rect 425973 164731 426039 164732
rect 426390 162757 426450 164870
rect 423995 162756 424061 162757
rect 423995 162692 423996 162756
rect 424060 162692 424061 162756
rect 423995 162691 424061 162692
rect 425283 162756 425349 162757
rect 425283 162692 425284 162756
rect 425348 162692 425349 162756
rect 425283 162691 425349 162692
rect 426387 162756 426453 162757
rect 426387 162692 426388 162756
rect 426452 162692 426453 162756
rect 426387 162691 426453 162692
rect 423234 153718 423266 153954
rect 423502 153718 423586 153954
rect 423822 153718 423854 153954
rect 423234 153634 423854 153718
rect 423234 153398 423266 153634
rect 423502 153398 423586 153634
rect 423822 153398 423854 153634
rect 423234 145308 423854 153398
rect 426954 157674 427574 163000
rect 427678 162213 427738 164870
rect 428230 164870 428348 164930
rect 428696 164930 428756 165106
rect 429784 164930 429844 165106
rect 431008 164930 431068 165106
rect 428696 164870 428842 164930
rect 428230 164253 428290 164870
rect 428227 164252 428293 164253
rect 428227 164188 428228 164252
rect 428292 164188 428293 164252
rect 428227 164187 428293 164188
rect 428782 162757 428842 164870
rect 429702 164870 429844 164930
rect 430990 164870 431068 164930
rect 431144 164930 431204 165106
rect 432232 164930 432292 165106
rect 431144 164870 431234 164930
rect 429702 162757 429762 164870
rect 430990 164253 431050 164870
rect 430987 164252 431053 164253
rect 430987 164188 430988 164252
rect 431052 164188 431053 164252
rect 430987 164187 431053 164188
rect 431174 162757 431234 164870
rect 432094 164870 432292 164930
rect 433320 164930 433380 165106
rect 433592 164930 433652 165106
rect 433320 164870 433442 164930
rect 432094 164250 432154 164870
rect 431726 164190 432154 164250
rect 431726 162757 431786 164190
rect 433382 162757 433442 164870
rect 433566 164870 433652 164930
rect 428779 162756 428845 162757
rect 428779 162692 428780 162756
rect 428844 162692 428845 162756
rect 428779 162691 428845 162692
rect 429699 162756 429765 162757
rect 429699 162692 429700 162756
rect 429764 162692 429765 162756
rect 429699 162691 429765 162692
rect 431171 162756 431237 162757
rect 431171 162692 431172 162756
rect 431236 162692 431237 162756
rect 431171 162691 431237 162692
rect 431723 162756 431789 162757
rect 431723 162692 431724 162756
rect 431788 162692 431789 162756
rect 431723 162691 431789 162692
rect 433379 162756 433445 162757
rect 433379 162692 433380 162756
rect 433444 162692 433445 162756
rect 433379 162691 433445 162692
rect 433566 162213 433626 164870
rect 434408 164797 434468 165106
rect 435768 164930 435828 165106
rect 436040 164930 436100 165106
rect 435768 164870 435834 164930
rect 434405 164796 434471 164797
rect 434405 164732 434406 164796
rect 434470 164732 434471 164796
rect 434405 164731 434471 164732
rect 427675 162212 427741 162213
rect 427675 162148 427676 162212
rect 427740 162148 427741 162212
rect 427675 162147 427741 162148
rect 433563 162212 433629 162213
rect 433563 162148 433564 162212
rect 433628 162148 433629 162212
rect 433563 162147 433629 162148
rect 426954 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 427574 157674
rect 426954 157354 427574 157438
rect 426954 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 427574 157354
rect 426954 145308 427574 157118
rect 433794 147454 434414 163000
rect 435774 162757 435834 164870
rect 435958 164870 436100 164930
rect 435958 162757 436018 164870
rect 436992 164661 437052 165106
rect 438080 164661 438140 165106
rect 438488 164930 438548 165106
rect 439168 164930 439228 165106
rect 440936 164930 440996 165106
rect 443520 164930 443580 165106
rect 445968 164930 446028 165106
rect 438488 164870 438594 164930
rect 436989 164660 437055 164661
rect 436989 164596 436990 164660
rect 437054 164596 437055 164660
rect 436989 164595 437055 164596
rect 438077 164660 438143 164661
rect 438077 164596 438078 164660
rect 438142 164596 438143 164660
rect 438077 164595 438143 164596
rect 435771 162756 435837 162757
rect 435771 162692 435772 162756
rect 435836 162692 435837 162756
rect 435771 162691 435837 162692
rect 435955 162756 436021 162757
rect 435955 162692 435956 162756
rect 436020 162692 436021 162756
rect 435955 162691 436021 162692
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 145308 434414 146898
rect 437514 151174 438134 163000
rect 438534 162757 438594 164870
rect 439086 164870 439228 164930
rect 440926 164870 440996 164930
rect 443502 164870 443580 164930
rect 445894 164870 446028 164930
rect 448280 164930 448340 165106
rect 448280 164870 448346 164930
rect 439086 162757 439146 164870
rect 440926 162757 440986 164870
rect 438531 162756 438597 162757
rect 438531 162692 438532 162756
rect 438596 162692 438597 162756
rect 438531 162691 438597 162692
rect 439083 162756 439149 162757
rect 439083 162692 439084 162756
rect 439148 162692 439149 162756
rect 439083 162691 439149 162692
rect 440923 162756 440989 162757
rect 440923 162692 440924 162756
rect 440988 162692 440989 162756
rect 440923 162691 440989 162692
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 145308 438134 150618
rect 441234 154894 441854 163000
rect 443502 162757 443562 164870
rect 443499 162756 443565 162757
rect 443499 162692 443500 162756
rect 443564 162692 443565 162756
rect 443499 162691 443565 162692
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 145308 441854 154338
rect 444954 158614 445574 163000
rect 445894 162757 445954 164870
rect 448286 162757 448346 164870
rect 451000 164797 451060 165106
rect 450997 164796 451063 164797
rect 450997 164732 450998 164796
rect 451062 164732 451063 164796
rect 453448 164794 453508 165106
rect 455896 164930 455956 165106
rect 458480 164930 458540 165106
rect 450997 164731 451063 164732
rect 453438 164734 453508 164794
rect 455830 164870 455956 164930
rect 458406 164870 458540 164930
rect 460928 164930 460988 165106
rect 463512 164930 463572 165106
rect 465960 164930 466020 165106
rect 468544 164930 468604 165106
rect 470992 164930 471052 165106
rect 460928 164870 461042 164930
rect 445891 162756 445957 162757
rect 445891 162692 445892 162756
rect 445956 162692 445957 162756
rect 445891 162691 445957 162692
rect 448283 162756 448349 162757
rect 448283 162692 448284 162756
rect 448348 162692 448349 162756
rect 448283 162691 448349 162692
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 145308 445574 158058
rect 451794 148394 452414 163000
rect 453438 162757 453498 164734
rect 455830 163165 455890 164870
rect 455827 163164 455893 163165
rect 455827 163100 455828 163164
rect 455892 163100 455893 163164
rect 455827 163099 455893 163100
rect 453435 162756 453501 162757
rect 453435 162692 453436 162756
rect 453500 162692 453501 162756
rect 453435 162691 453501 162692
rect 451794 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 452414 148394
rect 451794 148074 452414 148158
rect 451794 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 452414 148074
rect 451794 145308 452414 147838
rect 455514 152114 456134 163000
rect 458406 162757 458466 164870
rect 458403 162756 458469 162757
rect 458403 162692 458404 162756
rect 458468 162692 458469 162756
rect 458403 162691 458469 162692
rect 455514 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 456134 152114
rect 455514 151794 456134 151878
rect 455514 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 456134 151794
rect 455514 145308 456134 151558
rect 459234 153954 459854 163000
rect 460982 162349 461042 164870
rect 462638 164870 463572 164930
rect 465950 164870 466020 164930
rect 468526 164870 468604 164930
rect 470918 164870 471052 164930
rect 473440 164930 473500 165106
rect 475888 164930 475948 165106
rect 478472 164930 478532 165106
rect 473440 164870 473554 164930
rect 462638 162485 462698 164870
rect 462635 162484 462701 162485
rect 462635 162420 462636 162484
rect 462700 162420 462701 162484
rect 462635 162419 462701 162420
rect 460979 162348 461045 162349
rect 460979 162284 460980 162348
rect 461044 162284 461045 162348
rect 460979 162283 461045 162284
rect 459234 153718 459266 153954
rect 459502 153718 459586 153954
rect 459822 153718 459854 153954
rect 459234 153634 459854 153718
rect 459234 153398 459266 153634
rect 459502 153398 459586 153634
rect 459822 153398 459854 153634
rect 459234 145308 459854 153398
rect 462954 157674 463574 163000
rect 465950 162621 466010 164870
rect 465947 162620 466013 162621
rect 465947 162556 465948 162620
rect 466012 162556 466013 162620
rect 465947 162555 466013 162556
rect 468526 161941 468586 164870
rect 470918 164250 470978 164870
rect 473494 164253 473554 164870
rect 475886 164870 475948 164930
rect 478462 164870 478532 164930
rect 475886 164253 475946 164870
rect 478462 164253 478522 164870
rect 480920 164661 480980 165106
rect 483368 164930 483428 165106
rect 485952 164930 486012 165106
rect 503224 164930 503284 165106
rect 483368 164870 483490 164930
rect 485952 164870 486066 164930
rect 480917 164660 480983 164661
rect 480917 164596 480918 164660
rect 480982 164596 480983 164660
rect 480917 164595 480983 164596
rect 470366 164190 470978 164250
rect 473491 164252 473557 164253
rect 470366 163845 470426 164190
rect 473491 164188 473492 164252
rect 473556 164188 473557 164252
rect 473491 164187 473557 164188
rect 475883 164252 475949 164253
rect 475883 164188 475884 164252
rect 475948 164188 475949 164252
rect 475883 164187 475949 164188
rect 478459 164252 478525 164253
rect 478459 164188 478460 164252
rect 478524 164188 478525 164252
rect 478459 164187 478525 164188
rect 483430 163981 483490 164870
rect 486006 164117 486066 164870
rect 503118 164870 503284 164930
rect 503360 164930 503420 165106
rect 503360 164870 503546 164930
rect 486003 164116 486069 164117
rect 486003 164052 486004 164116
rect 486068 164052 486069 164116
rect 486003 164051 486069 164052
rect 483427 163980 483493 163981
rect 483427 163916 483428 163980
rect 483492 163916 483493 163980
rect 483427 163915 483493 163916
rect 470363 163844 470429 163845
rect 470363 163780 470364 163844
rect 470428 163780 470429 163844
rect 470363 163779 470429 163780
rect 468523 161940 468589 161941
rect 468523 161876 468524 161940
rect 468588 161876 468589 161940
rect 468523 161875 468589 161876
rect 462954 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 463574 157674
rect 462954 157354 463574 157438
rect 462954 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 463574 157354
rect 462954 145308 463574 157118
rect 469794 147454 470414 163000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 145308 470414 146898
rect 473514 151174 474134 163000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 145308 474134 150618
rect 477234 154894 477854 163000
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 145308 477854 154338
rect 480954 158614 481574 163000
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 145308 481574 158058
rect 487794 148394 488414 163000
rect 487794 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 487794 148074 488414 148158
rect 487794 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 487794 145308 488414 147838
rect 491514 152114 492134 163000
rect 491514 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 491514 151794 492134 151878
rect 491514 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 491514 145308 492134 151558
rect 495234 153954 495854 163000
rect 495234 153718 495266 153954
rect 495502 153718 495586 153954
rect 495822 153718 495854 153954
rect 495234 153634 495854 153718
rect 495234 153398 495266 153634
rect 495502 153398 495586 153634
rect 495822 153398 495854 153634
rect 495234 145308 495854 153398
rect 498954 157674 499574 163000
rect 503118 162757 503178 164870
rect 503115 162756 503181 162757
rect 503115 162692 503116 162756
rect 503180 162692 503181 162756
rect 503115 162691 503181 162692
rect 503486 162621 503546 164870
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 503483 162620 503549 162621
rect 503483 162556 503484 162620
rect 503548 162556 503549 162620
rect 503483 162555 503549 162556
rect 498954 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 498954 157354 499574 157438
rect 498954 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 498954 145308 499574 157118
rect 505794 147454 506414 163000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 145308 506414 146898
rect 509514 151174 510134 163000
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 145308 510134 150618
rect 513234 154894 513854 163000
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 510843 146164 510909 146165
rect 510843 146100 510844 146164
rect 510908 146100 510909 146164
rect 510843 146099 510909 146100
rect 498515 144940 498581 144941
rect 498515 144876 498516 144940
rect 498580 144876 498581 144940
rect 498515 144875 498581 144876
rect 499803 144940 499869 144941
rect 499803 144876 499804 144940
rect 499868 144876 499869 144940
rect 499803 144875 499869 144876
rect 498518 143850 498578 144875
rect 499806 143850 499866 144875
rect 510846 143850 510906 146099
rect 513234 145308 513854 154338
rect 516954 158614 517574 163000
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 145308 517574 158058
rect 498464 143790 498578 143850
rect 499688 143790 499866 143850
rect 510840 143790 510906 143850
rect 498464 143202 498524 143790
rect 499688 143202 499748 143790
rect 510840 143202 510900 143790
rect 380272 129454 380620 129486
rect 380272 129218 380328 129454
rect 380564 129218 380620 129454
rect 380272 129134 380620 129218
rect 380272 128898 380328 129134
rect 380564 128898 380620 129134
rect 380272 128866 380620 128898
rect 516000 129454 516348 129486
rect 516000 129218 516056 129454
rect 516292 129218 516348 129454
rect 516000 129134 516348 129218
rect 516000 128898 516056 129134
rect 516292 128898 516348 129134
rect 516000 128866 516348 128898
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 380952 111454 381300 111486
rect 380952 111218 381008 111454
rect 381244 111218 381300 111454
rect 380952 111134 381300 111218
rect 380952 110898 381008 111134
rect 381244 110898 381300 111134
rect 380952 110866 381300 110898
rect 515320 111454 515668 111486
rect 515320 111218 515376 111454
rect 515612 111218 515668 111454
rect 515320 111134 515668 111218
rect 515320 110898 515376 111134
rect 515612 110898 515668 111134
rect 515320 110866 515668 110898
rect 380272 93454 380620 93486
rect 380272 93218 380328 93454
rect 380564 93218 380620 93454
rect 380272 93134 380620 93218
rect 380272 92898 380328 93134
rect 380564 92898 380620 93134
rect 380272 92866 380620 92898
rect 516000 93454 516348 93486
rect 516000 93218 516056 93454
rect 516292 93218 516348 93454
rect 516000 93134 516348 93218
rect 516000 92898 516056 93134
rect 516292 92898 516348 93134
rect 516000 92866 516348 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 380952 75454 381300 75486
rect 380952 75218 381008 75454
rect 381244 75218 381300 75454
rect 380952 75134 381300 75218
rect 380952 74898 381008 75134
rect 381244 74898 381300 75134
rect 380952 74866 381300 74898
rect 515320 75454 515668 75486
rect 515320 75218 515376 75454
rect 515612 75218 515668 75454
rect 515320 75134 515668 75218
rect 515320 74898 515376 75134
rect 515612 74898 515668 75134
rect 515320 74866 515668 74898
rect 396056 59805 396116 60106
rect 397144 59805 397204 60106
rect 396053 59804 396119 59805
rect 396053 59740 396054 59804
rect 396118 59740 396119 59804
rect 396053 59739 396119 59740
rect 397141 59804 397207 59805
rect 397141 59740 397142 59804
rect 397206 59740 397207 59804
rect 397141 59739 397207 59740
rect 398232 59530 398292 60106
rect 399592 59666 399652 60106
rect 400544 59666 400604 60106
rect 399526 59606 399652 59666
rect 400446 59606 400604 59666
rect 398232 59470 398298 59530
rect 398238 58173 398298 59470
rect 398235 58172 398301 58173
rect 398235 58108 398236 58172
rect 398300 58108 398301 58172
rect 398235 58107 398301 58108
rect 379794 57454 380414 58000
rect 379099 57220 379165 57221
rect 379099 57156 379100 57220
rect 379164 57156 379165 57220
rect 379099 57155 379165 57156
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 378731 57084 378797 57085
rect 378731 57020 378732 57084
rect 378796 57020 378797 57084
rect 378731 57019 378797 57020
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 377443 55180 377509 55181
rect 377443 55116 377444 55180
rect 377508 55116 377509 55180
rect 377443 55115 377509 55116
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 399526 57901 399586 59606
rect 400446 57901 400506 59606
rect 401768 59530 401828 60106
rect 403128 59669 403188 60106
rect 404216 59669 404276 60106
rect 403125 59668 403191 59669
rect 403125 59604 403126 59668
rect 403190 59604 403191 59668
rect 403125 59603 403191 59604
rect 404213 59668 404279 59669
rect 404213 59604 404214 59668
rect 404278 59604 404279 59668
rect 404213 59603 404279 59604
rect 405440 59530 405500 60106
rect 406528 59530 406588 60106
rect 401734 59470 401828 59530
rect 405414 59470 405500 59530
rect 406518 59470 406588 59530
rect 407616 59530 407676 60106
rect 408296 59530 408356 60106
rect 408704 59530 408764 60106
rect 410064 59530 410124 60106
rect 407616 59470 407682 59530
rect 408296 59470 408418 59530
rect 408704 59470 408786 59530
rect 401734 58173 401794 59470
rect 405414 58173 405474 59470
rect 401731 58172 401797 58173
rect 401731 58108 401732 58172
rect 401796 58108 401797 58172
rect 401731 58107 401797 58108
rect 405411 58172 405477 58173
rect 405411 58108 405412 58172
rect 405476 58108 405477 58172
rect 405411 58107 405477 58108
rect 399523 57900 399589 57901
rect 399523 57836 399524 57900
rect 399588 57836 399589 57900
rect 399523 57835 399589 57836
rect 400443 57900 400509 57901
rect 400443 57836 400444 57900
rect 400508 57836 400509 57900
rect 400443 57835 400509 57836
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 406518 57901 406578 59470
rect 407622 57901 407682 59470
rect 408358 57901 408418 59470
rect 408726 57901 408786 59470
rect 410014 59470 410124 59530
rect 410744 59530 410804 60106
rect 411288 59530 411348 60106
rect 412376 59530 412436 60106
rect 413464 59669 413524 60106
rect 413461 59668 413527 59669
rect 413461 59604 413462 59668
rect 413526 59604 413527 59668
rect 413461 59603 413527 59604
rect 413600 59530 413660 60106
rect 410744 59470 410810 59530
rect 411288 59470 411362 59530
rect 412376 59470 412466 59530
rect 406515 57900 406581 57901
rect 406515 57836 406516 57900
rect 406580 57836 406581 57900
rect 406515 57835 406581 57836
rect 407619 57900 407685 57901
rect 407619 57836 407620 57900
rect 407684 57836 407685 57900
rect 407619 57835 407685 57836
rect 408355 57900 408421 57901
rect 408355 57836 408356 57900
rect 408420 57836 408421 57900
rect 408355 57835 408421 57836
rect 408723 57900 408789 57901
rect 408723 57836 408724 57900
rect 408788 57836 408789 57900
rect 408723 57835 408789 57836
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 410014 57901 410074 59470
rect 410011 57900 410077 57901
rect 410011 57836 410012 57900
rect 410076 57836 410077 57900
rect 410011 57835 410077 57836
rect 410750 56541 410810 59470
rect 411302 56949 411362 59470
rect 412406 57901 412466 59470
rect 413510 59470 413660 59530
rect 414552 59530 414612 60106
rect 415912 59530 415972 60106
rect 414552 59470 414674 59530
rect 412403 57900 412469 57901
rect 412403 57836 412404 57900
rect 412468 57836 412469 57900
rect 412403 57835 412469 57836
rect 413510 57085 413570 59470
rect 414614 57901 414674 59470
rect 415534 59470 415972 59530
rect 416048 59530 416108 60106
rect 417000 59805 417060 60106
rect 416997 59804 417063 59805
rect 416997 59740 416998 59804
rect 417062 59740 417063 59804
rect 416997 59739 417063 59740
rect 418088 59533 418148 60106
rect 418496 59805 418556 60106
rect 418493 59804 418559 59805
rect 418493 59740 418494 59804
rect 418558 59740 418559 59804
rect 418493 59739 418559 59740
rect 418088 59532 418173 59533
rect 416048 59470 416146 59530
rect 418088 59470 418108 59532
rect 415534 57901 415594 59470
rect 416086 58173 416146 59470
rect 418107 59468 418108 59470
rect 418172 59468 418173 59532
rect 419448 59530 419508 60106
rect 418107 59467 418173 59468
rect 419398 59470 419508 59530
rect 420672 59530 420732 60106
rect 421080 59530 421140 60106
rect 420672 59470 420746 59530
rect 419398 58445 419458 59470
rect 420686 59397 420746 59470
rect 421054 59470 421140 59530
rect 421760 59530 421820 60106
rect 422848 59805 422908 60106
rect 422845 59804 422911 59805
rect 422845 59740 422846 59804
rect 422910 59740 422911 59804
rect 422845 59739 422911 59740
rect 423528 59669 423588 60106
rect 423936 59805 423996 60106
rect 423933 59804 423999 59805
rect 423933 59740 423934 59804
rect 423998 59740 423999 59804
rect 423933 59739 423999 59740
rect 423525 59668 423591 59669
rect 423525 59604 423526 59668
rect 423590 59604 423591 59668
rect 423525 59603 423591 59604
rect 425296 59530 425356 60106
rect 421760 59470 421850 59530
rect 420683 59396 420749 59397
rect 420683 59332 420684 59396
rect 420748 59332 420749 59396
rect 420683 59331 420749 59332
rect 419395 58444 419461 58445
rect 419395 58380 419396 58444
rect 419460 58380 419461 58444
rect 419395 58379 419461 58380
rect 416083 58172 416149 58173
rect 416083 58108 416084 58172
rect 416148 58108 416149 58172
rect 416083 58107 416149 58108
rect 414611 57900 414677 57901
rect 414611 57836 414612 57900
rect 414676 57836 414677 57900
rect 414611 57835 414677 57836
rect 415531 57900 415597 57901
rect 415531 57836 415532 57900
rect 415596 57836 415597 57900
rect 415531 57835 415597 57836
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 413507 57084 413573 57085
rect 413507 57020 413508 57084
rect 413572 57020 413573 57084
rect 413507 57019 413573 57020
rect 411299 56948 411365 56949
rect 411299 56884 411300 56948
rect 411364 56884 411365 56948
rect 411299 56883 411365 56884
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 410747 56540 410813 56541
rect 410747 56476 410748 56540
rect 410812 56476 410813 56540
rect 410747 56475 410813 56476
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 421054 57221 421114 59470
rect 421790 59397 421850 59470
rect 425286 59470 425356 59530
rect 425976 59530 426036 60106
rect 426384 59530 426444 60106
rect 427608 59530 427668 60106
rect 428288 59530 428348 60106
rect 428696 59530 428756 60106
rect 429784 59530 429844 60106
rect 431008 59530 431068 60106
rect 425976 59470 426082 59530
rect 426384 59470 426450 59530
rect 427608 59470 427738 59530
rect 421787 59396 421853 59397
rect 421787 59332 421788 59396
rect 421852 59332 421853 59396
rect 421787 59331 421853 59332
rect 425286 58581 425346 59470
rect 426022 59397 426082 59470
rect 426019 59396 426085 59397
rect 426019 59332 426020 59396
rect 426084 59332 426085 59396
rect 426019 59331 426085 59332
rect 425283 58580 425349 58581
rect 425283 58516 425284 58580
rect 425348 58516 425349 58580
rect 425283 58515 425349 58516
rect 421051 57220 421117 57221
rect 421051 57156 421052 57220
rect 421116 57156 421117 57220
rect 421051 57155 421117 57156
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 426390 57901 426450 59470
rect 426387 57900 426453 57901
rect 426387 57836 426388 57900
rect 426452 57836 426453 57900
rect 426387 57835 426453 57836
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 427678 57901 427738 59470
rect 428230 59470 428348 59530
rect 428598 59470 428756 59530
rect 429702 59470 429844 59530
rect 430990 59470 431068 59530
rect 431144 59530 431204 60106
rect 432232 59530 432292 60106
rect 433320 59530 433380 60106
rect 433592 59530 433652 60106
rect 431144 59470 431234 59530
rect 432232 59470 432338 59530
rect 433320 59470 433442 59530
rect 428230 59397 428290 59470
rect 428227 59396 428293 59397
rect 428227 59332 428228 59396
rect 428292 59332 428293 59396
rect 428227 59331 428293 59332
rect 428598 57901 428658 59470
rect 429702 57901 429762 59470
rect 427675 57900 427741 57901
rect 427675 57836 427676 57900
rect 427740 57836 427741 57900
rect 427675 57835 427741 57836
rect 428595 57900 428661 57901
rect 428595 57836 428596 57900
rect 428660 57836 428661 57900
rect 428595 57835 428661 57836
rect 429699 57900 429765 57901
rect 429699 57836 429700 57900
rect 429764 57836 429765 57900
rect 429699 57835 429765 57836
rect 430990 57221 431050 59470
rect 431174 57901 431234 59470
rect 432278 57901 432338 59470
rect 433382 57901 433442 59470
rect 433566 59470 433652 59530
rect 434408 59530 434468 60106
rect 435768 59530 435828 60106
rect 436040 59530 436100 60106
rect 436992 59530 437052 60106
rect 434408 59470 434730 59530
rect 435768 59470 435834 59530
rect 433566 57901 433626 59470
rect 431171 57900 431237 57901
rect 431171 57836 431172 57900
rect 431236 57836 431237 57900
rect 431171 57835 431237 57836
rect 432275 57900 432341 57901
rect 432275 57836 432276 57900
rect 432340 57836 432341 57900
rect 432275 57835 432341 57836
rect 433379 57900 433445 57901
rect 433379 57836 433380 57900
rect 433444 57836 433445 57900
rect 433379 57835 433445 57836
rect 433563 57900 433629 57901
rect 433563 57836 433564 57900
rect 433628 57836 433629 57900
rect 433563 57835 433629 57836
rect 430987 57220 431053 57221
rect 430987 57156 430988 57220
rect 431052 57156 431053 57220
rect 430987 57155 431053 57156
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 434670 57221 434730 59470
rect 435774 57221 435834 59470
rect 435958 59470 436100 59530
rect 436878 59470 437052 59530
rect 438080 59530 438140 60106
rect 438488 59530 438548 60106
rect 439168 59530 439228 60106
rect 440936 59530 440996 60106
rect 443520 59530 443580 60106
rect 445968 59530 446028 60106
rect 438080 59470 438410 59530
rect 438488 59470 438594 59530
rect 435958 57901 436018 59470
rect 436878 57901 436938 59470
rect 435955 57900 436021 57901
rect 435955 57836 435956 57900
rect 436020 57836 436021 57900
rect 435955 57835 436021 57836
rect 436875 57900 436941 57901
rect 436875 57836 436876 57900
rect 436940 57836 436941 57900
rect 436875 57835 436941 57836
rect 434667 57220 434733 57221
rect 434667 57156 434668 57220
rect 434732 57156 434733 57220
rect 434667 57155 434733 57156
rect 435771 57220 435837 57221
rect 435771 57156 435772 57220
rect 435836 57156 435837 57220
rect 435771 57155 435837 57156
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 438350 57901 438410 59470
rect 438534 57901 438594 59470
rect 439086 59470 439228 59530
rect 440926 59470 440996 59530
rect 443502 59470 443580 59530
rect 445894 59470 446028 59530
rect 448280 59530 448340 60106
rect 451000 59530 451060 60106
rect 453448 59530 453508 60106
rect 448280 59470 448346 59530
rect 451000 59470 451106 59530
rect 439086 57901 439146 59470
rect 440926 57901 440986 59470
rect 438347 57900 438413 57901
rect 438347 57836 438348 57900
rect 438412 57836 438413 57900
rect 438347 57835 438413 57836
rect 438531 57900 438597 57901
rect 438531 57836 438532 57900
rect 438596 57836 438597 57900
rect 438531 57835 438597 57836
rect 439083 57900 439149 57901
rect 439083 57836 439084 57900
rect 439148 57836 439149 57900
rect 439083 57835 439149 57836
rect 440923 57900 440989 57901
rect 440923 57836 440924 57900
rect 440988 57836 440989 57900
rect 440923 57835 440989 57836
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 443502 57901 443562 59470
rect 443499 57900 443565 57901
rect 443499 57836 443500 57900
rect 443564 57836 443565 57900
rect 443499 57835 443565 57836
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 445894 57493 445954 59470
rect 448286 57901 448346 59470
rect 448283 57900 448349 57901
rect 448283 57836 448284 57900
rect 448348 57836 448349 57900
rect 448283 57835 448349 57836
rect 451046 57765 451106 59470
rect 453438 59470 453508 59530
rect 455896 59530 455956 60106
rect 458480 59530 458540 60106
rect 455896 59470 456442 59530
rect 453438 59397 453498 59470
rect 453435 59396 453501 59397
rect 453435 59332 453436 59396
rect 453500 59332 453501 59396
rect 453435 59331 453501 59332
rect 451043 57764 451109 57765
rect 451043 57700 451044 57764
rect 451108 57700 451109 57764
rect 451043 57699 451109 57700
rect 445891 57492 445957 57493
rect 445891 57428 445892 57492
rect 445956 57428 445957 57492
rect 445891 57427 445957 57428
rect 451794 57454 452414 58000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 456382 57357 456442 59470
rect 458406 59470 458540 59530
rect 460928 59530 460988 60106
rect 463512 59530 463572 60106
rect 465960 59530 466020 60106
rect 468544 59530 468604 60106
rect 470992 59530 471052 60106
rect 460928 59470 461042 59530
rect 463512 59470 463618 59530
rect 458406 58717 458466 59470
rect 458403 58716 458469 58717
rect 458403 58652 458404 58716
rect 458468 58652 458469 58716
rect 458403 58651 458469 58652
rect 456379 57356 456445 57357
rect 456379 57292 456380 57356
rect 456444 57292 456445 57356
rect 456379 57291 456445 57292
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 460982 57629 461042 59470
rect 463558 59397 463618 59470
rect 465950 59470 466020 59530
rect 468526 59470 468604 59530
rect 470918 59470 471052 59530
rect 473440 59530 473500 60106
rect 475888 59530 475948 60106
rect 478472 59530 478532 60106
rect 480920 59669 480980 60106
rect 480917 59668 480983 59669
rect 480917 59604 480918 59668
rect 480982 59604 480983 59668
rect 480917 59603 480983 59604
rect 473440 59470 473554 59530
rect 463555 59396 463621 59397
rect 463555 59332 463556 59396
rect 463620 59332 463621 59396
rect 463555 59331 463621 59332
rect 460979 57628 461045 57629
rect 460979 57564 460980 57628
rect 461044 57564 461045 57628
rect 460979 57563 461045 57564
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 465950 56677 466010 59470
rect 468526 59125 468586 59470
rect 468523 59124 468589 59125
rect 468523 59060 468524 59124
rect 468588 59060 468589 59124
rect 468523 59059 468589 59060
rect 465947 56676 466013 56677
rect 465947 56612 465948 56676
rect 466012 56612 466013 56676
rect 465947 56611 466013 56612
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 470918 57901 470978 59470
rect 473494 58989 473554 59470
rect 475886 59470 475948 59530
rect 478462 59470 478532 59530
rect 483368 59530 483428 60106
rect 485952 59530 486012 60106
rect 503224 59530 503284 60106
rect 483368 59470 483490 59530
rect 485952 59470 486066 59530
rect 473491 58988 473557 58989
rect 473491 58924 473492 58988
rect 473556 58924 473557 58988
rect 473491 58923 473557 58924
rect 475886 58853 475946 59470
rect 475883 58852 475949 58853
rect 475883 58788 475884 58852
rect 475948 58788 475949 58852
rect 475883 58787 475949 58788
rect 470915 57900 470981 57901
rect 470915 57836 470916 57900
rect 470980 57836 470981 57900
rect 470915 57835 470981 57836
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 478462 57901 478522 59470
rect 483430 59261 483490 59470
rect 486006 59261 486066 59470
rect 503118 59470 503284 59530
rect 503360 59530 503420 60106
rect 503360 59470 503546 59530
rect 483427 59260 483493 59261
rect 483427 59196 483428 59260
rect 483492 59196 483493 59260
rect 483427 59195 483493 59196
rect 486003 59260 486069 59261
rect 486003 59196 486004 59260
rect 486068 59196 486069 59260
rect 486003 59195 486069 59196
rect 478459 57900 478525 57901
rect 478459 57836 478460 57900
rect 478524 57836 478525 57900
rect 478459 57835 478525 57836
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 503118 57901 503178 59470
rect 503486 57901 503546 59470
rect 503115 57900 503181 57901
rect 503115 57836 503116 57900
rect 503180 57836 503181 57900
rect 503115 57835 503181 57836
rect 503483 57900 503549 57901
rect 503483 57836 503484 57900
rect 503548 57836 503549 57900
rect 503483 57835 503549 57836
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 79610 597218 79846 597454
rect 79610 596898 79846 597134
rect 110330 597218 110566 597454
rect 110330 596898 110566 597134
rect 64250 579218 64486 579454
rect 64250 578898 64486 579134
rect 94970 579218 95206 579454
rect 94970 578898 95206 579134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 59546 547878 59782 548114
rect 59866 547878 60102 548114
rect 59546 547558 59782 547794
rect 59866 547558 60102 547794
rect 63266 549718 63502 549954
rect 63586 549718 63822 549954
rect 63266 549398 63502 549634
rect 63586 549398 63822 549634
rect 66986 553438 67222 553674
rect 67306 553438 67542 553674
rect 66986 553118 67222 553354
rect 67306 553118 67542 553354
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 91826 544158 92062 544394
rect 92146 544158 92382 544394
rect 91826 543838 92062 544074
rect 92146 543838 92382 544074
rect 95546 547878 95782 548114
rect 95866 547878 96102 548114
rect 95546 547558 95782 547794
rect 95866 547558 96102 547794
rect 99266 549718 99502 549954
rect 99586 549718 99822 549954
rect 99266 549398 99502 549634
rect 99586 549398 99822 549634
rect 102986 553438 103222 553674
rect 103306 553438 103542 553674
rect 102986 553118 103222 553354
rect 103306 553118 103542 553354
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 127826 544158 128062 544394
rect 128146 544158 128382 544394
rect 127826 543838 128062 544074
rect 128146 543838 128382 544074
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 547878 131782 548114
rect 131866 547878 132102 548114
rect 131546 547558 131782 547794
rect 131866 547558 132102 547794
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 144250 615218 144486 615454
rect 144250 614898 144486 615134
rect 174970 615218 175206 615454
rect 174970 614898 175206 615134
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 159610 597218 159846 597454
rect 159610 596898 159846 597134
rect 190330 597218 190566 597454
rect 190330 596898 190566 597134
rect 144250 579218 144486 579454
rect 144250 578898 144486 579134
rect 174970 579218 175206 579454
rect 174970 578898 175206 579134
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 135266 549718 135502 549954
rect 135586 549718 135822 549954
rect 135266 549398 135502 549634
rect 135586 549398 135822 549634
rect 138986 553438 139222 553674
rect 139306 553438 139542 553674
rect 138986 553118 139222 553354
rect 139306 553118 139542 553354
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 544158 164062 544394
rect 164146 544158 164382 544394
rect 163826 543838 164062 544074
rect 164146 543838 164382 544074
rect 167546 547878 167782 548114
rect 167866 547878 168102 548114
rect 167546 547558 167782 547794
rect 167866 547558 168102 547794
rect 171266 549718 171502 549954
rect 171586 549718 171822 549954
rect 171266 549398 171502 549634
rect 171586 549398 171822 549634
rect 174986 553438 175222 553674
rect 175306 553438 175542 553674
rect 174986 553118 175222 553354
rect 175306 553118 175542 553354
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 544158 200062 544394
rect 200146 544158 200382 544394
rect 199826 543838 200062 544074
rect 200146 543838 200382 544074
rect 203546 547878 203782 548114
rect 203866 547878 204102 548114
rect 203546 547558 203782 547794
rect 203866 547558 204102 547794
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 549718 207502 549954
rect 207586 549718 207822 549954
rect 207266 549398 207502 549634
rect 207586 549398 207822 549634
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 224250 615218 224486 615454
rect 224250 614898 224486 615134
rect 254970 615218 255206 615454
rect 254970 614898 255206 615134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 239610 597218 239846 597454
rect 239610 596898 239846 597134
rect 270330 597218 270566 597454
rect 270330 596898 270566 597134
rect 224250 579218 224486 579454
rect 224250 578898 224486 579134
rect 254970 579218 255206 579454
rect 254970 578898 255206 579134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 553438 211222 553674
rect 211306 553438 211542 553674
rect 210986 553118 211222 553354
rect 211306 553118 211542 553354
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 544158 236062 544394
rect 236146 544158 236382 544394
rect 235826 543838 236062 544074
rect 236146 543838 236382 544074
rect 239546 547878 239782 548114
rect 239866 547878 240102 548114
rect 239546 547558 239782 547794
rect 239866 547558 240102 547794
rect 243266 549718 243502 549954
rect 243586 549718 243822 549954
rect 243266 549398 243502 549634
rect 243586 549398 243822 549634
rect 246986 553438 247222 553674
rect 247306 553438 247542 553674
rect 246986 553118 247222 553354
rect 247306 553118 247542 553354
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 544158 272062 544394
rect 272146 544158 272382 544394
rect 271826 543838 272062 544074
rect 272146 543838 272382 544074
rect 275546 547878 275782 548114
rect 275866 547878 276102 548114
rect 275546 547558 275782 547794
rect 275866 547558 276102 547794
rect 279266 549718 279502 549954
rect 279586 549718 279822 549954
rect 279266 549398 279502 549634
rect 279586 549398 279822 549634
rect 282986 553438 283222 553674
rect 283306 553438 283542 553674
rect 282986 553118 283222 553354
rect 283306 553118 283542 553354
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 79610 525218 79846 525454
rect 79610 524898 79846 525134
rect 110330 525218 110566 525454
rect 110330 524898 110566 525134
rect 141050 525218 141286 525454
rect 141050 524898 141286 525134
rect 171770 525218 172006 525454
rect 171770 524898 172006 525134
rect 202490 525218 202726 525454
rect 202490 524898 202726 525134
rect 233210 525218 233446 525454
rect 233210 524898 233446 525134
rect 263930 525218 264166 525454
rect 263930 524898 264166 525134
rect 294650 525218 294886 525454
rect 294650 524898 294886 525134
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 79610 489218 79846 489454
rect 79610 488898 79846 489134
rect 110330 489218 110566 489454
rect 110330 488898 110566 489134
rect 141050 489218 141286 489454
rect 141050 488898 141286 489134
rect 171770 489218 172006 489454
rect 171770 488898 172006 489134
rect 202490 489218 202726 489454
rect 202490 488898 202726 489134
rect 233210 489218 233446 489454
rect 233210 488898 233446 489134
rect 263930 489218 264166 489454
rect 263930 488898 264166 489134
rect 294650 489218 294886 489454
rect 294650 488898 294886 489134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 473998 59782 474234
rect 59866 473998 60102 474234
rect 59546 473678 59782 473914
rect 59866 473678 60102 473914
rect 63266 469842 63502 470078
rect 63586 469842 63822 470078
rect 63266 469522 63502 469758
rect 63586 469522 63822 469758
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 468902 81502 469138
rect 81586 468902 81822 469138
rect 81266 468582 81502 468818
rect 81586 468582 81822 468818
rect 84986 465318 85222 465554
rect 85306 465318 85542 465554
rect 84986 464998 85222 465234
rect 85306 464998 85542 465234
rect 91826 470278 92062 470514
rect 92146 470278 92382 470514
rect 91826 469958 92062 470194
rect 92146 469958 92382 470194
rect 95546 473998 95782 474234
rect 95866 473998 96102 474234
rect 95546 473678 95782 473914
rect 95866 473678 96102 473914
rect 99266 469842 99502 470078
rect 99586 469842 99822 470078
rect 99266 469522 99502 469758
rect 99586 469522 99822 469758
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 468902 117502 469138
rect 117586 468902 117822 469138
rect 117266 468582 117502 468818
rect 117586 468582 117822 468818
rect 120986 465318 121222 465554
rect 121306 465318 121542 465554
rect 120986 464998 121222 465234
rect 121306 464998 121542 465234
rect 127826 470278 128062 470514
rect 128146 470278 128382 470514
rect 127826 469958 128062 470194
rect 128146 469958 128382 470194
rect 131546 473998 131782 474234
rect 131866 473998 132102 474234
rect 131546 473678 131782 473914
rect 131866 473678 132102 473914
rect 135266 469842 135502 470078
rect 135586 469842 135822 470078
rect 135266 469522 135502 469758
rect 135586 469522 135822 469758
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 468902 153502 469138
rect 153586 468902 153822 469138
rect 153266 468582 153502 468818
rect 153586 468582 153822 468818
rect 156986 465318 157222 465554
rect 157306 465318 157542 465554
rect 156986 464998 157222 465234
rect 157306 464998 157542 465234
rect 163826 470278 164062 470514
rect 164146 470278 164382 470514
rect 163826 469958 164062 470194
rect 164146 469958 164382 470194
rect 167546 473998 167782 474234
rect 167866 473998 168102 474234
rect 167546 473678 167782 473914
rect 167866 473678 168102 473914
rect 171266 469842 171502 470078
rect 171586 469842 171822 470078
rect 171266 469522 171502 469758
rect 171586 469522 171822 469758
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 468902 189502 469138
rect 189586 468902 189822 469138
rect 189266 468582 189502 468818
rect 189586 468582 189822 468818
rect 192986 465318 193222 465554
rect 193306 465318 193542 465554
rect 192986 464998 193222 465234
rect 193306 464998 193542 465234
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 61008 399218 61244 399454
rect 61008 398898 61244 399134
rect 195376 399218 195612 399454
rect 195376 398898 195612 399134
rect 60328 381218 60564 381454
rect 60328 380898 60564 381134
rect 196056 381218 196292 381454
rect 196056 380898 196292 381134
rect 59546 365998 59782 366234
rect 59866 365998 60102 366234
rect 59546 365678 59782 365914
rect 59866 365678 60102 365914
rect 63266 369718 63502 369954
rect 63586 369718 63822 369954
rect 63266 369398 63502 369634
rect 63586 369398 63822 369634
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 84986 357318 85222 357554
rect 85306 357318 85542 357554
rect 84986 356998 85222 357234
rect 85306 356998 85542 357234
rect 91826 364158 92062 364394
rect 92146 364158 92382 364394
rect 91826 363838 92062 364074
rect 92146 363838 92382 364074
rect 95546 365998 95782 366234
rect 95866 365998 96102 366234
rect 95546 365678 95782 365914
rect 95866 365678 96102 365914
rect 99266 369718 99502 369954
rect 99586 369718 99822 369954
rect 99266 369398 99502 369634
rect 99586 369398 99822 369634
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 357318 121222 357554
rect 121306 357318 121542 357554
rect 120986 356998 121222 357234
rect 121306 356998 121542 357234
rect 127826 364158 128062 364394
rect 128146 364158 128382 364394
rect 127826 363838 128062 364074
rect 128146 363838 128382 364074
rect 131546 365998 131782 366234
rect 131866 365998 132102 366234
rect 131546 365678 131782 365914
rect 131866 365678 132102 365914
rect 135266 369718 135502 369954
rect 135586 369718 135822 369954
rect 135266 369398 135502 369634
rect 135586 369398 135822 369634
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 156986 357318 157222 357554
rect 157306 357318 157542 357554
rect 156986 356998 157222 357234
rect 157306 356998 157542 357234
rect 163826 364158 164062 364394
rect 164146 364158 164382 364394
rect 163826 363838 164062 364074
rect 164146 363838 164382 364074
rect 167546 365998 167782 366234
rect 167866 365998 168102 366234
rect 167546 365678 167782 365914
rect 167866 365678 168102 365914
rect 171266 369718 171502 369954
rect 171586 369718 171822 369954
rect 171266 369398 171502 369634
rect 171586 369398 171822 369634
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 192986 357318 193222 357554
rect 193306 357318 193542 357554
rect 192986 356998 193222 357234
rect 193306 356998 193542 357234
rect 60328 345218 60564 345454
rect 60328 344898 60564 345134
rect 196056 345218 196292 345454
rect 196056 344898 196292 345134
rect 61008 327218 61244 327454
rect 61008 326898 61244 327134
rect 195376 327218 195612 327454
rect 195376 326898 195612 327134
rect 60328 309218 60564 309454
rect 60328 308898 60564 309134
rect 196056 309218 196292 309454
rect 196056 308898 196292 309134
rect 61008 291218 61244 291454
rect 61008 290898 61244 291134
rect 195376 291218 195612 291454
rect 195376 290898 195612 291134
rect 60328 273218 60564 273454
rect 60328 272898 60564 273134
rect 196056 273218 196292 273454
rect 196056 272898 196292 273134
rect 59546 259878 59782 260114
rect 59866 259878 60102 260114
rect 59546 259558 59782 259794
rect 59866 259558 60102 259794
rect 63266 261718 63502 261954
rect 63586 261718 63822 261954
rect 63266 261398 63502 261634
rect 63586 261398 63822 261634
rect 66986 265438 67222 265674
rect 67306 265438 67542 265674
rect 66986 265118 67222 265354
rect 67306 265118 67542 265354
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 91826 256158 92062 256394
rect 92146 256158 92382 256394
rect 91826 255838 92062 256074
rect 92146 255838 92382 256074
rect 95546 259878 95782 260114
rect 95866 259878 96102 260114
rect 95546 259558 95782 259794
rect 95866 259558 96102 259794
rect 99266 261718 99502 261954
rect 99586 261718 99822 261954
rect 99266 261398 99502 261634
rect 99586 261398 99822 261634
rect 102986 265438 103222 265674
rect 103306 265438 103542 265674
rect 102986 265118 103222 265354
rect 103306 265118 103542 265354
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 127826 256158 128062 256394
rect 128146 256158 128382 256394
rect 127826 255838 128062 256074
rect 128146 255838 128382 256074
rect 131546 259878 131782 260114
rect 131866 259878 132102 260114
rect 131546 259558 131782 259794
rect 131866 259558 132102 259794
rect 135266 261718 135502 261954
rect 135586 261718 135822 261954
rect 135266 261398 135502 261634
rect 135586 261398 135822 261634
rect 138986 265438 139222 265674
rect 139306 265438 139542 265674
rect 138986 265118 139222 265354
rect 139306 265118 139542 265354
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 256158 164062 256394
rect 164146 256158 164382 256394
rect 163826 255838 164062 256074
rect 164146 255838 164382 256074
rect 167546 259878 167782 260114
rect 167866 259878 168102 260114
rect 167546 259558 167782 259794
rect 167866 259558 168102 259794
rect 171266 261718 171502 261954
rect 171586 261718 171822 261954
rect 171266 261398 171502 261634
rect 171586 261398 171822 261634
rect 174986 265438 175222 265674
rect 175306 265438 175542 265674
rect 174986 265118 175222 265354
rect 175306 265118 175542 265354
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 60328 237218 60564 237454
rect 60328 236898 60564 237134
rect 196056 237218 196292 237454
rect 196056 236898 196292 237134
rect 61008 219218 61244 219454
rect 61008 218898 61244 219134
rect 195376 219218 195612 219454
rect 195376 218898 195612 219134
rect 60328 201218 60564 201454
rect 60328 200898 60564 201134
rect 196056 201218 196292 201454
rect 196056 200898 196292 201134
rect 61008 183218 61244 183454
rect 61008 182898 61244 183134
rect 195376 183218 195612 183454
rect 195376 182898 195612 183134
rect 59546 151878 59782 152114
rect 59866 151878 60102 152114
rect 59546 151558 59782 151794
rect 59866 151558 60102 151794
rect 63266 153718 63502 153954
rect 63586 153718 63822 153954
rect 63266 153398 63502 153634
rect 63586 153398 63822 153634
rect 66986 157438 67222 157674
rect 67306 157438 67542 157674
rect 66986 157118 67222 157354
rect 67306 157118 67542 157354
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 148158 92062 148394
rect 92146 148158 92382 148394
rect 91826 147838 92062 148074
rect 92146 147838 92382 148074
rect 95546 151878 95782 152114
rect 95866 151878 96102 152114
rect 95546 151558 95782 151794
rect 95866 151558 96102 151794
rect 99266 153718 99502 153954
rect 99586 153718 99822 153954
rect 99266 153398 99502 153634
rect 99586 153398 99822 153634
rect 102986 157438 103222 157674
rect 103306 157438 103542 157674
rect 102986 157118 103222 157354
rect 103306 157118 103542 157354
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 127826 148158 128062 148394
rect 128146 148158 128382 148394
rect 127826 147838 128062 148074
rect 128146 147838 128382 148074
rect 131546 151878 131782 152114
rect 131866 151878 132102 152114
rect 131546 151558 131782 151794
rect 131866 151558 132102 151794
rect 135266 153718 135502 153954
rect 135586 153718 135822 153954
rect 135266 153398 135502 153634
rect 135586 153398 135822 153634
rect 138986 157438 139222 157674
rect 139306 157438 139542 157674
rect 138986 157118 139222 157354
rect 139306 157118 139542 157354
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 163826 148158 164062 148394
rect 164146 148158 164382 148394
rect 163826 147838 164062 148074
rect 164146 147838 164382 148074
rect 167546 151878 167782 152114
rect 167866 151878 168102 152114
rect 167546 151558 167782 151794
rect 167866 151558 168102 151794
rect 171266 153718 171502 153954
rect 171586 153718 171822 153954
rect 171266 153398 171502 153634
rect 171586 153398 171822 153634
rect 174986 157438 175222 157674
rect 175306 157438 175542 157674
rect 174986 157118 175222 157354
rect 175306 157118 175542 157354
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 60328 129218 60564 129454
rect 60328 128898 60564 129134
rect 196056 129218 196292 129454
rect 196056 128898 196292 129134
rect 61008 111218 61244 111454
rect 61008 110898 61244 111134
rect 195376 111218 195612 111454
rect 195376 110898 195612 111134
rect 60328 93218 60564 93454
rect 60328 92898 60564 93134
rect 196056 93218 196292 93454
rect 196056 92898 196292 93134
rect 61008 75218 61244 75454
rect 61008 74898 61244 75134
rect 195376 75218 195612 75454
rect 195376 74898 195612 75134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 199826 470278 200062 470514
rect 200146 470278 200382 470514
rect 199826 469958 200062 470194
rect 200146 469958 200382 470194
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 364158 200062 364394
rect 200146 364158 200382 364394
rect 199826 363838 200062 364074
rect 200146 363838 200382 364074
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 256158 200062 256394
rect 200146 256158 200382 256394
rect 199826 255838 200062 256074
rect 200146 255838 200382 256074
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 148158 200062 148394
rect 200146 148158 200382 148394
rect 199826 147838 200062 148074
rect 200146 147838 200382 148074
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 203546 473998 203782 474234
rect 203866 473998 204102 474234
rect 203546 473678 203782 473914
rect 203866 473678 204102 473914
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 365998 203782 366234
rect 203866 365998 204102 366234
rect 203546 365678 203782 365914
rect 203866 365678 204102 365914
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 259878 203782 260114
rect 203866 259878 204102 260114
rect 203546 259558 203782 259794
rect 203866 259558 204102 259794
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 151878 203782 152114
rect 203866 151878 204102 152114
rect 203546 151558 203782 151794
rect 203866 151558 204102 151794
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 207266 469842 207502 470078
rect 207586 469842 207822 470078
rect 207266 469522 207502 469758
rect 207586 469522 207822 469758
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 369718 207502 369954
rect 207586 369718 207822 369954
rect 207266 369398 207502 369634
rect 207586 369398 207822 369634
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 261718 207502 261954
rect 207586 261718 207822 261954
rect 207266 261398 207502 261634
rect 207586 261398 207822 261634
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 153718 207502 153954
rect 207586 153718 207822 153954
rect 207266 153398 207502 153634
rect 207586 153398 207822 153634
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 265438 211222 265674
rect 211306 265438 211542 265674
rect 210986 265118 211222 265354
rect 211306 265118 211542 265354
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 157438 211222 157674
rect 211306 157438 211542 157674
rect 210986 157118 211222 157354
rect 211306 157118 211542 157354
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 468902 225502 469138
rect 225586 468902 225822 469138
rect 225266 468582 225502 468818
rect 225586 468582 225822 468818
rect 228986 465318 229222 465554
rect 229306 465318 229542 465554
rect 228986 464998 229222 465234
rect 229306 464998 229542 465234
rect 235826 470278 236062 470514
rect 236146 470278 236382 470514
rect 235826 469958 236062 470194
rect 236146 469958 236382 470194
rect 239546 473998 239782 474234
rect 239866 473998 240102 474234
rect 239546 473678 239782 473914
rect 239866 473678 240102 473914
rect 243266 469842 243502 470078
rect 243586 469842 243822 470078
rect 243266 469522 243502 469758
rect 243586 469522 243822 469758
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 468902 261502 469138
rect 261586 468902 261822 469138
rect 261266 468582 261502 468818
rect 261586 468582 261822 468818
rect 264986 465318 265222 465554
rect 265306 465318 265542 465554
rect 264986 464998 265222 465234
rect 265306 464998 265542 465234
rect 271826 470278 272062 470514
rect 272146 470278 272382 470514
rect 271826 469958 272062 470194
rect 272146 469958 272382 470194
rect 275546 473998 275782 474234
rect 275866 473998 276102 474234
rect 275546 473678 275782 473914
rect 275866 473678 276102 473914
rect 279266 469842 279502 470078
rect 279586 469842 279822 470078
rect 279266 469522 279502 469758
rect 279586 469522 279822 469758
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 468902 297502 469138
rect 297586 468902 297822 469138
rect 297266 468582 297502 468818
rect 297586 468582 297822 468818
rect 300986 465318 301222 465554
rect 301306 465318 301542 465554
rect 300986 464998 301222 465234
rect 301306 464998 301542 465234
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 324250 615218 324486 615454
rect 324250 614898 324486 615134
rect 354970 615218 355206 615454
rect 354970 614898 355206 615134
rect 385690 615218 385926 615454
rect 385690 614898 385926 615134
rect 416410 615218 416646 615454
rect 416410 614898 416646 615134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 339610 597218 339846 597454
rect 339610 596898 339846 597134
rect 370330 597218 370566 597454
rect 370330 596898 370566 597134
rect 401050 597218 401286 597454
rect 401050 596898 401286 597134
rect 324250 579218 324486 579454
rect 324250 578898 324486 579134
rect 354970 579218 355206 579454
rect 354970 578898 355206 579134
rect 385690 579218 385926 579454
rect 385690 578898 385926 579134
rect 416410 579218 416646 579454
rect 416410 578898 416646 579134
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 339610 561218 339846 561454
rect 339610 560898 339846 561134
rect 370330 561218 370566 561454
rect 370330 560898 370566 561134
rect 401050 561218 401286 561454
rect 401050 560898 401286 561134
rect 324250 543218 324486 543454
rect 324250 542898 324486 543134
rect 354970 543218 355206 543454
rect 354970 542898 355206 543134
rect 385690 543218 385926 543454
rect 385690 542898 385926 543134
rect 416410 543218 416646 543454
rect 416410 542898 416646 543134
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 339610 525218 339846 525454
rect 339610 524898 339846 525134
rect 370330 525218 370566 525454
rect 370330 524898 370566 525134
rect 401050 525218 401286 525454
rect 401050 524898 401286 525134
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221008 399218 221244 399454
rect 221008 398898 221244 399134
rect 355376 399218 355612 399454
rect 355376 398898 355612 399134
rect 220328 381218 220564 381454
rect 220328 380898 220564 381134
rect 356056 381218 356292 381454
rect 356056 380898 356292 381134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 228986 357318 229222 357554
rect 229306 357318 229542 357554
rect 228986 356998 229222 357234
rect 229306 356998 229542 357234
rect 235826 364158 236062 364394
rect 236146 364158 236382 364394
rect 235826 363838 236062 364074
rect 236146 363838 236382 364074
rect 239546 365998 239782 366234
rect 239866 365998 240102 366234
rect 239546 365678 239782 365914
rect 239866 365678 240102 365914
rect 243266 369718 243502 369954
rect 243586 369718 243822 369954
rect 243266 369398 243502 369634
rect 243586 369398 243822 369634
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 264986 357318 265222 357554
rect 265306 357318 265542 357554
rect 264986 356998 265222 357234
rect 265306 356998 265542 357234
rect 271826 364158 272062 364394
rect 272146 364158 272382 364394
rect 271826 363838 272062 364074
rect 272146 363838 272382 364074
rect 275546 365998 275782 366234
rect 275866 365998 276102 366234
rect 275546 365678 275782 365914
rect 275866 365678 276102 365914
rect 279266 369718 279502 369954
rect 279586 369718 279822 369954
rect 279266 369398 279502 369634
rect 279586 369398 279822 369634
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 300986 357318 301222 357554
rect 301306 357318 301542 357554
rect 300986 356998 301222 357234
rect 301306 356998 301542 357234
rect 307826 364158 308062 364394
rect 308146 364158 308382 364394
rect 307826 363838 308062 364074
rect 308146 363838 308382 364074
rect 311546 365998 311782 366234
rect 311866 365998 312102 366234
rect 311546 365678 311782 365914
rect 311866 365678 312102 365914
rect 315266 369718 315502 369954
rect 315586 369718 315822 369954
rect 315266 369398 315502 369634
rect 315586 369398 315822 369634
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 336986 357318 337222 357554
rect 337306 357318 337542 357554
rect 336986 356998 337222 357234
rect 337306 356998 337542 357234
rect 343826 364158 344062 364394
rect 344146 364158 344382 364394
rect 343826 363838 344062 364074
rect 344146 363838 344382 364074
rect 347546 365998 347782 366234
rect 347866 365998 348102 366234
rect 347546 365678 347782 365914
rect 347866 365678 348102 365914
rect 351266 369718 351502 369954
rect 351586 369718 351822 369954
rect 351266 369398 351502 369634
rect 351586 369398 351822 369634
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 220328 345218 220564 345454
rect 220328 344898 220564 345134
rect 356056 345218 356292 345454
rect 356056 344898 356292 345134
rect 221008 327218 221244 327454
rect 221008 326898 221244 327134
rect 355376 327218 355612 327454
rect 355376 326898 355612 327134
rect 220328 309218 220564 309454
rect 220328 308898 220564 309134
rect 356056 309218 356292 309454
rect 356056 308898 356292 309134
rect 221008 291218 221244 291454
rect 221008 290898 221244 291134
rect 355376 291218 355612 291454
rect 355376 290898 355612 291134
rect 220328 273218 220564 273454
rect 220328 272898 220564 273134
rect 356056 273218 356292 273454
rect 356056 272898 356292 273134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 235826 256158 236062 256394
rect 236146 256158 236382 256394
rect 235826 255838 236062 256074
rect 236146 255838 236382 256074
rect 239546 259878 239782 260114
rect 239866 259878 240102 260114
rect 239546 259558 239782 259794
rect 239866 259558 240102 259794
rect 243266 261718 243502 261954
rect 243586 261718 243822 261954
rect 243266 261398 243502 261634
rect 243586 261398 243822 261634
rect 246986 265438 247222 265674
rect 247306 265438 247542 265674
rect 246986 265118 247222 265354
rect 247306 265118 247542 265354
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 271826 256158 272062 256394
rect 272146 256158 272382 256394
rect 271826 255838 272062 256074
rect 272146 255838 272382 256074
rect 275546 259878 275782 260114
rect 275866 259878 276102 260114
rect 275546 259558 275782 259794
rect 275866 259558 276102 259794
rect 279266 261718 279502 261954
rect 279586 261718 279822 261954
rect 279266 261398 279502 261634
rect 279586 261398 279822 261634
rect 282986 265438 283222 265674
rect 283306 265438 283542 265674
rect 282986 265118 283222 265354
rect 283306 265118 283542 265354
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 307826 256158 308062 256394
rect 308146 256158 308382 256394
rect 307826 255838 308062 256074
rect 308146 255838 308382 256074
rect 311546 259878 311782 260114
rect 311866 259878 312102 260114
rect 311546 259558 311782 259794
rect 311866 259558 312102 259794
rect 315266 261718 315502 261954
rect 315586 261718 315822 261954
rect 315266 261398 315502 261634
rect 315586 261398 315822 261634
rect 318986 265438 319222 265674
rect 319306 265438 319542 265674
rect 318986 265118 319222 265354
rect 319306 265118 319542 265354
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 343826 256158 344062 256394
rect 344146 256158 344382 256394
rect 343826 255838 344062 256074
rect 344146 255838 344382 256074
rect 347546 259878 347782 260114
rect 347866 259878 348102 260114
rect 347546 259558 347782 259794
rect 347866 259558 348102 259794
rect 351266 261718 351502 261954
rect 351586 261718 351822 261954
rect 351266 261398 351502 261634
rect 351586 261398 351822 261634
rect 354986 265438 355222 265674
rect 355306 265438 355542 265674
rect 354986 265118 355222 265354
rect 355306 265118 355542 265354
rect 220328 237218 220564 237454
rect 220328 236898 220564 237134
rect 356056 237218 356292 237454
rect 356056 236898 356292 237134
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 201218 220564 201454
rect 220328 200898 220564 201134
rect 356056 201218 356292 201454
rect 356056 200898 356292 201134
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 235826 148158 236062 148394
rect 236146 148158 236382 148394
rect 235826 147838 236062 148074
rect 236146 147838 236382 148074
rect 239546 151878 239782 152114
rect 239866 151878 240102 152114
rect 239546 151558 239782 151794
rect 239866 151558 240102 151794
rect 243266 153718 243502 153954
rect 243586 153718 243822 153954
rect 243266 153398 243502 153634
rect 243586 153398 243822 153634
rect 246986 157438 247222 157674
rect 247306 157438 247542 157674
rect 246986 157118 247222 157354
rect 247306 157118 247542 157354
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 271826 148158 272062 148394
rect 272146 148158 272382 148394
rect 271826 147838 272062 148074
rect 272146 147838 272382 148074
rect 275546 151878 275782 152114
rect 275866 151878 276102 152114
rect 275546 151558 275782 151794
rect 275866 151558 276102 151794
rect 279266 153718 279502 153954
rect 279586 153718 279822 153954
rect 279266 153398 279502 153634
rect 279586 153398 279822 153634
rect 282986 157438 283222 157674
rect 283306 157438 283542 157674
rect 282986 157118 283222 157354
rect 283306 157118 283542 157354
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 307826 148158 308062 148394
rect 308146 148158 308382 148394
rect 307826 147838 308062 148074
rect 308146 147838 308382 148074
rect 311546 151878 311782 152114
rect 311866 151878 312102 152114
rect 311546 151558 311782 151794
rect 311866 151558 312102 151794
rect 315266 153718 315502 153954
rect 315586 153718 315822 153954
rect 315266 153398 315502 153634
rect 315586 153398 315822 153634
rect 318986 157438 319222 157674
rect 319306 157438 319542 157674
rect 318986 157118 319222 157354
rect 319306 157118 319542 157354
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 343826 148158 344062 148394
rect 344146 148158 344382 148394
rect 343826 147838 344062 148074
rect 344146 147838 344382 148074
rect 347546 151878 347782 152114
rect 347866 151878 348102 152114
rect 347546 151558 347782 151794
rect 347866 151558 348102 151794
rect 351266 153718 351502 153954
rect 351586 153718 351822 153954
rect 351266 153398 351502 153634
rect 351586 153398 351822 153634
rect 354986 157438 355222 157674
rect 355306 157438 355542 157674
rect 354986 157118 355222 157354
rect 355306 157118 355542 157354
rect 220328 129218 220564 129454
rect 220328 128898 220564 129134
rect 356056 129218 356292 129454
rect 356056 128898 356292 129134
rect 221008 111218 221244 111454
rect 221008 110898 221244 111134
rect 355376 111218 355612 111454
rect 355376 110898 355612 111134
rect 220328 93218 220564 93454
rect 220328 92898 220564 93134
rect 356056 93218 356292 93454
rect 356056 92898 356292 93134
rect 221008 75218 221244 75454
rect 221008 74898 221244 75134
rect 355376 75218 355612 75454
rect 355376 74898 355612 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 357318 373222 357554
rect 373306 357318 373542 357554
rect 372986 356998 373222 357234
rect 373306 356998 373542 357234
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 479610 597218 479846 597454
rect 479610 596898 479846 597134
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 464250 579218 464486 579454
rect 464250 578898 464486 579134
rect 494970 579218 495206 579454
rect 494970 578898 495206 579134
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 380328 453218 380564 453454
rect 380328 452898 380564 453134
rect 516056 453218 516292 453454
rect 516056 452898 516292 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 381008 435218 381244 435454
rect 381008 434898 381244 435134
rect 515376 435218 515612 435454
rect 515376 434898 515612 435134
rect 380328 417218 380564 417454
rect 380328 416898 380564 417134
rect 516056 417218 516292 417454
rect 516056 416898 516292 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 381008 399218 381244 399454
rect 381008 398898 381244 399134
rect 515376 399218 515612 399454
rect 515376 398898 515612 399134
rect 380328 381218 380564 381454
rect 380328 380898 380564 381134
rect 516056 381218 516292 381454
rect 516056 380898 516292 381134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 379826 364158 380062 364394
rect 380146 364158 380382 364394
rect 379826 363838 380062 364074
rect 380146 363838 380382 364074
rect 383546 365998 383782 366234
rect 383866 365998 384102 366234
rect 383546 365678 383782 365914
rect 383866 365678 384102 365914
rect 387266 369718 387502 369954
rect 387586 369718 387822 369954
rect 387266 369398 387502 369634
rect 387586 369398 387822 369634
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 408986 357318 409222 357554
rect 409306 357318 409542 357554
rect 408986 356998 409222 357234
rect 409306 356998 409542 357234
rect 415826 364158 416062 364394
rect 416146 364158 416382 364394
rect 415826 363838 416062 364074
rect 416146 363838 416382 364074
rect 419546 365998 419782 366234
rect 419866 365998 420102 366234
rect 419546 365678 419782 365914
rect 419866 365678 420102 365914
rect 423266 369718 423502 369954
rect 423586 369718 423822 369954
rect 423266 369398 423502 369634
rect 423586 369398 423822 369634
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 444986 357318 445222 357554
rect 445306 357318 445542 357554
rect 444986 356998 445222 357234
rect 445306 356998 445542 357234
rect 451826 364158 452062 364394
rect 452146 364158 452382 364394
rect 451826 363838 452062 364074
rect 452146 363838 452382 364074
rect 455546 365998 455782 366234
rect 455866 365998 456102 366234
rect 455546 365678 455782 365914
rect 455866 365678 456102 365914
rect 459266 369718 459502 369954
rect 459586 369718 459822 369954
rect 459266 369398 459502 369634
rect 459586 369398 459822 369634
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 480986 357318 481222 357554
rect 481306 357318 481542 357554
rect 480986 356998 481222 357234
rect 481306 356998 481542 357234
rect 487826 364158 488062 364394
rect 488146 364158 488382 364394
rect 487826 363838 488062 364074
rect 488146 363838 488382 364074
rect 491546 365998 491782 366234
rect 491866 365998 492102 366234
rect 491546 365678 491782 365914
rect 491866 365678 492102 365914
rect 495266 369718 495502 369954
rect 495586 369718 495822 369954
rect 495266 369398 495502 369634
rect 495586 369398 495822 369634
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 516986 357318 517222 357554
rect 517306 357318 517542 357554
rect 516986 356998 517222 357234
rect 517306 356998 517542 357234
rect 380328 345218 380564 345454
rect 380328 344898 380564 345134
rect 516056 345218 516292 345454
rect 516056 344898 516292 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 381008 327218 381244 327454
rect 381008 326898 381244 327134
rect 515376 327218 515612 327454
rect 515376 326898 515612 327134
rect 380328 309218 380564 309454
rect 380328 308898 380564 309134
rect 516056 309218 516292 309454
rect 516056 308898 516292 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 381008 291218 381244 291454
rect 381008 290898 381244 291134
rect 515376 291218 515612 291454
rect 515376 290898 515612 291134
rect 380328 273218 380564 273454
rect 380328 272898 380564 273134
rect 516056 273218 516292 273454
rect 516056 272898 516292 273134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 379826 256158 380062 256394
rect 380146 256158 380382 256394
rect 379826 255838 380062 256074
rect 380146 255838 380382 256074
rect 383546 259878 383782 260114
rect 383866 259878 384102 260114
rect 383546 259558 383782 259794
rect 383866 259558 384102 259794
rect 387266 261718 387502 261954
rect 387586 261718 387822 261954
rect 387266 261398 387502 261634
rect 387586 261398 387822 261634
rect 390986 265438 391222 265674
rect 391306 265438 391542 265674
rect 390986 265118 391222 265354
rect 391306 265118 391542 265354
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 415826 256158 416062 256394
rect 416146 256158 416382 256394
rect 415826 255838 416062 256074
rect 416146 255838 416382 256074
rect 419546 259878 419782 260114
rect 419866 259878 420102 260114
rect 419546 259558 419782 259794
rect 419866 259558 420102 259794
rect 423266 261718 423502 261954
rect 423586 261718 423822 261954
rect 423266 261398 423502 261634
rect 423586 261398 423822 261634
rect 426986 265438 427222 265674
rect 427306 265438 427542 265674
rect 426986 265118 427222 265354
rect 427306 265118 427542 265354
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 451826 256158 452062 256394
rect 452146 256158 452382 256394
rect 451826 255838 452062 256074
rect 452146 255838 452382 256074
rect 455546 259878 455782 260114
rect 455866 259878 456102 260114
rect 455546 259558 455782 259794
rect 455866 259558 456102 259794
rect 459266 261718 459502 261954
rect 459586 261718 459822 261954
rect 459266 261398 459502 261634
rect 459586 261398 459822 261634
rect 462986 265438 463222 265674
rect 463306 265438 463542 265674
rect 462986 265118 463222 265354
rect 463306 265118 463542 265354
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 487826 256158 488062 256394
rect 488146 256158 488382 256394
rect 487826 255838 488062 256074
rect 488146 255838 488382 256074
rect 491546 259878 491782 260114
rect 491866 259878 492102 260114
rect 491546 259558 491782 259794
rect 491866 259558 492102 259794
rect 495266 261718 495502 261954
rect 495586 261718 495822 261954
rect 495266 261398 495502 261634
rect 495586 261398 495822 261634
rect 498986 265438 499222 265674
rect 499306 265438 499542 265674
rect 498986 265118 499222 265354
rect 499306 265118 499542 265354
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 380328 237218 380564 237454
rect 380328 236898 380564 237134
rect 516056 237218 516292 237454
rect 516056 236898 516292 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 381008 219218 381244 219454
rect 381008 218898 381244 219134
rect 515376 219218 515612 219454
rect 515376 218898 515612 219134
rect 380328 201218 380564 201454
rect 380328 200898 380564 201134
rect 516056 201218 516292 201454
rect 516056 200898 516292 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 381008 183218 381244 183454
rect 381008 182898 381244 183134
rect 515376 183218 515612 183454
rect 515376 182898 515612 183134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 379826 148158 380062 148394
rect 380146 148158 380382 148394
rect 379826 147838 380062 148074
rect 380146 147838 380382 148074
rect 383546 151878 383782 152114
rect 383866 151878 384102 152114
rect 383546 151558 383782 151794
rect 383866 151558 384102 151794
rect 387266 153718 387502 153954
rect 387586 153718 387822 153954
rect 387266 153398 387502 153634
rect 387586 153398 387822 153634
rect 390986 157438 391222 157674
rect 391306 157438 391542 157674
rect 390986 157118 391222 157354
rect 391306 157118 391542 157354
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 415826 148158 416062 148394
rect 416146 148158 416382 148394
rect 415826 147838 416062 148074
rect 416146 147838 416382 148074
rect 419546 151878 419782 152114
rect 419866 151878 420102 152114
rect 419546 151558 419782 151794
rect 419866 151558 420102 151794
rect 423266 153718 423502 153954
rect 423586 153718 423822 153954
rect 423266 153398 423502 153634
rect 423586 153398 423822 153634
rect 426986 157438 427222 157674
rect 427306 157438 427542 157674
rect 426986 157118 427222 157354
rect 427306 157118 427542 157354
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 148158 452062 148394
rect 452146 148158 452382 148394
rect 451826 147838 452062 148074
rect 452146 147838 452382 148074
rect 455546 151878 455782 152114
rect 455866 151878 456102 152114
rect 455546 151558 455782 151794
rect 455866 151558 456102 151794
rect 459266 153718 459502 153954
rect 459586 153718 459822 153954
rect 459266 153398 459502 153634
rect 459586 153398 459822 153634
rect 462986 157438 463222 157674
rect 463306 157438 463542 157674
rect 462986 157118 463222 157354
rect 463306 157118 463542 157354
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 148158 488062 148394
rect 488146 148158 488382 148394
rect 487826 147838 488062 148074
rect 488146 147838 488382 148074
rect 491546 151878 491782 152114
rect 491866 151878 492102 152114
rect 491546 151558 491782 151794
rect 491866 151558 492102 151794
rect 495266 153718 495502 153954
rect 495586 153718 495822 153954
rect 495266 153398 495502 153634
rect 495586 153398 495822 153634
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 498986 157438 499222 157674
rect 499306 157438 499542 157674
rect 498986 157118 499222 157354
rect 499306 157118 499542 157354
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 380328 129218 380564 129454
rect 380328 128898 380564 129134
rect 516056 129218 516292 129454
rect 516056 128898 516292 129134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 381008 111218 381244 111454
rect 381008 110898 381244 111134
rect 515376 111218 515612 111454
rect 515376 110898 515612 111134
rect 380328 93218 380564 93454
rect 380328 92898 380564 93134
rect 516056 93218 516292 93454
rect 516056 92898 516292 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 381008 75218 381244 75454
rect 381008 74898 381244 75134
rect 515376 75218 515612 75454
rect 515376 74898 515612 75134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 144250 615454
rect 144486 615218 174970 615454
rect 175206 615218 224250 615454
rect 224486 615218 254970 615454
rect 255206 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 324250 615454
rect 324486 615218 354970 615454
rect 355206 615218 385690 615454
rect 385926 615218 416410 615454
rect 416646 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 144250 615134
rect 144486 614898 174970 615134
rect 175206 614898 224250 615134
rect 224486 614898 254970 615134
rect 255206 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 324250 615134
rect 324486 614898 354970 615134
rect 355206 614898 385690 615134
rect 385926 614898 416410 615134
rect 416646 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 79610 597454
rect 79846 597218 110330 597454
rect 110566 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 159610 597454
rect 159846 597218 190330 597454
rect 190566 597218 239610 597454
rect 239846 597218 270330 597454
rect 270566 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 339610 597454
rect 339846 597218 370330 597454
rect 370566 597218 401050 597454
rect 401286 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 479610 597454
rect 479846 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 79610 597134
rect 79846 596898 110330 597134
rect 110566 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 159610 597134
rect 159846 596898 190330 597134
rect 190566 596898 239610 597134
rect 239846 596898 270330 597134
rect 270566 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 339610 597134
rect 339846 596898 370330 597134
rect 370566 596898 401050 597134
rect 401286 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 479610 597134
rect 479846 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64250 579454
rect 64486 579218 94970 579454
rect 95206 579218 144250 579454
rect 144486 579218 174970 579454
rect 175206 579218 224250 579454
rect 224486 579218 254970 579454
rect 255206 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 324250 579454
rect 324486 579218 354970 579454
rect 355206 579218 385690 579454
rect 385926 579218 416410 579454
rect 416646 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 464250 579454
rect 464486 579218 494970 579454
rect 495206 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64250 579134
rect 64486 578898 94970 579134
rect 95206 578898 144250 579134
rect 144486 578898 174970 579134
rect 175206 578898 224250 579134
rect 224486 578898 254970 579134
rect 255206 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 324250 579134
rect 324486 578898 354970 579134
rect 355206 578898 385690 579134
rect 385926 578898 416410 579134
rect 416646 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 464250 579134
rect 464486 578898 494970 579134
rect 495206 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 339610 561454
rect 339846 561218 370330 561454
rect 370566 561218 401050 561454
rect 401286 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 339610 561134
rect 339846 560898 370330 561134
rect 370566 560898 401050 561134
rect 401286 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect 66954 553674 283574 553706
rect 66954 553438 66986 553674
rect 67222 553438 67306 553674
rect 67542 553438 102986 553674
rect 103222 553438 103306 553674
rect 103542 553438 138986 553674
rect 139222 553438 139306 553674
rect 139542 553438 174986 553674
rect 175222 553438 175306 553674
rect 175542 553438 210986 553674
rect 211222 553438 211306 553674
rect 211542 553438 246986 553674
rect 247222 553438 247306 553674
rect 247542 553438 282986 553674
rect 283222 553438 283306 553674
rect 283542 553438 283574 553674
rect 66954 553354 283574 553438
rect 66954 553118 66986 553354
rect 67222 553118 67306 553354
rect 67542 553118 102986 553354
rect 103222 553118 103306 553354
rect 103542 553118 138986 553354
rect 139222 553118 139306 553354
rect 139542 553118 174986 553354
rect 175222 553118 175306 553354
rect 175542 553118 210986 553354
rect 211222 553118 211306 553354
rect 211542 553118 246986 553354
rect 247222 553118 247306 553354
rect 247542 553118 282986 553354
rect 283222 553118 283306 553354
rect 283542 553118 283574 553354
rect 66954 553086 283574 553118
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect 63234 549954 279854 549986
rect 63234 549718 63266 549954
rect 63502 549718 63586 549954
rect 63822 549718 99266 549954
rect 99502 549718 99586 549954
rect 99822 549718 135266 549954
rect 135502 549718 135586 549954
rect 135822 549718 171266 549954
rect 171502 549718 171586 549954
rect 171822 549718 207266 549954
rect 207502 549718 207586 549954
rect 207822 549718 243266 549954
rect 243502 549718 243586 549954
rect 243822 549718 279266 549954
rect 279502 549718 279586 549954
rect 279822 549718 279854 549954
rect 63234 549634 279854 549718
rect 63234 549398 63266 549634
rect 63502 549398 63586 549634
rect 63822 549398 99266 549634
rect 99502 549398 99586 549634
rect 99822 549398 135266 549634
rect 135502 549398 135586 549634
rect 135822 549398 171266 549634
rect 171502 549398 171586 549634
rect 171822 549398 207266 549634
rect 207502 549398 207586 549634
rect 207822 549398 243266 549634
rect 243502 549398 243586 549634
rect 243822 549398 279266 549634
rect 279502 549398 279586 549634
rect 279822 549398 279854 549634
rect 63234 549366 279854 549398
rect 59514 548114 276134 548146
rect 59514 547878 59546 548114
rect 59782 547878 59866 548114
rect 60102 547878 95546 548114
rect 95782 547878 95866 548114
rect 96102 547878 131546 548114
rect 131782 547878 131866 548114
rect 132102 547878 167546 548114
rect 167782 547878 167866 548114
rect 168102 547878 203546 548114
rect 203782 547878 203866 548114
rect 204102 547878 239546 548114
rect 239782 547878 239866 548114
rect 240102 547878 275546 548114
rect 275782 547878 275866 548114
rect 276102 547878 276134 548114
rect 59514 547794 276134 547878
rect 59514 547558 59546 547794
rect 59782 547558 59866 547794
rect 60102 547558 95546 547794
rect 95782 547558 95866 547794
rect 96102 547558 131546 547794
rect 131782 547558 131866 547794
rect 132102 547558 167546 547794
rect 167782 547558 167866 547794
rect 168102 547558 203546 547794
rect 203782 547558 203866 547794
rect 204102 547558 239546 547794
rect 239782 547558 239866 547794
rect 240102 547558 275546 547794
rect 275782 547558 275866 547794
rect 276102 547558 276134 547794
rect 59514 547526 276134 547558
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect 91794 544394 272414 544426
rect 91794 544158 91826 544394
rect 92062 544158 92146 544394
rect 92382 544158 127826 544394
rect 128062 544158 128146 544394
rect 128382 544158 163826 544394
rect 164062 544158 164146 544394
rect 164382 544158 199826 544394
rect 200062 544158 200146 544394
rect 200382 544158 235826 544394
rect 236062 544158 236146 544394
rect 236382 544158 271826 544394
rect 272062 544158 272146 544394
rect 272382 544158 272414 544394
rect 91794 544074 272414 544158
rect 91794 543838 91826 544074
rect 92062 543838 92146 544074
rect 92382 543838 127826 544074
rect 128062 543838 128146 544074
rect 128382 543838 163826 544074
rect 164062 543838 164146 544074
rect 164382 543838 199826 544074
rect 200062 543838 200146 544074
rect 200382 543838 235826 544074
rect 236062 543838 236146 544074
rect 236382 543838 271826 544074
rect 272062 543838 272146 544074
rect 272382 543838 272414 544074
rect 91794 543806 272414 543838
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 324250 543454
rect 324486 543218 354970 543454
rect 355206 543218 385690 543454
rect 385926 543218 416410 543454
rect 416646 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 324250 543134
rect 324486 542898 354970 543134
rect 355206 542898 385690 543134
rect 385926 542898 416410 543134
rect 416646 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 79610 525454
rect 79846 525218 110330 525454
rect 110566 525218 141050 525454
rect 141286 525218 171770 525454
rect 172006 525218 202490 525454
rect 202726 525218 233210 525454
rect 233446 525218 263930 525454
rect 264166 525218 294650 525454
rect 294886 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 339610 525454
rect 339846 525218 370330 525454
rect 370566 525218 401050 525454
rect 401286 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 79610 525134
rect 79846 524898 110330 525134
rect 110566 524898 141050 525134
rect 141286 524898 171770 525134
rect 172006 524898 202490 525134
rect 202726 524898 233210 525134
rect 233446 524898 263930 525134
rect 264166 524898 294650 525134
rect 294886 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 339610 525134
rect 339846 524898 370330 525134
rect 370566 524898 401050 525134
rect 401286 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 79610 489454
rect 79846 489218 110330 489454
rect 110566 489218 141050 489454
rect 141286 489218 171770 489454
rect 172006 489218 202490 489454
rect 202726 489218 233210 489454
rect 233446 489218 263930 489454
rect 264166 489218 294650 489454
rect 294886 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 79610 489134
rect 79846 488898 110330 489134
rect 110566 488898 141050 489134
rect 141286 488898 171770 489134
rect 172006 488898 202490 489134
rect 202726 488898 233210 489134
rect 233446 488898 263930 489134
rect 264166 488898 294650 489134
rect 294886 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect 59514 474234 276134 474266
rect 59514 473998 59546 474234
rect 59782 473998 59866 474234
rect 60102 473998 95546 474234
rect 95782 473998 95866 474234
rect 96102 473998 131546 474234
rect 131782 473998 131866 474234
rect 132102 473998 167546 474234
rect 167782 473998 167866 474234
rect 168102 473998 203546 474234
rect 203782 473998 203866 474234
rect 204102 473998 239546 474234
rect 239782 473998 239866 474234
rect 240102 473998 275546 474234
rect 275782 473998 275866 474234
rect 276102 473998 276134 474234
rect 59514 473914 276134 473998
rect 59514 473678 59546 473914
rect 59782 473678 59866 473914
rect 60102 473678 95546 473914
rect 95782 473678 95866 473914
rect 96102 473678 131546 473914
rect 131782 473678 131866 473914
rect 132102 473678 167546 473914
rect 167782 473678 167866 473914
rect 168102 473678 203546 473914
rect 203782 473678 203866 473914
rect 204102 473678 239546 473914
rect 239782 473678 239866 473914
rect 240102 473678 275546 473914
rect 275782 473678 275866 473914
rect 276102 473678 276134 473914
rect 59514 473646 276134 473678
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect 91794 470514 272414 470546
rect 91794 470278 91826 470514
rect 92062 470278 92146 470514
rect 92382 470278 127826 470514
rect 128062 470278 128146 470514
rect 128382 470278 163826 470514
rect 164062 470278 164146 470514
rect 164382 470278 199826 470514
rect 200062 470278 200146 470514
rect 200382 470278 235826 470514
rect 236062 470278 236146 470514
rect 236382 470278 271826 470514
rect 272062 470278 272146 470514
rect 272382 470278 272414 470514
rect 91794 470194 272414 470278
rect 91794 470110 91826 470194
rect 63234 470078 91826 470110
rect 63234 469842 63266 470078
rect 63502 469842 63586 470078
rect 63822 469958 91826 470078
rect 92062 469958 92146 470194
rect 92382 470078 127826 470194
rect 92382 469958 99266 470078
rect 63822 469842 99266 469958
rect 99502 469842 99586 470078
rect 99822 469958 127826 470078
rect 128062 469958 128146 470194
rect 128382 470078 163826 470194
rect 128382 469958 135266 470078
rect 99822 469842 135266 469958
rect 135502 469842 135586 470078
rect 135822 469958 163826 470078
rect 164062 469958 164146 470194
rect 164382 470078 199826 470194
rect 164382 469958 171266 470078
rect 135822 469842 171266 469958
rect 171502 469842 171586 470078
rect 171822 469958 199826 470078
rect 200062 469958 200146 470194
rect 200382 470078 235826 470194
rect 200382 469958 207266 470078
rect 171822 469842 207266 469958
rect 207502 469842 207586 470078
rect 207822 469958 235826 470078
rect 236062 469958 236146 470194
rect 236382 470078 271826 470194
rect 236382 469958 243266 470078
rect 207822 469842 243266 469958
rect 243502 469842 243586 470078
rect 243822 469958 271826 470078
rect 272062 469958 272146 470194
rect 272382 470110 272414 470194
rect 272382 470078 279854 470110
rect 272382 469958 279266 470078
rect 243822 469842 279266 469958
rect 279502 469842 279586 470078
rect 279822 469842 279854 470078
rect 63234 469758 279854 469842
rect 63234 469522 63266 469758
rect 63502 469522 63586 469758
rect 63822 469522 99266 469758
rect 99502 469522 99586 469758
rect 99822 469522 135266 469758
rect 135502 469522 135586 469758
rect 135822 469522 171266 469758
rect 171502 469522 171586 469758
rect 171822 469522 207266 469758
rect 207502 469522 207586 469758
rect 207822 469522 243266 469758
rect 243502 469522 243586 469758
rect 243822 469522 279266 469758
rect 279502 469522 279586 469758
rect 279822 469522 279854 469758
rect 63234 469490 279854 469522
rect 81234 469138 297854 469170
rect 81234 468902 81266 469138
rect 81502 468902 81586 469138
rect 81822 468902 117266 469138
rect 117502 468902 117586 469138
rect 117822 468902 153266 469138
rect 153502 468902 153586 469138
rect 153822 468902 189266 469138
rect 189502 468902 189586 469138
rect 189822 468902 225266 469138
rect 225502 468902 225586 469138
rect 225822 468902 261266 469138
rect 261502 468902 261586 469138
rect 261822 468902 297266 469138
rect 297502 468902 297586 469138
rect 297822 468902 297854 469138
rect 81234 468818 297854 468902
rect 81234 468582 81266 468818
rect 81502 468582 81586 468818
rect 81822 468582 117266 468818
rect 117502 468582 117586 468818
rect 117822 468582 153266 468818
rect 153502 468582 153586 468818
rect 153822 468582 189266 468818
rect 189502 468582 189586 468818
rect 189822 468582 225266 468818
rect 225502 468582 225586 468818
rect 225822 468582 261266 468818
rect 261502 468582 261586 468818
rect 261822 468582 297266 468818
rect 297502 468582 297586 468818
rect 297822 468582 297854 468818
rect 81234 468550 297854 468582
rect 84954 465554 301574 465586
rect 84954 465318 84986 465554
rect 85222 465318 85306 465554
rect 85542 465318 120986 465554
rect 121222 465318 121306 465554
rect 121542 465318 156986 465554
rect 157222 465318 157306 465554
rect 157542 465318 192986 465554
rect 193222 465318 193306 465554
rect 193542 465318 228986 465554
rect 229222 465318 229306 465554
rect 229542 465318 264986 465554
rect 265222 465318 265306 465554
rect 265542 465318 300986 465554
rect 301222 465318 301306 465554
rect 301542 465318 301574 465554
rect 84954 465234 301574 465318
rect 84954 464998 84986 465234
rect 85222 464998 85306 465234
rect 85542 464998 120986 465234
rect 121222 464998 121306 465234
rect 121542 464998 156986 465234
rect 157222 464998 157306 465234
rect 157542 464998 192986 465234
rect 193222 464998 193306 465234
rect 193542 464998 228986 465234
rect 229222 464998 229306 465234
rect 229542 464998 264986 465234
rect 265222 464998 265306 465234
rect 265542 464998 300986 465234
rect 301222 464998 301306 465234
rect 301542 464998 301574 465234
rect 84954 464966 301574 464998
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 380328 453454
rect 380564 453218 516056 453454
rect 516292 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 380328 453134
rect 380564 452898 516056 453134
rect 516292 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 381008 435454
rect 381244 435218 515376 435454
rect 515612 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 381008 435134
rect 381244 434898 515376 435134
rect 515612 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 380328 417454
rect 380564 417218 516056 417454
rect 516292 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 380328 417134
rect 380564 416898 516056 417134
rect 516292 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 61008 399454
rect 61244 399218 195376 399454
rect 195612 399218 221008 399454
rect 221244 399218 355376 399454
rect 355612 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 381008 399454
rect 381244 399218 515376 399454
rect 515612 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 61008 399134
rect 61244 398898 195376 399134
rect 195612 398898 221008 399134
rect 221244 398898 355376 399134
rect 355612 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 381008 399134
rect 381244 398898 515376 399134
rect 515612 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 60328 381454
rect 60564 381218 196056 381454
rect 196292 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 220328 381454
rect 220564 381218 356056 381454
rect 356292 381218 380328 381454
rect 380564 381218 516056 381454
rect 516292 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 60328 381134
rect 60564 380898 196056 381134
rect 196292 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 220328 381134
rect 220564 380898 356056 381134
rect 356292 380898 380328 381134
rect 380564 380898 516056 381134
rect 516292 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect 63234 369954 495854 369986
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 63234 369634 495854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 63234 369366 495854 369398
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect 59514 366234 492134 366266
rect 59514 365998 59546 366234
rect 59782 365998 59866 366234
rect 60102 365998 95546 366234
rect 95782 365998 95866 366234
rect 96102 365998 131546 366234
rect 131782 365998 131866 366234
rect 132102 365998 167546 366234
rect 167782 365998 167866 366234
rect 168102 365998 203546 366234
rect 203782 365998 203866 366234
rect 204102 365998 239546 366234
rect 239782 365998 239866 366234
rect 240102 365998 275546 366234
rect 275782 365998 275866 366234
rect 276102 365998 311546 366234
rect 311782 365998 311866 366234
rect 312102 365998 347546 366234
rect 347782 365998 347866 366234
rect 348102 365998 383546 366234
rect 383782 365998 383866 366234
rect 384102 365998 419546 366234
rect 419782 365998 419866 366234
rect 420102 365998 455546 366234
rect 455782 365998 455866 366234
rect 456102 365998 491546 366234
rect 491782 365998 491866 366234
rect 492102 365998 492134 366234
rect 59514 365914 492134 365998
rect 59514 365678 59546 365914
rect 59782 365678 59866 365914
rect 60102 365678 95546 365914
rect 95782 365678 95866 365914
rect 96102 365678 131546 365914
rect 131782 365678 131866 365914
rect 132102 365678 167546 365914
rect 167782 365678 167866 365914
rect 168102 365678 203546 365914
rect 203782 365678 203866 365914
rect 204102 365678 239546 365914
rect 239782 365678 239866 365914
rect 240102 365678 275546 365914
rect 275782 365678 275866 365914
rect 276102 365678 311546 365914
rect 311782 365678 311866 365914
rect 312102 365678 347546 365914
rect 347782 365678 347866 365914
rect 348102 365678 383546 365914
rect 383782 365678 383866 365914
rect 384102 365678 419546 365914
rect 419782 365678 419866 365914
rect 420102 365678 455546 365914
rect 455782 365678 455866 365914
rect 456102 365678 491546 365914
rect 491782 365678 491866 365914
rect 492102 365678 492134 365914
rect 59514 365646 492134 365678
rect 91794 364394 488414 364426
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 91794 364074 488414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 91794 363806 488414 363838
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect 84954 357554 517574 357586
rect 84954 357318 84986 357554
rect 85222 357318 85306 357554
rect 85542 357318 120986 357554
rect 121222 357318 121306 357554
rect 121542 357318 156986 357554
rect 157222 357318 157306 357554
rect 157542 357318 192986 357554
rect 193222 357318 193306 357554
rect 193542 357318 228986 357554
rect 229222 357318 229306 357554
rect 229542 357318 264986 357554
rect 265222 357318 265306 357554
rect 265542 357318 300986 357554
rect 301222 357318 301306 357554
rect 301542 357318 336986 357554
rect 337222 357318 337306 357554
rect 337542 357318 372986 357554
rect 373222 357318 373306 357554
rect 373542 357318 408986 357554
rect 409222 357318 409306 357554
rect 409542 357318 444986 357554
rect 445222 357318 445306 357554
rect 445542 357318 480986 357554
rect 481222 357318 481306 357554
rect 481542 357318 516986 357554
rect 517222 357318 517306 357554
rect 517542 357318 517574 357554
rect 84954 357234 517574 357318
rect 84954 356998 84986 357234
rect 85222 356998 85306 357234
rect 85542 356998 120986 357234
rect 121222 356998 121306 357234
rect 121542 356998 156986 357234
rect 157222 356998 157306 357234
rect 157542 356998 192986 357234
rect 193222 356998 193306 357234
rect 193542 356998 228986 357234
rect 229222 356998 229306 357234
rect 229542 356998 264986 357234
rect 265222 356998 265306 357234
rect 265542 356998 300986 357234
rect 301222 356998 301306 357234
rect 301542 356998 336986 357234
rect 337222 356998 337306 357234
rect 337542 356998 372986 357234
rect 373222 356998 373306 357234
rect 373542 356998 408986 357234
rect 409222 356998 409306 357234
rect 409542 356998 444986 357234
rect 445222 356998 445306 357234
rect 445542 356998 480986 357234
rect 481222 356998 481306 357234
rect 481542 356998 516986 357234
rect 517222 356998 517306 357234
rect 517542 356998 517574 357234
rect 84954 356966 517574 356998
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 60328 345454
rect 60564 345218 196056 345454
rect 196292 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 220328 345454
rect 220564 345218 356056 345454
rect 356292 345218 380328 345454
rect 380564 345218 516056 345454
rect 516292 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 60328 345134
rect 60564 344898 196056 345134
rect 196292 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 220328 345134
rect 220564 344898 356056 345134
rect 356292 344898 380328 345134
rect 380564 344898 516056 345134
rect 516292 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 61008 327454
rect 61244 327218 195376 327454
rect 195612 327218 221008 327454
rect 221244 327218 355376 327454
rect 355612 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 381008 327454
rect 381244 327218 515376 327454
rect 515612 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 61008 327134
rect 61244 326898 195376 327134
rect 195612 326898 221008 327134
rect 221244 326898 355376 327134
rect 355612 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 381008 327134
rect 381244 326898 515376 327134
rect 515612 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 60328 309454
rect 60564 309218 196056 309454
rect 196292 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 220328 309454
rect 220564 309218 356056 309454
rect 356292 309218 380328 309454
rect 380564 309218 516056 309454
rect 516292 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 60328 309134
rect 60564 308898 196056 309134
rect 196292 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 220328 309134
rect 220564 308898 356056 309134
rect 356292 308898 380328 309134
rect 380564 308898 516056 309134
rect 516292 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 61008 291454
rect 61244 291218 195376 291454
rect 195612 291218 221008 291454
rect 221244 291218 355376 291454
rect 355612 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 381008 291454
rect 381244 291218 515376 291454
rect 515612 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 61008 291134
rect 61244 290898 195376 291134
rect 195612 290898 221008 291134
rect 221244 290898 355376 291134
rect 355612 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 381008 291134
rect 381244 290898 515376 291134
rect 515612 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 60328 273454
rect 60564 273218 196056 273454
rect 196292 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 220328 273454
rect 220564 273218 356056 273454
rect 356292 273218 380328 273454
rect 380564 273218 516056 273454
rect 516292 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 60328 273134
rect 60564 272898 196056 273134
rect 196292 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 220328 273134
rect 220564 272898 356056 273134
rect 356292 272898 380328 273134
rect 380564 272898 516056 273134
rect 516292 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect 66954 265674 499574 265706
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 66954 265354 499574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 66954 265086 499574 265118
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect 63234 261954 495854 261986
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 63234 261634 495854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 63234 261366 495854 261398
rect 59514 260114 492134 260146
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 59514 259794 492134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 59514 259526 492134 259558
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect 91794 256394 488414 256426
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 91794 256074 488414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 91794 255806 488414 255838
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 60328 237454
rect 60564 237218 196056 237454
rect 196292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 220328 237454
rect 220564 237218 356056 237454
rect 356292 237218 380328 237454
rect 380564 237218 516056 237454
rect 516292 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 60328 237134
rect 60564 236898 196056 237134
rect 196292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 220328 237134
rect 220564 236898 356056 237134
rect 356292 236898 380328 237134
rect 380564 236898 516056 237134
rect 516292 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 61008 219454
rect 61244 219218 195376 219454
rect 195612 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 381008 219454
rect 381244 219218 515376 219454
rect 515612 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 61008 219134
rect 61244 218898 195376 219134
rect 195612 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 381008 219134
rect 381244 218898 515376 219134
rect 515612 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 60328 201454
rect 60564 201218 196056 201454
rect 196292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 220328 201454
rect 220564 201218 356056 201454
rect 356292 201218 380328 201454
rect 380564 201218 516056 201454
rect 516292 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 60328 201134
rect 60564 200898 196056 201134
rect 196292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 220328 201134
rect 220564 200898 356056 201134
rect 356292 200898 380328 201134
rect 380564 200898 516056 201134
rect 516292 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 61008 183454
rect 61244 183218 195376 183454
rect 195612 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 381008 183454
rect 381244 183218 515376 183454
rect 515612 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 61008 183134
rect 61244 182898 195376 183134
rect 195612 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 381008 183134
rect 381244 182898 515376 183134
rect 515612 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect 66954 157674 499574 157706
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 66954 157354 499574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 66954 157086 499574 157118
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect 63234 153954 495854 153986
rect 63234 153718 63266 153954
rect 63502 153718 63586 153954
rect 63822 153718 99266 153954
rect 99502 153718 99586 153954
rect 99822 153718 135266 153954
rect 135502 153718 135586 153954
rect 135822 153718 171266 153954
rect 171502 153718 171586 153954
rect 171822 153718 207266 153954
rect 207502 153718 207586 153954
rect 207822 153718 243266 153954
rect 243502 153718 243586 153954
rect 243822 153718 279266 153954
rect 279502 153718 279586 153954
rect 279822 153718 315266 153954
rect 315502 153718 315586 153954
rect 315822 153718 351266 153954
rect 351502 153718 351586 153954
rect 351822 153718 387266 153954
rect 387502 153718 387586 153954
rect 387822 153718 423266 153954
rect 423502 153718 423586 153954
rect 423822 153718 459266 153954
rect 459502 153718 459586 153954
rect 459822 153718 495266 153954
rect 495502 153718 495586 153954
rect 495822 153718 495854 153954
rect 63234 153634 495854 153718
rect 63234 153398 63266 153634
rect 63502 153398 63586 153634
rect 63822 153398 99266 153634
rect 99502 153398 99586 153634
rect 99822 153398 135266 153634
rect 135502 153398 135586 153634
rect 135822 153398 171266 153634
rect 171502 153398 171586 153634
rect 171822 153398 207266 153634
rect 207502 153398 207586 153634
rect 207822 153398 243266 153634
rect 243502 153398 243586 153634
rect 243822 153398 279266 153634
rect 279502 153398 279586 153634
rect 279822 153398 315266 153634
rect 315502 153398 315586 153634
rect 315822 153398 351266 153634
rect 351502 153398 351586 153634
rect 351822 153398 387266 153634
rect 387502 153398 387586 153634
rect 387822 153398 423266 153634
rect 423502 153398 423586 153634
rect 423822 153398 459266 153634
rect 459502 153398 459586 153634
rect 459822 153398 495266 153634
rect 495502 153398 495586 153634
rect 495822 153398 495854 153634
rect 63234 153366 495854 153398
rect 59514 152114 492134 152146
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 59514 151794 492134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 59514 151526 492134 151558
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect 91794 148394 488414 148426
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 91794 148074 488414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 91794 147806 488414 147838
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 60328 129454
rect 60564 129218 196056 129454
rect 196292 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 220328 129454
rect 220564 129218 356056 129454
rect 356292 129218 380328 129454
rect 380564 129218 516056 129454
rect 516292 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 60328 129134
rect 60564 128898 196056 129134
rect 196292 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 220328 129134
rect 220564 128898 356056 129134
rect 356292 128898 380328 129134
rect 380564 128898 516056 129134
rect 516292 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 61008 111454
rect 61244 111218 195376 111454
rect 195612 111218 221008 111454
rect 221244 111218 355376 111454
rect 355612 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 381008 111454
rect 381244 111218 515376 111454
rect 515612 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 61008 111134
rect 61244 110898 195376 111134
rect 195612 110898 221008 111134
rect 221244 110898 355376 111134
rect 355612 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 381008 111134
rect 381244 110898 515376 111134
rect 515612 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 60328 93454
rect 60564 93218 196056 93454
rect 196292 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 220328 93454
rect 220564 93218 356056 93454
rect 356292 93218 380328 93454
rect 380564 93218 516056 93454
rect 516292 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 60328 93134
rect 60564 92898 196056 93134
rect 196292 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 220328 93134
rect 220564 92898 356056 93134
rect 356292 92898 380328 93134
rect 380564 92898 516056 93134
rect 516292 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 61008 75454
rect 61244 75218 195376 75454
rect 195612 75218 221008 75454
rect 221244 75218 355376 75454
rect 355612 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 381008 75454
rect 381244 75218 515376 75454
rect 515612 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 61008 75134
rect 61244 74898 195376 75134
rect 195612 74898 221008 75134
rect 221244 74898 355376 75134
rect 355612 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 381008 75134
rect 381244 74898 515376 75134
rect 515612 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst1
timestamp 0
transform 1 0 60000 0 1 165000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst2
timestamp 0
transform 1 0 60000 0 1 270000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst0
timestamp 0
transform 1 0 380000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst1
timestamp 0
transform 1 0 380000 0 1 165000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst2
timestamp 0
transform 1 0 380000 0 1 270000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst3
timestamp 0
transform 1 0 380000 0 1 375000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 375000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst1
timestamp 0
transform 1 0 220000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst2
timestamp 0
transform 1 0 220000 0 1 165000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst3
timestamp 0
transform 1 0 220000 0 1 270000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst4
timestamp 0
transform 1 0 220000 0 1 375000
box 0 0 136620 83308
use VerySimpleCPU_core  inst_agent_1
timestamp 0
transform 1 0 60000 0 1 560000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_codemaker
timestamp 0
transform 1 0 220000 0 1 560000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_control_tower
timestamp 0
transform 1 0 140000 0 1 560000
box 0 0 60955 63099
use main_controller  inst_main_controller
timestamp 0
transform 1 0 60000 0 1 480000
box 0 0 240000 60000
use main_memory  inst_main_memory
timestamp 0
transform 1 0 320000 0 1 520000
box 0 0 108889 111033
use uart  inst_uart
timestamp 0
transform 1 0 460000 0 1 570000
box 0 0 50000 50000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 145308 74414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 145308 110414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 145308 146414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 145308 182414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 145308 218414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 145308 254414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 145308 290414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 145308 326414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 145308 398414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 145308 434414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 145308 470414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 145308 506414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 250308 74414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 250308 110414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 250308 146414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 250308 182414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 250308 218414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 250308 254414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 250308 290414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 250308 326414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 250308 398414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 250308 434414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 250308 470414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 250308 506414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 355308 74414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 355308 110414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 355308 146414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 355308 182414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 355308 218414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 355308 254414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 355308 290414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 355308 326414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 355308 398414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 355308 434414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 355308 470414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 355308 506414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 460308 74414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 460308 110414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 460308 146414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 460308 182414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 460308 218414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 460308 254414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 460308 290414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 460308 326414 518000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 518000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 460308 398414 518000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 542000 74414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 542000 110414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 542000 146414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 542000 182414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 542000 218414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 542000 254414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 460308 470414 568000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 460308 506414 568000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 625099 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 625099 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 625099 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 625099 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 625099 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 625099 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 542000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 633033 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 633033 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 633033 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 460308 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 622000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 622000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 145308 78134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 145308 114134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 145308 150134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 145308 186134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 145308 222134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 145308 258134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 145308 294134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 145308 330134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 145308 402134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 145308 438134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 145308 474134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 145308 510134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 250308 78134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 250308 114134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 250308 150134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 250308 186134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 250308 222134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 250308 258134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 250308 294134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 250308 330134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 250308 402134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 250308 438134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 250308 474134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 250308 510134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 355308 78134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 355308 114134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 355308 150134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 355308 186134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 355308 222134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 355308 258134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 355308 294134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 355308 330134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 355308 402134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 355308 438134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 355308 474134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 355308 510134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 460308 78134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 460308 114134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 460308 150134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 460308 186134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 460308 222134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 460308 258134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 460308 294134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 460308 330134 518000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 518000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 460308 402134 518000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 542000 78134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 542000 114134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 542000 150134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 542000 186134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 542000 222134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 542000 258134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 460308 474134 568000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 460308 510134 568000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 625099 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 625099 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 625099 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 625099 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 625099 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 625099 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 542000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 633033 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 633033 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 633033 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 460308 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 622000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 622000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s 81234 468550 297854 469170 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 145308 81854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 145308 117854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 145308 153854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 145308 189854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 145308 225854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 145308 261854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 145308 297854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 145308 333854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 145308 405854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 145308 441854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 145308 477854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 145308 513854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 250308 81854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 250308 117854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 250308 153854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 250308 189854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 250308 225854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 250308 261854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 250308 297854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 250308 333854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 250308 405854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 250308 441854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 250308 477854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 250308 513854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 355308 81854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 355308 117854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 355308 153854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 355308 189854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 355308 225854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 355308 261854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 355308 297854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 355308 333854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 355308 405854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 355308 441854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 355308 477854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 355308 513854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 460308 81854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 460308 117854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 460308 153854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 460308 189854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 460308 225854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 460308 261854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 460308 297854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 460308 333854 518000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 518000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 460308 405854 518000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 542000 81854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 542000 117854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 542000 153854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 542000 189854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 542000 225854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 542000 261854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 460308 477854 568000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 625099 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 625099 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 625099 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 625099 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 625099 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 625099 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 542000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 633033 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 633033 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 633033 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 460308 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 622000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 460308 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s 84954 356966 517574 357586 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s 84954 464966 301574 465586 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 145308 85574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 145308 121574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 145308 157574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 145308 193574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 145308 229574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 145308 265574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 145308 301574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 145308 337574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 145308 409574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 145308 445574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 145308 481574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 145308 517574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 250308 85574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 250308 121574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 250308 157574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 250308 193574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 250308 229574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 250308 265574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 250308 301574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 250308 337574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 250308 409574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 250308 445574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 250308 481574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 250308 517574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 355308 85574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 355308 121574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 355308 157574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 355308 193574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 355308 229574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 355308 265574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 355308 301574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 355308 337574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 355308 409574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 355308 445574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 355308 481574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 355308 517574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 460308 85574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 460308 121574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 460308 157574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 460308 193574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 460308 229574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 460308 265574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 460308 301574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 460308 337574 518000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 518000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 460308 409574 518000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 542000 85574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 542000 121574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 542000 157574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 542000 193574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 542000 229574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 542000 265574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 460308 481574 568000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 625099 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 625099 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 625099 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 625099 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 625099 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 625099 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 542000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 633033 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 633033 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 633033 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 460308 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 622000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 460308 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 153366 495854 153986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 261366 495854 261986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 369366 495854 369986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 469490 279854 470110 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 549366 279854 549986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 145308 63854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 145308 99854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 145308 135854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 145308 171854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 145308 243854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 145308 279854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 145308 315854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 145308 351854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 145308 387854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 145308 423854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 145308 459854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 145308 495854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 250308 63854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 250308 99854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 250308 135854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 250308 171854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 250308 243854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 250308 279854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 250308 315854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 250308 351854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 250308 387854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 250308 423854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 250308 459854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 250308 495854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 355308 63854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 355308 99854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 355308 135854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 355308 171854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 355308 243854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 355308 279854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 355308 315854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 355308 351854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 355308 387854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 355308 423854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 355308 459854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 355308 495854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 460308 63854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 460308 99854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 460308 135854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 460308 171854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 460308 243854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 460308 279854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 460308 351854 518000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 460308 387854 518000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 460308 423854 518000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 542000 63854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 542000 99854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 542000 171854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 542000 243854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 542000 279854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 460308 459854 568000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 460308 495854 568000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 625099 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 625099 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 542000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 625099 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 542000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 625099 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 625099 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 460308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 633033 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 633033 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 633033 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 622000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 622000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 157086 499574 157706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 265086 499574 265706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 553086 283574 553706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 145308 67574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 145308 103574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 145308 139574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 145308 175574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 145308 247574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 145308 283574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 145308 319574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 145308 355574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 145308 391574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 145308 427574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 145308 463574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 145308 499574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 250308 67574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 250308 103574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 250308 139574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 250308 175574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 250308 247574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 250308 283574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 250308 319574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 250308 355574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 250308 391574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 250308 427574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 250308 463574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 250308 499574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 355308 67574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 355308 103574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 355308 139574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 355308 175574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 355308 247574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 355308 283574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 355308 319574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 355308 355574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 355308 391574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 355308 427574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 355308 463574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 355308 499574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 460308 67574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 460308 103574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 460308 139574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 460308 175574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 460308 247574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 460308 283574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 460308 319574 518000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 460308 355574 518000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 460308 391574 518000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 460308 427574 518000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 542000 67574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 542000 103574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 542000 139574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 542000 175574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 542000 247574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 542000 283574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 460308 463574 568000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 460308 499574 568000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 625099 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 625099 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 625099 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 625099 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 542000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 625099 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 625099 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 633033 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 633033 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 633033 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 633033 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 622000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 622000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 147806 488414 148426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 255806 488414 256426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 363806 488414 364426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 469926 272414 470546 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 543806 272414 544426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 145308 92414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 145308 128414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 145308 164414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 145308 236414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 145308 272414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 145308 308414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 145308 344414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 145308 380414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 145308 416414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 145308 452414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 145308 488414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 250308 92414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 250308 128414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 250308 164414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 250308 236414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 250308 272414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 250308 308414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 250308 344414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 250308 380414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 250308 416414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 250308 452414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 250308 488414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 355308 92414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 355308 128414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 355308 164414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 355308 236414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 355308 272414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 355308 308414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 355308 344414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 355308 380414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 355308 416414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 355308 452414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 355308 488414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 460308 92414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 460308 128414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 460308 164414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 460308 236414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 460308 272414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 460308 344414 518000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 460308 380414 518000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 460308 416414 518000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 542000 92414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 542000 164414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 542000 200414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 542000 236414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 542000 272414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 460308 488414 568000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 625099 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 542000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 625099 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 625099 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 625099 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 625099 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 460308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 633033 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 633033 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 633033 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 460308 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 622000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 151526 492134 152146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 259526 492134 260146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 365646 492134 366266 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 473646 276134 474266 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 547526 276134 548146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 145308 60134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 145308 96134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 145308 132134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 145308 168134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 145308 240134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 145308 276134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 145308 312134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 145308 348134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 145308 384134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 145308 420134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 145308 456134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 145308 492134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 250308 60134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 250308 96134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 250308 132134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 250308 168134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 250308 240134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 250308 276134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 250308 312134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 250308 348134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 250308 384134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 250308 420134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 250308 456134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 250308 492134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 355308 60134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 355308 96134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 355308 132134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 355308 168134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 355308 240134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 355308 276134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 355308 312134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 355308 348134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 355308 384134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 355308 420134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 355308 456134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 355308 492134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 460308 60134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 460308 96134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 460308 132134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 460308 168134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 460308 240134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 460308 276134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 460308 348134 518000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 460308 384134 518000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 460308 420134 518000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 542000 60134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 542000 96134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 542000 168134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 542000 240134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 542000 276134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 460308 492134 568000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 625099 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 625099 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 542000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 625099 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 542000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 625099 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 625099 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 460308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 633033 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 633033 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 633033 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 460308 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 622000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
