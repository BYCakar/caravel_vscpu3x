magic
tech sky130A
magscale 1 2
timestamp 1655556856
<< obsli1 >>
rect 61104 279159 509800 424401
<< obsm1 >>
rect 566 3408 580414 700392
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 580410 703610
rect 572 536 580410 703464
rect 710 480 1590 536
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6374 536
rect 6598 480 7570 536
rect 7794 480 8674 536
rect 8898 480 9870 536
rect 10094 480 11066 536
rect 11290 480 12262 536
rect 12486 480 13458 536
rect 13682 480 14654 536
rect 14878 480 15850 536
rect 16074 480 16954 536
rect 17178 480 18150 536
rect 18374 480 19346 536
rect 19570 480 20542 536
rect 20766 480 21738 536
rect 21962 480 22934 536
rect 23158 480 24130 536
rect 24354 480 25234 536
rect 25458 480 26430 536
rect 26654 480 27626 536
rect 27850 480 28822 536
rect 29046 480 30018 536
rect 30242 480 31214 536
rect 31438 480 32318 536
rect 32542 480 33514 536
rect 33738 480 34710 536
rect 34934 480 35906 536
rect 36130 480 37102 536
rect 37326 480 38298 536
rect 38522 480 39494 536
rect 39718 480 40598 536
rect 40822 480 41794 536
rect 42018 480 42990 536
rect 43214 480 44186 536
rect 44410 480 45382 536
rect 45606 480 46578 536
rect 46802 480 47774 536
rect 47998 480 48878 536
rect 49102 480 50074 536
rect 50298 480 51270 536
rect 51494 480 52466 536
rect 52690 480 53662 536
rect 53886 480 54858 536
rect 55082 480 55962 536
rect 56186 480 57158 536
rect 57382 480 58354 536
rect 58578 480 59550 536
rect 59774 480 60746 536
rect 60970 480 61942 536
rect 62166 480 63138 536
rect 63362 480 64242 536
rect 64466 480 65438 536
rect 65662 480 66634 536
rect 66858 480 67830 536
rect 68054 480 69026 536
rect 69250 480 70222 536
rect 70446 480 71418 536
rect 71642 480 72522 536
rect 72746 480 73718 536
rect 73942 480 74914 536
rect 75138 480 76110 536
rect 76334 480 77306 536
rect 77530 480 78502 536
rect 78726 480 79606 536
rect 79830 480 80802 536
rect 81026 480 81998 536
rect 82222 480 83194 536
rect 83418 480 84390 536
rect 84614 480 85586 536
rect 85810 480 86782 536
rect 87006 480 87886 536
rect 88110 480 89082 536
rect 89306 480 90278 536
rect 90502 480 91474 536
rect 91698 480 92670 536
rect 92894 480 93866 536
rect 94090 480 95062 536
rect 95286 480 96166 536
rect 96390 480 97362 536
rect 97586 480 98558 536
rect 98782 480 99754 536
rect 99978 480 100950 536
rect 101174 480 102146 536
rect 102370 480 103250 536
rect 103474 480 104446 536
rect 104670 480 105642 536
rect 105866 480 106838 536
rect 107062 480 108034 536
rect 108258 480 109230 536
rect 109454 480 110426 536
rect 110650 480 111530 536
rect 111754 480 112726 536
rect 112950 480 113922 536
rect 114146 480 115118 536
rect 115342 480 116314 536
rect 116538 480 117510 536
rect 117734 480 118706 536
rect 118930 480 119810 536
rect 120034 480 121006 536
rect 121230 480 122202 536
rect 122426 480 123398 536
rect 123622 480 124594 536
rect 124818 480 125790 536
rect 126014 480 126894 536
rect 127118 480 128090 536
rect 128314 480 129286 536
rect 129510 480 130482 536
rect 130706 480 131678 536
rect 131902 480 132874 536
rect 133098 480 134070 536
rect 134294 480 135174 536
rect 135398 480 136370 536
rect 136594 480 137566 536
rect 137790 480 138762 536
rect 138986 480 139958 536
rect 140182 480 141154 536
rect 141378 480 142350 536
rect 142574 480 143454 536
rect 143678 480 144650 536
rect 144874 480 145846 536
rect 146070 480 147042 536
rect 147266 480 148238 536
rect 148462 480 149434 536
rect 149658 480 150538 536
rect 150762 480 151734 536
rect 151958 480 152930 536
rect 153154 480 154126 536
rect 154350 480 155322 536
rect 155546 480 156518 536
rect 156742 480 157714 536
rect 157938 480 158818 536
rect 159042 480 160014 536
rect 160238 480 161210 536
rect 161434 480 162406 536
rect 162630 480 163602 536
rect 163826 480 164798 536
rect 165022 480 165994 536
rect 166218 480 167098 536
rect 167322 480 168294 536
rect 168518 480 169490 536
rect 169714 480 170686 536
rect 170910 480 171882 536
rect 172106 480 173078 536
rect 173302 480 174182 536
rect 174406 480 175378 536
rect 175602 480 176574 536
rect 176798 480 177770 536
rect 177994 480 178966 536
rect 179190 480 180162 536
rect 180386 480 181358 536
rect 181582 480 182462 536
rect 182686 480 183658 536
rect 183882 480 184854 536
rect 185078 480 186050 536
rect 186274 480 187246 536
rect 187470 480 188442 536
rect 188666 480 189638 536
rect 189862 480 190742 536
rect 190966 480 191938 536
rect 192162 480 193134 536
rect 193358 480 194330 536
rect 194554 480 195526 536
rect 195750 480 196722 536
rect 196946 480 197826 536
rect 198050 480 199022 536
rect 199246 480 200218 536
rect 200442 480 201414 536
rect 201638 480 202610 536
rect 202834 480 203806 536
rect 204030 480 205002 536
rect 205226 480 206106 536
rect 206330 480 207302 536
rect 207526 480 208498 536
rect 208722 480 209694 536
rect 209918 480 210890 536
rect 211114 480 212086 536
rect 212310 480 213282 536
rect 213506 480 214386 536
rect 214610 480 215582 536
rect 215806 480 216778 536
rect 217002 480 217974 536
rect 218198 480 219170 536
rect 219394 480 220366 536
rect 220590 480 221470 536
rect 221694 480 222666 536
rect 222890 480 223862 536
rect 224086 480 225058 536
rect 225282 480 226254 536
rect 226478 480 227450 536
rect 227674 480 228646 536
rect 228870 480 229750 536
rect 229974 480 230946 536
rect 231170 480 232142 536
rect 232366 480 233338 536
rect 233562 480 234534 536
rect 234758 480 235730 536
rect 235954 480 236926 536
rect 237150 480 238030 536
rect 238254 480 239226 536
rect 239450 480 240422 536
rect 240646 480 241618 536
rect 241842 480 242814 536
rect 243038 480 244010 536
rect 244234 480 245114 536
rect 245338 480 246310 536
rect 246534 480 247506 536
rect 247730 480 248702 536
rect 248926 480 249898 536
rect 250122 480 251094 536
rect 251318 480 252290 536
rect 252514 480 253394 536
rect 253618 480 254590 536
rect 254814 480 255786 536
rect 256010 480 256982 536
rect 257206 480 258178 536
rect 258402 480 259374 536
rect 259598 480 260570 536
rect 260794 480 261674 536
rect 261898 480 262870 536
rect 263094 480 264066 536
rect 264290 480 265262 536
rect 265486 480 266458 536
rect 266682 480 267654 536
rect 267878 480 268758 536
rect 268982 480 269954 536
rect 270178 480 271150 536
rect 271374 480 272346 536
rect 272570 480 273542 536
rect 273766 480 274738 536
rect 274962 480 275934 536
rect 276158 480 277038 536
rect 277262 480 278234 536
rect 278458 480 279430 536
rect 279654 480 280626 536
rect 280850 480 281822 536
rect 282046 480 283018 536
rect 283242 480 284214 536
rect 284438 480 285318 536
rect 285542 480 286514 536
rect 286738 480 287710 536
rect 287934 480 288906 536
rect 289130 480 290102 536
rect 290326 480 291298 536
rect 291522 480 292494 536
rect 292718 480 293598 536
rect 293822 480 294794 536
rect 295018 480 295990 536
rect 296214 480 297186 536
rect 297410 480 298382 536
rect 298606 480 299578 536
rect 299802 480 300682 536
rect 300906 480 301878 536
rect 302102 480 303074 536
rect 303298 480 304270 536
rect 304494 480 305466 536
rect 305690 480 306662 536
rect 306886 480 307858 536
rect 308082 480 308962 536
rect 309186 480 310158 536
rect 310382 480 311354 536
rect 311578 480 312550 536
rect 312774 480 313746 536
rect 313970 480 314942 536
rect 315166 480 316138 536
rect 316362 480 317242 536
rect 317466 480 318438 536
rect 318662 480 319634 536
rect 319858 480 320830 536
rect 321054 480 322026 536
rect 322250 480 323222 536
rect 323446 480 324326 536
rect 324550 480 325522 536
rect 325746 480 326718 536
rect 326942 480 327914 536
rect 328138 480 329110 536
rect 329334 480 330306 536
rect 330530 480 331502 536
rect 331726 480 332606 536
rect 332830 480 333802 536
rect 334026 480 334998 536
rect 335222 480 336194 536
rect 336418 480 337390 536
rect 337614 480 338586 536
rect 338810 480 339782 536
rect 340006 480 340886 536
rect 341110 480 342082 536
rect 342306 480 343278 536
rect 343502 480 344474 536
rect 344698 480 345670 536
rect 345894 480 346866 536
rect 347090 480 347970 536
rect 348194 480 349166 536
rect 349390 480 350362 536
rect 350586 480 351558 536
rect 351782 480 352754 536
rect 352978 480 353950 536
rect 354174 480 355146 536
rect 355370 480 356250 536
rect 356474 480 357446 536
rect 357670 480 358642 536
rect 358866 480 359838 536
rect 360062 480 361034 536
rect 361258 480 362230 536
rect 362454 480 363426 536
rect 363650 480 364530 536
rect 364754 480 365726 536
rect 365950 480 366922 536
rect 367146 480 368118 536
rect 368342 480 369314 536
rect 369538 480 370510 536
rect 370734 480 371614 536
rect 371838 480 372810 536
rect 373034 480 374006 536
rect 374230 480 375202 536
rect 375426 480 376398 536
rect 376622 480 377594 536
rect 377818 480 378790 536
rect 379014 480 379894 536
rect 380118 480 381090 536
rect 381314 480 382286 536
rect 382510 480 383482 536
rect 383706 480 384678 536
rect 384902 480 385874 536
rect 386098 480 387070 536
rect 387294 480 388174 536
rect 388398 480 389370 536
rect 389594 480 390566 536
rect 390790 480 391762 536
rect 391986 480 392958 536
rect 393182 480 394154 536
rect 394378 480 395258 536
rect 395482 480 396454 536
rect 396678 480 397650 536
rect 397874 480 398846 536
rect 399070 480 400042 536
rect 400266 480 401238 536
rect 401462 480 402434 536
rect 402658 480 403538 536
rect 403762 480 404734 536
rect 404958 480 405930 536
rect 406154 480 407126 536
rect 407350 480 408322 536
rect 408546 480 409518 536
rect 409742 480 410714 536
rect 410938 480 411818 536
rect 412042 480 413014 536
rect 413238 480 414210 536
rect 414434 480 415406 536
rect 415630 480 416602 536
rect 416826 480 417798 536
rect 418022 480 418902 536
rect 419126 480 420098 536
rect 420322 480 421294 536
rect 421518 480 422490 536
rect 422714 480 423686 536
rect 423910 480 424882 536
rect 425106 480 426078 536
rect 426302 480 427182 536
rect 427406 480 428378 536
rect 428602 480 429574 536
rect 429798 480 430770 536
rect 430994 480 431966 536
rect 432190 480 433162 536
rect 433386 480 434358 536
rect 434582 480 435462 536
rect 435686 480 436658 536
rect 436882 480 437854 536
rect 438078 480 439050 536
rect 439274 480 440246 536
rect 440470 480 441442 536
rect 441666 480 442546 536
rect 442770 480 443742 536
rect 443966 480 444938 536
rect 445162 480 446134 536
rect 446358 480 447330 536
rect 447554 480 448526 536
rect 448750 480 449722 536
rect 449946 480 450826 536
rect 451050 480 452022 536
rect 452246 480 453218 536
rect 453442 480 454414 536
rect 454638 480 455610 536
rect 455834 480 456806 536
rect 457030 480 458002 536
rect 458226 480 459106 536
rect 459330 480 460302 536
rect 460526 480 461498 536
rect 461722 480 462694 536
rect 462918 480 463890 536
rect 464114 480 465086 536
rect 465310 480 466190 536
rect 466414 480 467386 536
rect 467610 480 468582 536
rect 468806 480 469778 536
rect 470002 480 470974 536
rect 471198 480 472170 536
rect 472394 480 473366 536
rect 473590 480 474470 536
rect 474694 480 475666 536
rect 475890 480 476862 536
rect 477086 480 478058 536
rect 478282 480 479254 536
rect 479478 480 480450 536
rect 480674 480 481646 536
rect 481870 480 482750 536
rect 482974 480 483946 536
rect 484170 480 485142 536
rect 485366 480 486338 536
rect 486562 480 487534 536
rect 487758 480 488730 536
rect 488954 480 489834 536
rect 490058 480 491030 536
rect 491254 480 492226 536
rect 492450 480 493422 536
rect 493646 480 494618 536
rect 494842 480 495814 536
rect 496038 480 497010 536
rect 497234 480 498114 536
rect 498338 480 499310 536
rect 499534 480 500506 536
rect 500730 480 501702 536
rect 501926 480 502898 536
rect 503122 480 504094 536
rect 504318 480 505290 536
rect 505514 480 506394 536
rect 506618 480 507590 536
rect 507814 480 508786 536
rect 509010 480 509982 536
rect 510206 480 511178 536
rect 511402 480 512374 536
rect 512598 480 513478 536
rect 513702 480 514674 536
rect 514898 480 515870 536
rect 516094 480 517066 536
rect 517290 480 518262 536
rect 518486 480 519458 536
rect 519682 480 520654 536
rect 520878 480 521758 536
rect 521982 480 522954 536
rect 523178 480 524150 536
rect 524374 480 525346 536
rect 525570 480 526542 536
rect 526766 480 527738 536
rect 527962 480 528934 536
rect 529158 480 530038 536
rect 530262 480 531234 536
rect 531458 480 532430 536
rect 532654 480 533626 536
rect 533850 480 534822 536
rect 535046 480 536018 536
rect 536242 480 537122 536
rect 537346 480 538318 536
rect 538542 480 539514 536
rect 539738 480 540710 536
rect 540934 480 541906 536
rect 542130 480 543102 536
rect 543326 480 544298 536
rect 544522 480 545402 536
rect 545626 480 546598 536
rect 546822 480 547794 536
rect 548018 480 548990 536
rect 549214 480 550186 536
rect 550410 480 551382 536
rect 551606 480 552578 536
rect 552802 480 553682 536
rect 553906 480 554878 536
rect 555102 480 556074 536
rect 556298 480 557270 536
rect 557494 480 558466 536
rect 558690 480 559662 536
rect 559886 480 560766 536
rect 560990 480 561962 536
rect 562186 480 563158 536
rect 563382 480 564354 536
rect 564578 480 565550 536
rect 565774 480 566746 536
rect 566970 480 567942 536
rect 568166 480 569046 536
rect 569270 480 570242 536
rect 570466 480 571438 536
rect 571662 480 572634 536
rect 572858 480 573830 536
rect 574054 480 575026 536
rect 575250 480 576222 536
rect 576446 480 577326 536
rect 577550 480 578522 536
rect 578746 480 579718 536
rect 579942 480 580410 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 480 697540 583586 700365
rect 560 697404 583586 697540
rect 560 697140 583440 697404
rect 480 697004 583440 697140
rect 480 684484 583586 697004
rect 560 684084 583586 684484
rect 480 684076 583586 684084
rect 480 683676 583440 684076
rect 480 671428 583586 683676
rect 560 671028 583586 671428
rect 480 670884 583586 671028
rect 480 670484 583440 670884
rect 480 658372 583586 670484
rect 560 657972 583586 658372
rect 480 657556 583586 657972
rect 480 657156 583440 657556
rect 480 645316 583586 657156
rect 560 644916 583586 645316
rect 480 644228 583586 644916
rect 480 643828 583440 644228
rect 480 632260 583586 643828
rect 560 631860 583586 632260
rect 480 631036 583586 631860
rect 480 630636 583440 631036
rect 480 619340 583586 630636
rect 560 618940 583586 619340
rect 480 617708 583586 618940
rect 480 617308 583440 617708
rect 480 606284 583586 617308
rect 560 605884 583586 606284
rect 480 604380 583586 605884
rect 480 603980 583440 604380
rect 480 593228 583586 603980
rect 560 592828 583586 593228
rect 480 591188 583586 592828
rect 480 590788 583440 591188
rect 480 580172 583586 590788
rect 560 579772 583586 580172
rect 480 577860 583586 579772
rect 480 577460 583440 577860
rect 480 567116 583586 577460
rect 560 566716 583586 567116
rect 480 564532 583586 566716
rect 480 564132 583440 564532
rect 480 554060 583586 564132
rect 560 553660 583586 554060
rect 480 551340 583586 553660
rect 480 550940 583440 551340
rect 480 541004 583586 550940
rect 560 540604 583586 541004
rect 480 538012 583586 540604
rect 480 537612 583440 538012
rect 480 528084 583586 537612
rect 560 527684 583586 528084
rect 480 524684 583586 527684
rect 480 524284 583440 524684
rect 480 515028 583586 524284
rect 560 514628 583586 515028
rect 480 511492 583586 514628
rect 480 511092 583440 511492
rect 480 501972 583586 511092
rect 560 501572 583586 501972
rect 480 498164 583586 501572
rect 480 497764 583440 498164
rect 480 488916 583586 497764
rect 560 488516 583586 488916
rect 480 484836 583586 488516
rect 480 484436 583440 484836
rect 480 475860 583586 484436
rect 560 475460 583586 475860
rect 480 471644 583586 475460
rect 480 471244 583440 471644
rect 480 462804 583586 471244
rect 560 462404 583586 462804
rect 480 458316 583586 462404
rect 480 457916 583440 458316
rect 480 449748 583586 457916
rect 560 449348 583586 449748
rect 480 444988 583586 449348
rect 480 444588 583440 444988
rect 480 436828 583586 444588
rect 560 436428 583586 436828
rect 480 431796 583586 436428
rect 480 431396 583440 431796
rect 480 423772 583586 431396
rect 560 423372 583586 423772
rect 480 418468 583586 423372
rect 480 418068 583440 418468
rect 480 410716 583586 418068
rect 560 410316 583586 410716
rect 480 405140 583586 410316
rect 480 404740 583440 405140
rect 480 397660 583586 404740
rect 560 397260 583586 397660
rect 480 391948 583586 397260
rect 480 391548 583440 391948
rect 480 384604 583586 391548
rect 560 384204 583586 384604
rect 480 378620 583586 384204
rect 480 378220 583440 378620
rect 480 371548 583586 378220
rect 560 371148 583586 371548
rect 480 365292 583586 371148
rect 480 364892 583440 365292
rect 480 358628 583586 364892
rect 560 358228 583586 358628
rect 480 352100 583586 358228
rect 480 351700 583440 352100
rect 480 345572 583586 351700
rect 560 345172 583586 345572
rect 480 338772 583586 345172
rect 480 338372 583440 338772
rect 480 332516 583586 338372
rect 560 332116 583586 332516
rect 480 325444 583586 332116
rect 480 325044 583440 325444
rect 480 319460 583586 325044
rect 560 319060 583586 319460
rect 480 312252 583586 319060
rect 480 311852 583440 312252
rect 480 306404 583586 311852
rect 560 306004 583586 306404
rect 480 298924 583586 306004
rect 480 298524 583440 298924
rect 480 293348 583586 298524
rect 560 292948 583586 293348
rect 480 285596 583586 292948
rect 480 285196 583440 285596
rect 480 280292 583586 285196
rect 560 279892 583586 280292
rect 480 272404 583586 279892
rect 480 272004 583440 272404
rect 480 267372 583586 272004
rect 560 266972 583586 267372
rect 480 259076 583586 266972
rect 480 258676 583440 259076
rect 480 254316 583586 258676
rect 560 253916 583586 254316
rect 480 245748 583586 253916
rect 480 245348 583440 245748
rect 480 241260 583586 245348
rect 560 240860 583586 241260
rect 480 232556 583586 240860
rect 480 232156 583440 232556
rect 480 228204 583586 232156
rect 560 227804 583586 228204
rect 480 219228 583586 227804
rect 480 218828 583440 219228
rect 480 215148 583586 218828
rect 560 214748 583586 215148
rect 480 205900 583586 214748
rect 480 205500 583440 205900
rect 480 202092 583586 205500
rect 560 201692 583586 202092
rect 480 192708 583586 201692
rect 480 192308 583440 192708
rect 480 189036 583586 192308
rect 560 188636 583586 189036
rect 480 179380 583586 188636
rect 480 178980 583440 179380
rect 480 176116 583586 178980
rect 560 175716 583586 176116
rect 480 166052 583586 175716
rect 480 165652 583440 166052
rect 480 163060 583586 165652
rect 560 162660 583586 163060
rect 480 152860 583586 162660
rect 480 152460 583440 152860
rect 480 150004 583586 152460
rect 560 149604 583586 150004
rect 480 139532 583586 149604
rect 480 139132 583440 139532
rect 480 136948 583586 139132
rect 560 136548 583586 136948
rect 480 126204 583586 136548
rect 480 125804 583440 126204
rect 480 123892 583586 125804
rect 560 123492 583586 123892
rect 480 113012 583586 123492
rect 480 112612 583440 113012
rect 480 110836 583586 112612
rect 560 110436 583586 110836
rect 480 99684 583586 110436
rect 480 99284 583440 99684
rect 480 97780 583586 99284
rect 560 97380 583586 97780
rect 480 86356 583586 97380
rect 480 85956 583440 86356
rect 480 84860 583586 85956
rect 560 84460 583586 84860
rect 480 73164 583586 84460
rect 480 72764 583440 73164
rect 480 71804 583586 72764
rect 560 71404 583586 71804
rect 480 59836 583586 71404
rect 480 59436 583440 59836
rect 480 58748 583586 59436
rect 560 58348 583586 58748
rect 480 46508 583586 58348
rect 480 46108 583440 46508
rect 480 45692 583586 46108
rect 560 45292 583586 45692
rect 480 33316 583586 45292
rect 480 32916 583440 33316
rect 480 32636 583586 32916
rect 560 32236 583586 32636
rect 480 19988 583586 32236
rect 480 19588 583440 19988
rect 480 19580 583586 19588
rect 560 19180 583586 19580
rect 480 11595 583586 19180
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 -5734 9854 709670
rect 12954 -7654 13574 711590
rect 15794 -1894 16414 705830
rect 19514 -3814 20134 707750
rect 23234 -5734 23854 709670
rect 26954 -7654 27574 711590
rect 29794 -1894 30414 705830
rect 33514 -3814 34134 707750
rect 37234 -5734 37854 709670
rect 40954 -7654 41574 711590
rect 43794 -1894 44414 705830
rect 47514 -3814 48134 707750
rect 51234 -5734 51854 709670
rect 54954 -7654 55574 711590
rect 57794 645308 58414 705830
rect 61514 645308 62134 707750
rect 65234 645308 65854 709670
rect 68954 645308 69574 711590
rect 71794 645308 72414 705830
rect 75514 645308 76134 707750
rect 79234 645308 79854 709670
rect 82954 645308 83574 711590
rect 85794 645308 86414 705830
rect 89514 645308 90134 707750
rect 93234 645308 93854 709670
rect 96954 645308 97574 711590
rect 99794 645308 100414 705830
rect 103514 645308 104134 707750
rect 107234 645308 107854 709670
rect 110954 645308 111574 711590
rect 113794 645308 114414 705830
rect 117514 645308 118134 707750
rect 121234 645308 121854 709670
rect 124954 645308 125574 711590
rect 127794 645308 128414 705830
rect 131514 645308 132134 707750
rect 135234 645308 135854 709670
rect 138954 645308 139574 711590
rect 141794 645308 142414 705830
rect 145514 645308 146134 707750
rect 149234 645308 149854 709670
rect 152954 645308 153574 711590
rect 155794 645308 156414 705830
rect 159514 645308 160134 707750
rect 163234 645308 163854 709670
rect 166954 645308 167574 711590
rect 169794 645308 170414 705830
rect 173514 645308 174134 707750
rect 177234 645308 177854 709670
rect 180954 645308 181574 711590
rect 183794 645308 184414 705830
rect 187514 645308 188134 707750
rect 191234 645308 191854 709670
rect 194954 645308 195574 711590
rect 197794 645308 198414 705830
rect 57794 538308 58414 558000
rect 61514 538308 62134 558000
rect 65234 538308 65854 558000
rect 68954 538308 69574 558000
rect 71794 538308 72414 558000
rect 75514 538308 76134 558000
rect 79234 538308 79854 558000
rect 82954 538308 83574 558000
rect 85794 538308 86414 558000
rect 89514 538308 90134 558000
rect 93234 538308 93854 558000
rect 96954 538308 97574 558000
rect 99794 538308 100414 558000
rect 103514 538308 104134 558000
rect 107234 538308 107854 558000
rect 110954 538308 111574 558000
rect 113794 538308 114414 558000
rect 117514 538308 118134 558000
rect 121234 538308 121854 558000
rect 124954 538308 125574 558000
rect 127794 538308 128414 558000
rect 131514 538308 132134 558000
rect 135234 538308 135854 558000
rect 138954 538308 139574 558000
rect 141794 538308 142414 558000
rect 145514 538308 146134 558000
rect 149234 538308 149854 558000
rect 152954 538308 153574 558000
rect 155794 538308 156414 558000
rect 159514 538308 160134 558000
rect 163234 538308 163854 558000
rect 166954 538308 167574 558000
rect 169794 538308 170414 558000
rect 173514 538308 174134 558000
rect 177234 538308 177854 558000
rect 180954 538308 181574 558000
rect 183794 538308 184414 558000
rect 187514 538308 188134 558000
rect 191234 538308 191854 558000
rect 194954 538308 195574 558000
rect 197794 538308 198414 558000
rect 57794 427033 58414 451000
rect 61514 427033 62134 451000
rect 65234 427033 65854 451000
rect 68954 427033 69574 451000
rect 71794 427033 72414 451000
rect 75514 427033 76134 451000
rect 79234 427033 79854 451000
rect 82954 427033 83574 451000
rect 85794 427033 86414 451000
rect 89514 427033 90134 451000
rect 93234 427033 93854 451000
rect 96954 427033 97574 451000
rect 99794 427033 100414 451000
rect 103514 427033 104134 451000
rect 107234 427033 107854 451000
rect 110954 427033 111574 451000
rect 113794 427033 114414 451000
rect 117514 427033 118134 451000
rect 121234 427033 121854 451000
rect 124954 427033 125574 451000
rect 127794 427033 128414 451000
rect 131514 427033 132134 451000
rect 135234 427033 135854 451000
rect 138954 427033 139574 451000
rect 141794 427033 142414 451000
rect 145514 427033 146134 451000
rect 149234 427033 149854 451000
rect 152954 427033 153574 451000
rect 155794 427033 156414 451000
rect 159514 427033 160134 451000
rect 163234 427033 163854 451000
rect 166954 427033 167574 451000
rect 169794 427033 170414 451000
rect 57794 252308 58414 312000
rect 61514 252308 62134 312000
rect 65234 252308 65854 312000
rect 68954 252308 69574 312000
rect 71794 252308 72414 312000
rect 75514 252308 76134 312000
rect 79234 252308 79854 312000
rect 82954 252308 83574 312000
rect 85794 252308 86414 312000
rect 89514 252308 90134 312000
rect 93234 252308 93854 312000
rect 96954 252308 97574 312000
rect 99794 252308 100414 312000
rect 103514 252308 104134 312000
rect 107234 252308 107854 312000
rect 110954 252308 111574 312000
rect 113794 252308 114414 312000
rect 117514 252308 118134 312000
rect 121234 252308 121854 312000
rect 124954 252308 125574 312000
rect 127794 252308 128414 312000
rect 131514 252308 132134 312000
rect 135234 252308 135854 312000
rect 138954 252308 139574 312000
rect 141794 252308 142414 312000
rect 145514 252308 146134 312000
rect 149234 252308 149854 312000
rect 152954 252308 153574 312000
rect 155794 252308 156414 312000
rect 159514 252308 160134 312000
rect 163234 252308 163854 312000
rect 166954 252308 167574 312000
rect 169794 252308 170414 312000
rect 173514 252308 174134 451000
rect 177234 252308 177854 451000
rect 180954 252308 181574 451000
rect 183794 252308 184414 451000
rect 187514 252308 188134 451000
rect 191234 252308 191854 451000
rect 194954 252308 195574 451000
rect 197794 426000 198414 451000
rect 201514 426000 202134 707750
rect 205234 426000 205854 709670
rect 208954 426000 209574 711590
rect 211794 426000 212414 705830
rect 215514 426000 216134 707750
rect 219234 645308 219854 709670
rect 222954 645308 223574 711590
rect 225794 645308 226414 705830
rect 229514 645308 230134 707750
rect 233234 645308 233854 709670
rect 236954 645308 237574 711590
rect 239794 645308 240414 705830
rect 243514 645308 244134 707750
rect 247234 645308 247854 709670
rect 250954 645308 251574 711590
rect 253794 645308 254414 705830
rect 257514 645308 258134 707750
rect 261234 645308 261854 709670
rect 264954 645308 265574 711590
rect 267794 645308 268414 705830
rect 271514 645308 272134 707750
rect 275234 645308 275854 709670
rect 278954 645308 279574 711590
rect 281794 645308 282414 705830
rect 285514 645308 286134 707750
rect 289234 645308 289854 709670
rect 292954 645308 293574 711590
rect 295794 645308 296414 705830
rect 299514 645308 300134 707750
rect 303234 645308 303854 709670
rect 306954 645308 307574 711590
rect 309794 645308 310414 705830
rect 313514 645308 314134 707750
rect 317234 645308 317854 709670
rect 320954 645308 321574 711590
rect 323794 645308 324414 705830
rect 327514 645308 328134 707750
rect 331234 645308 331854 709670
rect 334954 645308 335574 711590
rect 337794 645308 338414 705830
rect 341514 645308 342134 707750
rect 345234 645308 345854 709670
rect 348954 645308 349574 711590
rect 351794 645308 352414 705830
rect 355514 645308 356134 707750
rect 219234 538308 219854 558000
rect 222954 538308 223574 558000
rect 225794 538308 226414 558000
rect 229514 538308 230134 558000
rect 233234 538308 233854 558000
rect 236954 538308 237574 558000
rect 239794 538308 240414 558000
rect 243514 538308 244134 558000
rect 247234 538308 247854 558000
rect 250954 538308 251574 558000
rect 253794 538308 254414 558000
rect 257514 538308 258134 558000
rect 261234 538308 261854 558000
rect 264954 538308 265574 558000
rect 267794 538308 268414 558000
rect 271514 538308 272134 558000
rect 275234 538308 275854 558000
rect 278954 538308 279574 558000
rect 281794 538308 282414 558000
rect 285514 538308 286134 558000
rect 289234 538308 289854 558000
rect 292954 538308 293574 558000
rect 295794 538308 296414 558000
rect 299514 538308 300134 558000
rect 303234 538308 303854 558000
rect 306954 538308 307574 558000
rect 309794 538308 310414 558000
rect 313514 538308 314134 558000
rect 317234 538308 317854 558000
rect 320954 538308 321574 558000
rect 323794 538308 324414 558000
rect 327514 538308 328134 558000
rect 331234 538308 331854 558000
rect 334954 538308 335574 558000
rect 337794 538308 338414 558000
rect 341514 538308 342134 558000
rect 345234 538308 345854 558000
rect 348954 538308 349574 558000
rect 351794 538308 352414 558000
rect 355514 538308 356134 558000
rect 219234 426000 219854 451000
rect 222954 426000 223574 451000
rect 225794 426000 226414 451000
rect 229514 426000 230134 451000
rect 233234 426000 233854 451000
rect 236954 426000 237574 451000
rect 239794 426000 240414 451000
rect 243514 426000 244134 451000
rect 247234 426000 247854 451000
rect 250954 426000 251574 451000
rect 253794 426000 254414 451000
rect 257514 426000 258134 451000
rect 261234 426000 261854 451000
rect 264954 426000 265574 451000
rect 267794 426000 268414 451000
rect 271514 426000 272134 451000
rect 275234 426000 275854 451000
rect 278954 426000 279574 451000
rect 281794 426000 282414 451000
rect 285514 426000 286134 451000
rect 289234 426000 289854 451000
rect 292954 426000 293574 451000
rect 295794 426000 296414 451000
rect 299514 426000 300134 451000
rect 303234 426000 303854 451000
rect 306954 426000 307574 451000
rect 309794 426000 310414 451000
rect 313514 426000 314134 451000
rect 317234 426000 317854 451000
rect 320954 426000 321574 451000
rect 197794 252308 198414 275000
rect 57794 145308 58414 165000
rect 61514 145308 62134 165000
rect 65234 145308 65854 165000
rect 68954 145308 69574 165000
rect 71794 145308 72414 165000
rect 75514 145308 76134 165000
rect 79234 145308 79854 165000
rect 82954 145308 83574 165000
rect 85794 145308 86414 165000
rect 89514 145308 90134 165000
rect 93234 145308 93854 165000
rect 96954 145308 97574 165000
rect 99794 145308 100414 165000
rect 103514 145308 104134 165000
rect 107234 145308 107854 165000
rect 110954 145308 111574 165000
rect 113794 145308 114414 165000
rect 117514 145308 118134 165000
rect 121234 145308 121854 165000
rect 124954 145308 125574 165000
rect 127794 145308 128414 165000
rect 131514 145308 132134 165000
rect 135234 145308 135854 165000
rect 138954 145308 139574 165000
rect 141794 145308 142414 165000
rect 145514 145308 146134 165000
rect 149234 145308 149854 165000
rect 152954 145308 153574 165000
rect 155794 145308 156414 165000
rect 159514 145308 160134 165000
rect 163234 145308 163854 165000
rect 166954 145308 167574 165000
rect 169794 145308 170414 165000
rect 173514 145308 174134 165000
rect 177234 145308 177854 165000
rect 180954 145308 181574 165000
rect 183794 145308 184414 165000
rect 187514 145308 188134 165000
rect 191234 145308 191854 165000
rect 194954 145308 195574 165000
rect 197794 145308 198414 165000
rect 57794 -1894 58414 58000
rect 61514 -3814 62134 58000
rect 65234 -5734 65854 58000
rect 68954 -7654 69574 58000
rect 71794 -1894 72414 58000
rect 75514 -3814 76134 58000
rect 79234 -5734 79854 58000
rect 82954 -7654 83574 58000
rect 85794 -1894 86414 58000
rect 89514 -3814 90134 58000
rect 93234 -5734 93854 58000
rect 96954 -7654 97574 58000
rect 99794 -1894 100414 58000
rect 103514 -3814 104134 58000
rect 107234 -5734 107854 58000
rect 110954 -7654 111574 58000
rect 113794 -1894 114414 58000
rect 117514 -3814 118134 58000
rect 121234 -5734 121854 58000
rect 124954 -7654 125574 58000
rect 127794 -1894 128414 58000
rect 131514 -3814 132134 58000
rect 135234 -5734 135854 58000
rect 138954 -7654 139574 58000
rect 141794 -1894 142414 58000
rect 145514 -3814 146134 58000
rect 149234 -5734 149854 58000
rect 152954 -7654 153574 58000
rect 155794 -1894 156414 58000
rect 159514 -3814 160134 58000
rect 163234 -5734 163854 58000
rect 166954 -7654 167574 58000
rect 169794 -1894 170414 58000
rect 173514 -3814 174134 58000
rect 177234 -5734 177854 58000
rect 180954 -7654 181574 58000
rect 183794 -1894 184414 58000
rect 187514 -3814 188134 58000
rect 191234 -5734 191854 58000
rect 194954 -7654 195574 58000
rect 197794 -1894 198414 58000
rect 201514 -3814 202134 275000
rect 205234 -5734 205854 275000
rect 208954 -7654 209574 275000
rect 211794 -1894 212414 275000
rect 215514 -3814 216134 275000
rect 219234 252308 219854 275000
rect 222954 252308 223574 275000
rect 225794 252308 226414 275000
rect 229514 252308 230134 275000
rect 233234 252308 233854 275000
rect 236954 252308 237574 275000
rect 239794 252308 240414 275000
rect 243514 252308 244134 275000
rect 247234 252308 247854 275000
rect 250954 252308 251574 275000
rect 253794 252308 254414 275000
rect 257514 252308 258134 275000
rect 261234 252308 261854 275000
rect 264954 252308 265574 275000
rect 267794 252308 268414 275000
rect 271514 252308 272134 275000
rect 275234 252308 275854 275000
rect 278954 252308 279574 275000
rect 281794 252308 282414 275000
rect 285514 252308 286134 275000
rect 289234 252308 289854 275000
rect 292954 252308 293574 275000
rect 295794 252308 296414 275000
rect 299514 252308 300134 275000
rect 303234 252308 303854 275000
rect 306954 252308 307574 275000
rect 309794 252308 310414 275000
rect 313514 252308 314134 275000
rect 317234 252308 317854 275000
rect 320954 252308 321574 275000
rect 323794 252308 324414 451000
rect 327514 252308 328134 451000
rect 331234 252308 331854 451000
rect 334954 252308 335574 451000
rect 337794 252308 338414 451000
rect 341514 252308 342134 451000
rect 345234 252308 345854 451000
rect 348954 252308 349574 451000
rect 351794 252308 352414 451000
rect 355514 252308 356134 451000
rect 359234 429099 359854 709670
rect 362954 429099 363574 711590
rect 365794 429099 366414 705830
rect 369514 429099 370134 707750
rect 373234 429099 373854 709670
rect 376954 429099 377574 711590
rect 379794 645308 380414 705830
rect 383514 645308 384134 707750
rect 387234 645308 387854 709670
rect 390954 645308 391574 711590
rect 393794 645308 394414 705830
rect 397514 645308 398134 707750
rect 401234 645308 401854 709670
rect 404954 645308 405574 711590
rect 407794 645308 408414 705830
rect 411514 645308 412134 707750
rect 415234 645308 415854 709670
rect 418954 645308 419574 711590
rect 421794 645308 422414 705830
rect 425514 645308 426134 707750
rect 429234 645308 429854 709670
rect 432954 645308 433574 711590
rect 435794 645308 436414 705830
rect 439514 645308 440134 707750
rect 443234 645308 443854 709670
rect 446954 645308 447574 711590
rect 449794 645308 450414 705830
rect 453514 645308 454134 707750
rect 457234 645308 457854 709670
rect 460954 645308 461574 711590
rect 463794 645308 464414 705830
rect 467514 645308 468134 707750
rect 471234 645308 471854 709670
rect 474954 645308 475574 711590
rect 477794 645308 478414 705830
rect 481514 645308 482134 707750
rect 485234 645308 485854 709670
rect 488954 645308 489574 711590
rect 491794 645308 492414 705830
rect 495514 645308 496134 707750
rect 499234 645308 499854 709670
rect 502954 645308 503574 711590
rect 505794 645308 506414 705830
rect 509514 645308 510134 707750
rect 513234 645308 513854 709670
rect 516954 645308 517574 711590
rect 379794 538308 380414 558000
rect 383514 538308 384134 558000
rect 387234 538308 387854 558000
rect 390954 538308 391574 558000
rect 393794 538308 394414 558000
rect 397514 538308 398134 558000
rect 401234 538308 401854 558000
rect 404954 538308 405574 558000
rect 407794 538308 408414 558000
rect 411514 538308 412134 558000
rect 415234 538308 415854 558000
rect 418954 538308 419574 558000
rect 421794 538308 422414 558000
rect 425514 538308 426134 558000
rect 429234 538308 429854 558000
rect 432954 538308 433574 558000
rect 435794 538308 436414 558000
rect 439514 538308 440134 558000
rect 443234 538308 443854 558000
rect 446954 538308 447574 558000
rect 449794 538308 450414 558000
rect 453514 538308 454134 558000
rect 457234 538308 457854 558000
rect 460954 538308 461574 558000
rect 463794 538308 464414 558000
rect 467514 538308 468134 558000
rect 471234 538308 471854 558000
rect 474954 538308 475574 558000
rect 477794 538308 478414 558000
rect 481514 538308 482134 558000
rect 485234 538308 485854 558000
rect 488954 538308 489574 558000
rect 491794 538308 492414 558000
rect 495514 538308 496134 558000
rect 499234 538308 499854 558000
rect 502954 538308 503574 558000
rect 505794 538308 506414 558000
rect 509514 538308 510134 558000
rect 513234 538308 513854 558000
rect 516954 538308 517574 558000
rect 379794 429099 380414 451000
rect 383514 429099 384134 451000
rect 387234 429099 387854 451000
rect 390954 429099 391574 451000
rect 393794 429099 394414 451000
rect 397514 429099 398134 451000
rect 401234 429099 401854 451000
rect 404954 429099 405574 451000
rect 407794 429099 408414 451000
rect 411514 429099 412134 451000
rect 415234 429099 415854 451000
rect 418954 429099 419574 451000
rect 421794 429099 422414 451000
rect 359234 342099 359854 362000
rect 362954 342099 363574 362000
rect 365794 342099 366414 362000
rect 369514 342099 370134 362000
rect 373234 342099 373854 362000
rect 376954 342099 377574 362000
rect 379794 342099 380414 362000
rect 383514 342099 384134 362000
rect 387234 342099 387854 362000
rect 390954 342099 391574 362000
rect 393794 342099 394414 362000
rect 397514 342099 398134 362000
rect 401234 342099 401854 362000
rect 404954 342099 405574 362000
rect 407794 342099 408414 362000
rect 411514 342099 412134 362000
rect 415234 342099 415854 362000
rect 418954 342099 419574 362000
rect 421794 342099 422414 362000
rect 219234 145308 219854 165000
rect 222954 145308 223574 165000
rect 225794 145308 226414 165000
rect 229514 145308 230134 165000
rect 233234 145308 233854 165000
rect 236954 145308 237574 165000
rect 239794 145308 240414 165000
rect 243514 145308 244134 165000
rect 247234 145308 247854 165000
rect 250954 145308 251574 165000
rect 253794 145308 254414 165000
rect 257514 145308 258134 165000
rect 261234 145308 261854 165000
rect 264954 145308 265574 165000
rect 267794 145308 268414 165000
rect 271514 145308 272134 165000
rect 275234 145308 275854 165000
rect 278954 145308 279574 165000
rect 281794 145308 282414 165000
rect 285514 145308 286134 165000
rect 289234 145308 289854 165000
rect 292954 145308 293574 165000
rect 295794 145308 296414 165000
rect 299514 145308 300134 165000
rect 303234 145308 303854 165000
rect 306954 145308 307574 165000
rect 309794 145308 310414 165000
rect 313514 145308 314134 165000
rect 317234 145308 317854 165000
rect 320954 145308 321574 165000
rect 323794 145308 324414 165000
rect 327514 145308 328134 165000
rect 331234 145308 331854 165000
rect 334954 145308 335574 165000
rect 337794 145308 338414 165000
rect 341514 145308 342134 165000
rect 345234 145308 345854 165000
rect 348954 145308 349574 165000
rect 351794 145308 352414 165000
rect 355514 145308 356134 165000
rect 219234 -5734 219854 58000
rect 222954 -7654 223574 58000
rect 225794 -1894 226414 58000
rect 229514 -3814 230134 58000
rect 233234 -5734 233854 58000
rect 236954 -7654 237574 58000
rect 239794 -1894 240414 58000
rect 243514 -3814 244134 58000
rect 247234 -5734 247854 58000
rect 250954 -7654 251574 58000
rect 253794 -1894 254414 58000
rect 257514 -3814 258134 58000
rect 261234 -5734 261854 58000
rect 264954 -7654 265574 58000
rect 267794 -1894 268414 58000
rect 271514 -3814 272134 58000
rect 275234 -5734 275854 58000
rect 278954 -7654 279574 58000
rect 281794 -1894 282414 58000
rect 285514 -3814 286134 58000
rect 289234 -5734 289854 58000
rect 292954 -7654 293574 58000
rect 295794 -1894 296414 58000
rect 299514 -3814 300134 58000
rect 303234 -5734 303854 58000
rect 306954 -7654 307574 58000
rect 309794 -1894 310414 58000
rect 313514 -3814 314134 58000
rect 317234 -5734 317854 58000
rect 320954 -7654 321574 58000
rect 323794 -1894 324414 58000
rect 327514 -3814 328134 58000
rect 331234 -5734 331854 58000
rect 334954 -7654 335574 58000
rect 337794 -1894 338414 58000
rect 341514 -3814 342134 58000
rect 345234 -5734 345854 58000
rect 348954 -7654 349574 58000
rect 351794 -1894 352414 58000
rect 355514 -3814 356134 58000
rect 359234 -5734 359854 275000
rect 362954 -7654 363574 275000
rect 365794 -1894 366414 275000
rect 369514 -3814 370134 275000
rect 373234 -5734 373854 275000
rect 376954 -7654 377574 275000
rect 379794 252308 380414 275000
rect 383514 252308 384134 275000
rect 387234 252308 387854 275000
rect 390954 252308 391574 275000
rect 393794 252308 394414 275000
rect 397514 252308 398134 275000
rect 401234 252308 401854 275000
rect 404954 252308 405574 275000
rect 407794 252308 408414 275000
rect 411514 252308 412134 275000
rect 415234 252308 415854 275000
rect 418954 252308 419574 275000
rect 421794 252308 422414 275000
rect 425514 252308 426134 451000
rect 429234 252308 429854 451000
rect 432954 252308 433574 451000
rect 435794 252308 436414 451000
rect 439514 252308 440134 451000
rect 443234 252308 443854 451000
rect 446954 252308 447574 451000
rect 449794 429099 450414 451000
rect 453514 429099 454134 451000
rect 457234 429099 457854 451000
rect 460954 429099 461574 451000
rect 463794 429099 464414 451000
rect 467514 429099 468134 451000
rect 471234 429099 471854 451000
rect 474954 429099 475574 451000
rect 477794 429099 478414 451000
rect 481514 429099 482134 451000
rect 485234 429099 485854 451000
rect 488954 429099 489574 451000
rect 491794 429099 492414 451000
rect 495514 429099 496134 451000
rect 499234 429099 499854 451000
rect 502954 429099 503574 451000
rect 505794 429099 506414 451000
rect 509514 429099 510134 451000
rect 449794 252308 450414 362000
rect 453514 252308 454134 362000
rect 457234 252308 457854 362000
rect 460954 329000 461574 362000
rect 463794 329000 464414 362000
rect 467514 329000 468134 362000
rect 471234 329000 471854 362000
rect 474954 329000 475574 362000
rect 477794 329000 478414 362000
rect 481514 329000 482134 362000
rect 485234 329000 485854 362000
rect 488954 329000 489574 362000
rect 491794 329000 492414 362000
rect 495514 329000 496134 362000
rect 499234 329000 499854 362000
rect 502954 329000 503574 362000
rect 505794 329000 506414 362000
rect 509514 329000 510134 362000
rect 460954 252308 461574 275000
rect 463794 252308 464414 275000
rect 467514 252308 468134 275000
rect 471234 252308 471854 275000
rect 474954 252308 475574 275000
rect 477794 252308 478414 275000
rect 481514 252308 482134 275000
rect 485234 252308 485854 275000
rect 488954 252308 489574 275000
rect 491794 252308 492414 275000
rect 495514 252308 496134 275000
rect 499234 252308 499854 275000
rect 502954 252308 503574 275000
rect 505794 252308 506414 275000
rect 509514 252308 510134 275000
rect 513234 252308 513854 451000
rect 516954 252308 517574 451000
rect 379794 145308 380414 165000
rect 383514 145308 384134 165000
rect 387234 145308 387854 165000
rect 390954 145308 391574 165000
rect 393794 145308 394414 165000
rect 397514 145308 398134 165000
rect 401234 145308 401854 165000
rect 404954 145308 405574 165000
rect 407794 145308 408414 165000
rect 411514 145308 412134 165000
rect 415234 145308 415854 165000
rect 418954 145308 419574 165000
rect 421794 145308 422414 165000
rect 425514 145308 426134 165000
rect 429234 145308 429854 165000
rect 432954 145308 433574 165000
rect 435794 145308 436414 165000
rect 439514 145308 440134 165000
rect 443234 145308 443854 165000
rect 446954 145308 447574 165000
rect 449794 145308 450414 165000
rect 453514 145308 454134 165000
rect 457234 145308 457854 165000
rect 460954 145308 461574 165000
rect 463794 145308 464414 165000
rect 467514 145308 468134 165000
rect 471234 145308 471854 165000
rect 474954 145308 475574 165000
rect 477794 145308 478414 165000
rect 481514 145308 482134 165000
rect 485234 145308 485854 165000
rect 488954 145308 489574 165000
rect 491794 145308 492414 165000
rect 495514 145308 496134 165000
rect 499234 145308 499854 165000
rect 502954 145308 503574 165000
rect 505794 145308 506414 165000
rect 509514 145308 510134 165000
rect 513234 145308 513854 165000
rect 516954 145308 517574 165000
rect 379794 -1894 380414 58000
rect 383514 -3814 384134 58000
rect 387234 -5734 387854 58000
rect 390954 -7654 391574 58000
rect 393794 -1894 394414 58000
rect 397514 -3814 398134 58000
rect 401234 -5734 401854 58000
rect 404954 -7654 405574 58000
rect 407794 -1894 408414 58000
rect 411514 -3814 412134 58000
rect 415234 -5734 415854 58000
rect 418954 -7654 419574 58000
rect 421794 -1894 422414 58000
rect 425514 -3814 426134 58000
rect 429234 -5734 429854 58000
rect 432954 -7654 433574 58000
rect 435794 -1894 436414 58000
rect 439514 -3814 440134 58000
rect 443234 -5734 443854 58000
rect 446954 -7654 447574 58000
rect 449794 -1894 450414 58000
rect 453514 -3814 454134 58000
rect 457234 -5734 457854 58000
rect 460954 -7654 461574 58000
rect 463794 -1894 464414 58000
rect 467514 -3814 468134 58000
rect 471234 -5734 471854 58000
rect 474954 -7654 475574 58000
rect 477794 -1894 478414 58000
rect 481514 -3814 482134 58000
rect 485234 -5734 485854 58000
rect 488954 -7654 489574 58000
rect 491794 -1894 492414 58000
rect 495514 -3814 496134 58000
rect 499234 -5734 499854 58000
rect 502954 -7654 503574 58000
rect 505794 -1894 506414 58000
rect 509514 -3814 510134 58000
rect 513234 -5734 513854 58000
rect 516954 -7654 517574 58000
rect 519794 -1894 520414 705830
rect 523514 -3814 524134 707750
rect 527234 -5734 527854 709670
rect 530954 -7654 531574 711590
rect 533794 -1894 534414 705830
rect 537514 -3814 538134 707750
rect 541234 -5734 541854 709670
rect 544954 -7654 545574 711590
rect 547794 -1894 548414 705830
rect 551514 -3814 552134 707750
rect 555234 -5734 555854 709670
rect 558954 -7654 559574 711590
rect 561794 -1894 562414 705830
rect 565514 -3814 566134 707750
rect 569234 -5734 569854 709670
rect 572954 -7654 573574 711590
rect 575794 -1894 576414 705830
rect 579514 -3814 580134 707750
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 57099 645228 57714 700365
rect 58494 645228 61434 700365
rect 62214 645228 65154 700365
rect 65934 645228 68874 700365
rect 69654 645228 71714 700365
rect 72494 645228 75434 700365
rect 76214 645228 79154 700365
rect 79934 645228 82874 700365
rect 83654 645228 85714 700365
rect 86494 645228 89434 700365
rect 90214 645228 93154 700365
rect 93934 645228 96874 700365
rect 97654 645228 99714 700365
rect 100494 645228 103434 700365
rect 104214 645228 107154 700365
rect 107934 645228 110874 700365
rect 111654 645228 113714 700365
rect 114494 645228 117434 700365
rect 118214 645228 121154 700365
rect 121934 645228 124874 700365
rect 125654 645228 127714 700365
rect 128494 645228 131434 700365
rect 132214 645228 135154 700365
rect 135934 645228 138874 700365
rect 139654 645228 141714 700365
rect 142494 645228 145434 700365
rect 146214 645228 149154 700365
rect 149934 645228 152874 700365
rect 153654 645228 155714 700365
rect 156494 645228 159434 700365
rect 160214 645228 163154 700365
rect 163934 645228 166874 700365
rect 167654 645228 169714 700365
rect 170494 645228 173434 700365
rect 174214 645228 177154 700365
rect 177934 645228 180874 700365
rect 181654 645228 183714 700365
rect 184494 645228 187434 700365
rect 188214 645228 191154 700365
rect 191934 645228 194874 700365
rect 195654 645228 197714 700365
rect 198494 645228 201434 700365
rect 57099 558080 201434 645228
rect 57099 538228 57714 558080
rect 58494 538228 61434 558080
rect 62214 538228 65154 558080
rect 65934 538228 68874 558080
rect 69654 538228 71714 558080
rect 72494 538228 75434 558080
rect 76214 538228 79154 558080
rect 79934 538228 82874 558080
rect 83654 538228 85714 558080
rect 86494 538228 89434 558080
rect 90214 538228 93154 558080
rect 93934 538228 96874 558080
rect 97654 538228 99714 558080
rect 100494 538228 103434 558080
rect 104214 538228 107154 558080
rect 107934 538228 110874 558080
rect 111654 538228 113714 558080
rect 114494 538228 117434 558080
rect 118214 538228 121154 558080
rect 121934 538228 124874 558080
rect 125654 538228 127714 558080
rect 128494 538228 131434 558080
rect 132214 538228 135154 558080
rect 135934 538228 138874 558080
rect 139654 538228 141714 558080
rect 142494 538228 145434 558080
rect 146214 538228 149154 558080
rect 149934 538228 152874 558080
rect 153654 538228 155714 558080
rect 156494 538228 159434 558080
rect 160214 538228 163154 558080
rect 163934 538228 166874 558080
rect 167654 538228 169714 558080
rect 170494 538228 173434 558080
rect 174214 538228 177154 558080
rect 177934 538228 180874 558080
rect 181654 538228 183714 558080
rect 184494 538228 187434 558080
rect 188214 538228 191154 558080
rect 191934 538228 194874 558080
rect 195654 538228 197714 558080
rect 198494 538228 201434 558080
rect 57099 451080 201434 538228
rect 57099 426953 57714 451080
rect 58494 426953 61434 451080
rect 62214 426953 65154 451080
rect 65934 426953 68874 451080
rect 69654 426953 71714 451080
rect 72494 426953 75434 451080
rect 76214 426953 79154 451080
rect 79934 426953 82874 451080
rect 83654 426953 85714 451080
rect 86494 426953 89434 451080
rect 90214 426953 93154 451080
rect 93934 426953 96874 451080
rect 97654 426953 99714 451080
rect 100494 426953 103434 451080
rect 104214 426953 107154 451080
rect 107934 426953 110874 451080
rect 111654 426953 113714 451080
rect 114494 426953 117434 451080
rect 118214 426953 121154 451080
rect 121934 426953 124874 451080
rect 125654 426953 127714 451080
rect 128494 426953 131434 451080
rect 132214 426953 135154 451080
rect 135934 426953 138874 451080
rect 139654 426953 141714 451080
rect 142494 426953 145434 451080
rect 146214 426953 149154 451080
rect 149934 426953 152874 451080
rect 153654 426953 155714 451080
rect 156494 426953 159434 451080
rect 160214 426953 163154 451080
rect 163934 426953 166874 451080
rect 167654 426953 169714 451080
rect 170494 426953 173434 451080
rect 57099 312080 173434 426953
rect 57099 252228 57714 312080
rect 58494 252228 61434 312080
rect 62214 252228 65154 312080
rect 65934 252228 68874 312080
rect 69654 252228 71714 312080
rect 72494 252228 75434 312080
rect 76214 252228 79154 312080
rect 79934 252228 82874 312080
rect 83654 252228 85714 312080
rect 86494 252228 89434 312080
rect 90214 252228 93154 312080
rect 93934 252228 96874 312080
rect 97654 252228 99714 312080
rect 100494 252228 103434 312080
rect 104214 252228 107154 312080
rect 107934 252228 110874 312080
rect 111654 252228 113714 312080
rect 114494 252228 117434 312080
rect 118214 252228 121154 312080
rect 121934 252228 124874 312080
rect 125654 252228 127714 312080
rect 128494 252228 131434 312080
rect 132214 252228 135154 312080
rect 135934 252228 138874 312080
rect 139654 252228 141714 312080
rect 142494 252228 145434 312080
rect 146214 252228 149154 312080
rect 149934 252228 152874 312080
rect 153654 252228 155714 312080
rect 156494 252228 159434 312080
rect 160214 252228 163154 312080
rect 163934 252228 166874 312080
rect 167654 252228 169714 312080
rect 170494 252228 173434 312080
rect 174214 252228 177154 451080
rect 177934 252228 180874 451080
rect 181654 252228 183714 451080
rect 184494 252228 187434 451080
rect 188214 252228 191154 451080
rect 191934 252228 194874 451080
rect 195654 425920 197714 451080
rect 198494 425920 201434 451080
rect 202214 425920 205154 700365
rect 205934 425920 208874 700365
rect 209654 425920 211714 700365
rect 212494 425920 215434 700365
rect 216214 645228 219154 700365
rect 219934 645228 222874 700365
rect 223654 645228 225714 700365
rect 226494 645228 229434 700365
rect 230214 645228 233154 700365
rect 233934 645228 236874 700365
rect 237654 645228 239714 700365
rect 240494 645228 243434 700365
rect 244214 645228 247154 700365
rect 247934 645228 250874 700365
rect 251654 645228 253714 700365
rect 254494 645228 257434 700365
rect 258214 645228 261154 700365
rect 261934 645228 264874 700365
rect 265654 645228 267714 700365
rect 268494 645228 271434 700365
rect 272214 645228 275154 700365
rect 275934 645228 278874 700365
rect 279654 645228 281714 700365
rect 282494 645228 285434 700365
rect 286214 645228 289154 700365
rect 289934 645228 292874 700365
rect 293654 645228 295714 700365
rect 296494 645228 299434 700365
rect 300214 645228 303154 700365
rect 303934 645228 306874 700365
rect 307654 645228 309714 700365
rect 310494 645228 313434 700365
rect 314214 645228 317154 700365
rect 317934 645228 320874 700365
rect 321654 645228 323714 700365
rect 324494 645228 327434 700365
rect 328214 645228 331154 700365
rect 331934 645228 334874 700365
rect 335654 645228 337714 700365
rect 338494 645228 341434 700365
rect 342214 645228 345154 700365
rect 345934 645228 348874 700365
rect 349654 645228 351714 700365
rect 352494 645228 355434 700365
rect 356214 645228 359154 700365
rect 216214 558080 359154 645228
rect 216214 538228 219154 558080
rect 219934 538228 222874 558080
rect 223654 538228 225714 558080
rect 226494 538228 229434 558080
rect 230214 538228 233154 558080
rect 233934 538228 236874 558080
rect 237654 538228 239714 558080
rect 240494 538228 243434 558080
rect 244214 538228 247154 558080
rect 247934 538228 250874 558080
rect 251654 538228 253714 558080
rect 254494 538228 257434 558080
rect 258214 538228 261154 558080
rect 261934 538228 264874 558080
rect 265654 538228 267714 558080
rect 268494 538228 271434 558080
rect 272214 538228 275154 558080
rect 275934 538228 278874 558080
rect 279654 538228 281714 558080
rect 282494 538228 285434 558080
rect 286214 538228 289154 558080
rect 289934 538228 292874 558080
rect 293654 538228 295714 558080
rect 296494 538228 299434 558080
rect 300214 538228 303154 558080
rect 303934 538228 306874 558080
rect 307654 538228 309714 558080
rect 310494 538228 313434 558080
rect 314214 538228 317154 558080
rect 317934 538228 320874 558080
rect 321654 538228 323714 558080
rect 324494 538228 327434 558080
rect 328214 538228 331154 558080
rect 331934 538228 334874 558080
rect 335654 538228 337714 558080
rect 338494 538228 341434 558080
rect 342214 538228 345154 558080
rect 345934 538228 348874 558080
rect 349654 538228 351714 558080
rect 352494 538228 355434 558080
rect 356214 538228 359154 558080
rect 216214 451080 359154 538228
rect 216214 425920 219154 451080
rect 219934 425920 222874 451080
rect 223654 425920 225714 451080
rect 226494 425920 229434 451080
rect 230214 425920 233154 451080
rect 233934 425920 236874 451080
rect 237654 425920 239714 451080
rect 240494 425920 243434 451080
rect 244214 425920 247154 451080
rect 247934 425920 250874 451080
rect 251654 425920 253714 451080
rect 254494 425920 257434 451080
rect 258214 425920 261154 451080
rect 261934 425920 264874 451080
rect 265654 425920 267714 451080
rect 268494 425920 271434 451080
rect 272214 425920 275154 451080
rect 275934 425920 278874 451080
rect 279654 425920 281714 451080
rect 282494 425920 285434 451080
rect 286214 425920 289154 451080
rect 289934 425920 292874 451080
rect 293654 425920 295714 451080
rect 296494 425920 299434 451080
rect 300214 425920 303154 451080
rect 303934 425920 306874 451080
rect 307654 425920 309714 451080
rect 310494 425920 313434 451080
rect 314214 425920 317154 451080
rect 317934 425920 320874 451080
rect 321654 425920 323714 451080
rect 195654 275080 323714 425920
rect 195654 252228 197714 275080
rect 198494 252228 201434 275080
rect 57099 165080 201434 252228
rect 57099 145228 57714 165080
rect 58494 145228 61434 165080
rect 62214 145228 65154 165080
rect 65934 145228 68874 165080
rect 69654 145228 71714 165080
rect 72494 145228 75434 165080
rect 76214 145228 79154 165080
rect 79934 145228 82874 165080
rect 83654 145228 85714 165080
rect 86494 145228 89434 165080
rect 90214 145228 93154 165080
rect 93934 145228 96874 165080
rect 97654 145228 99714 165080
rect 100494 145228 103434 165080
rect 104214 145228 107154 165080
rect 107934 145228 110874 165080
rect 111654 145228 113714 165080
rect 114494 145228 117434 165080
rect 118214 145228 121154 165080
rect 121934 145228 124874 165080
rect 125654 145228 127714 165080
rect 128494 145228 131434 165080
rect 132214 145228 135154 165080
rect 135934 145228 138874 165080
rect 139654 145228 141714 165080
rect 142494 145228 145434 165080
rect 146214 145228 149154 165080
rect 149934 145228 152874 165080
rect 153654 145228 155714 165080
rect 156494 145228 159434 165080
rect 160214 145228 163154 165080
rect 163934 145228 166874 165080
rect 167654 145228 169714 165080
rect 170494 145228 173434 165080
rect 174214 145228 177154 165080
rect 177934 145228 180874 165080
rect 181654 145228 183714 165080
rect 184494 145228 187434 165080
rect 188214 145228 191154 165080
rect 191934 145228 194874 165080
rect 195654 145228 197714 165080
rect 198494 145228 201434 165080
rect 57099 58080 201434 145228
rect 57099 11595 57714 58080
rect 58494 11595 61434 58080
rect 62214 11595 65154 58080
rect 65934 11595 68874 58080
rect 69654 11595 71714 58080
rect 72494 11595 75434 58080
rect 76214 11595 79154 58080
rect 79934 11595 82874 58080
rect 83654 11595 85714 58080
rect 86494 11595 89434 58080
rect 90214 11595 93154 58080
rect 93934 11595 96874 58080
rect 97654 11595 99714 58080
rect 100494 11595 103434 58080
rect 104214 11595 107154 58080
rect 107934 11595 110874 58080
rect 111654 11595 113714 58080
rect 114494 11595 117434 58080
rect 118214 11595 121154 58080
rect 121934 11595 124874 58080
rect 125654 11595 127714 58080
rect 128494 11595 131434 58080
rect 132214 11595 135154 58080
rect 135934 11595 138874 58080
rect 139654 11595 141714 58080
rect 142494 11595 145434 58080
rect 146214 11595 149154 58080
rect 149934 11595 152874 58080
rect 153654 11595 155714 58080
rect 156494 11595 159434 58080
rect 160214 11595 163154 58080
rect 163934 11595 166874 58080
rect 167654 11595 169714 58080
rect 170494 11595 173434 58080
rect 174214 11595 177154 58080
rect 177934 11595 180874 58080
rect 181654 11595 183714 58080
rect 184494 11595 187434 58080
rect 188214 11595 191154 58080
rect 191934 11595 194874 58080
rect 195654 11595 197714 58080
rect 198494 11595 201434 58080
rect 202214 11595 205154 275080
rect 205934 11595 208874 275080
rect 209654 11595 211714 275080
rect 212494 11595 215434 275080
rect 216214 252228 219154 275080
rect 219934 252228 222874 275080
rect 223654 252228 225714 275080
rect 226494 252228 229434 275080
rect 230214 252228 233154 275080
rect 233934 252228 236874 275080
rect 237654 252228 239714 275080
rect 240494 252228 243434 275080
rect 244214 252228 247154 275080
rect 247934 252228 250874 275080
rect 251654 252228 253714 275080
rect 254494 252228 257434 275080
rect 258214 252228 261154 275080
rect 261934 252228 264874 275080
rect 265654 252228 267714 275080
rect 268494 252228 271434 275080
rect 272214 252228 275154 275080
rect 275934 252228 278874 275080
rect 279654 252228 281714 275080
rect 282494 252228 285434 275080
rect 286214 252228 289154 275080
rect 289934 252228 292874 275080
rect 293654 252228 295714 275080
rect 296494 252228 299434 275080
rect 300214 252228 303154 275080
rect 303934 252228 306874 275080
rect 307654 252228 309714 275080
rect 310494 252228 313434 275080
rect 314214 252228 317154 275080
rect 317934 252228 320874 275080
rect 321654 252228 323714 275080
rect 324494 252228 327434 451080
rect 328214 252228 331154 451080
rect 331934 252228 334874 451080
rect 335654 252228 337714 451080
rect 338494 252228 341434 451080
rect 342214 252228 345154 451080
rect 345934 252228 348874 451080
rect 349654 252228 351714 451080
rect 352494 252228 355434 451080
rect 356214 429019 359154 451080
rect 359934 429019 362874 700365
rect 363654 429019 365714 700365
rect 366494 429019 369434 700365
rect 370214 429019 373154 700365
rect 373934 429019 376874 700365
rect 377654 645228 379714 700365
rect 380494 645228 383434 700365
rect 384214 645228 387154 700365
rect 387934 645228 390874 700365
rect 391654 645228 393714 700365
rect 394494 645228 397434 700365
rect 398214 645228 401154 700365
rect 401934 645228 404874 700365
rect 405654 645228 407714 700365
rect 408494 645228 411434 700365
rect 412214 645228 415154 700365
rect 415934 645228 418874 700365
rect 419654 645228 421714 700365
rect 422494 645228 425434 700365
rect 426214 645228 429154 700365
rect 429934 645228 432874 700365
rect 433654 645228 435714 700365
rect 436494 645228 439434 700365
rect 440214 645228 443154 700365
rect 443934 645228 446874 700365
rect 447654 645228 449714 700365
rect 450494 645228 453434 700365
rect 454214 645228 457154 700365
rect 457934 645228 460874 700365
rect 461654 645228 463714 700365
rect 464494 645228 467434 700365
rect 468214 645228 471154 700365
rect 471934 645228 474874 700365
rect 475654 645228 477714 700365
rect 478494 645228 481434 700365
rect 482214 645228 485154 700365
rect 485934 645228 488874 700365
rect 489654 645228 491714 700365
rect 492494 645228 495434 700365
rect 496214 645228 499154 700365
rect 499934 645228 502874 700365
rect 503654 645228 505714 700365
rect 506494 645228 509434 700365
rect 510214 645228 513154 700365
rect 513934 645228 516496 700365
rect 377654 558080 516496 645228
rect 377654 538228 379714 558080
rect 380494 538228 383434 558080
rect 384214 538228 387154 558080
rect 387934 538228 390874 558080
rect 391654 538228 393714 558080
rect 394494 538228 397434 558080
rect 398214 538228 401154 558080
rect 401934 538228 404874 558080
rect 405654 538228 407714 558080
rect 408494 538228 411434 558080
rect 412214 538228 415154 558080
rect 415934 538228 418874 558080
rect 419654 538228 421714 558080
rect 422494 538228 425434 558080
rect 426214 538228 429154 558080
rect 429934 538228 432874 558080
rect 433654 538228 435714 558080
rect 436494 538228 439434 558080
rect 440214 538228 443154 558080
rect 443934 538228 446874 558080
rect 447654 538228 449714 558080
rect 450494 538228 453434 558080
rect 454214 538228 457154 558080
rect 457934 538228 460874 558080
rect 461654 538228 463714 558080
rect 464494 538228 467434 558080
rect 468214 538228 471154 558080
rect 471934 538228 474874 558080
rect 475654 538228 477714 558080
rect 478494 538228 481434 558080
rect 482214 538228 485154 558080
rect 485934 538228 488874 558080
rect 489654 538228 491714 558080
rect 492494 538228 495434 558080
rect 496214 538228 499154 558080
rect 499934 538228 502874 558080
rect 503654 538228 505714 558080
rect 506494 538228 509434 558080
rect 510214 538228 513154 558080
rect 513934 538228 516496 558080
rect 377654 451080 516496 538228
rect 377654 429019 379714 451080
rect 380494 429019 383434 451080
rect 384214 429019 387154 451080
rect 387934 429019 390874 451080
rect 391654 429019 393714 451080
rect 394494 429019 397434 451080
rect 398214 429019 401154 451080
rect 401934 429019 404874 451080
rect 405654 429019 407714 451080
rect 408494 429019 411434 451080
rect 412214 429019 415154 451080
rect 415934 429019 418874 451080
rect 419654 429019 421714 451080
rect 422494 429019 425434 451080
rect 356214 362080 425434 429019
rect 356214 342019 359154 362080
rect 359934 342019 362874 362080
rect 363654 342019 365714 362080
rect 366494 342019 369434 362080
rect 370214 342019 373154 362080
rect 373934 342019 376874 362080
rect 377654 342019 379714 362080
rect 380494 342019 383434 362080
rect 384214 342019 387154 362080
rect 387934 342019 390874 362080
rect 391654 342019 393714 362080
rect 394494 342019 397434 362080
rect 398214 342019 401154 362080
rect 401934 342019 404874 362080
rect 405654 342019 407714 362080
rect 408494 342019 411434 362080
rect 412214 342019 415154 362080
rect 415934 342019 418874 362080
rect 419654 342019 421714 362080
rect 422494 342019 425434 362080
rect 356214 275080 425434 342019
rect 356214 252228 359154 275080
rect 216214 165080 359154 252228
rect 216214 145228 219154 165080
rect 219934 145228 222874 165080
rect 223654 145228 225714 165080
rect 226494 145228 229434 165080
rect 230214 145228 233154 165080
rect 233934 145228 236874 165080
rect 237654 145228 239714 165080
rect 240494 145228 243434 165080
rect 244214 145228 247154 165080
rect 247934 145228 250874 165080
rect 251654 145228 253714 165080
rect 254494 145228 257434 165080
rect 258214 145228 261154 165080
rect 261934 145228 264874 165080
rect 265654 145228 267714 165080
rect 268494 145228 271434 165080
rect 272214 145228 275154 165080
rect 275934 145228 278874 165080
rect 279654 145228 281714 165080
rect 282494 145228 285434 165080
rect 286214 145228 289154 165080
rect 289934 145228 292874 165080
rect 293654 145228 295714 165080
rect 296494 145228 299434 165080
rect 300214 145228 303154 165080
rect 303934 145228 306874 165080
rect 307654 145228 309714 165080
rect 310494 145228 313434 165080
rect 314214 145228 317154 165080
rect 317934 145228 320874 165080
rect 321654 145228 323714 165080
rect 324494 145228 327434 165080
rect 328214 145228 331154 165080
rect 331934 145228 334874 165080
rect 335654 145228 337714 165080
rect 338494 145228 341434 165080
rect 342214 145228 345154 165080
rect 345934 145228 348874 165080
rect 349654 145228 351714 165080
rect 352494 145228 355434 165080
rect 356214 145228 359154 165080
rect 216214 58080 359154 145228
rect 216214 11595 219154 58080
rect 219934 11595 222874 58080
rect 223654 11595 225714 58080
rect 226494 11595 229434 58080
rect 230214 11595 233154 58080
rect 233934 11595 236874 58080
rect 237654 11595 239714 58080
rect 240494 11595 243434 58080
rect 244214 11595 247154 58080
rect 247934 11595 250874 58080
rect 251654 11595 253714 58080
rect 254494 11595 257434 58080
rect 258214 11595 261154 58080
rect 261934 11595 264874 58080
rect 265654 11595 267714 58080
rect 268494 11595 271434 58080
rect 272214 11595 275154 58080
rect 275934 11595 278874 58080
rect 279654 11595 281714 58080
rect 282494 11595 285434 58080
rect 286214 11595 289154 58080
rect 289934 11595 292874 58080
rect 293654 11595 295714 58080
rect 296494 11595 299434 58080
rect 300214 11595 303154 58080
rect 303934 11595 306874 58080
rect 307654 11595 309714 58080
rect 310494 11595 313434 58080
rect 314214 11595 317154 58080
rect 317934 11595 320874 58080
rect 321654 11595 323714 58080
rect 324494 11595 327434 58080
rect 328214 11595 331154 58080
rect 331934 11595 334874 58080
rect 335654 11595 337714 58080
rect 338494 11595 341434 58080
rect 342214 11595 345154 58080
rect 345934 11595 348874 58080
rect 349654 11595 351714 58080
rect 352494 11595 355434 58080
rect 356214 11595 359154 58080
rect 359934 11595 362874 275080
rect 363654 11595 365714 275080
rect 366494 11595 369434 275080
rect 370214 11595 373154 275080
rect 373934 11595 376874 275080
rect 377654 252228 379714 275080
rect 380494 252228 383434 275080
rect 384214 252228 387154 275080
rect 387934 252228 390874 275080
rect 391654 252228 393714 275080
rect 394494 252228 397434 275080
rect 398214 252228 401154 275080
rect 401934 252228 404874 275080
rect 405654 252228 407714 275080
rect 408494 252228 411434 275080
rect 412214 252228 415154 275080
rect 415934 252228 418874 275080
rect 419654 252228 421714 275080
rect 422494 252228 425434 275080
rect 426214 252228 429154 451080
rect 429934 252228 432874 451080
rect 433654 252228 435714 451080
rect 436494 252228 439434 451080
rect 440214 252228 443154 451080
rect 443934 252228 446874 451080
rect 447654 429019 449714 451080
rect 450494 429019 453434 451080
rect 454214 429019 457154 451080
rect 457934 429019 460874 451080
rect 461654 429019 463714 451080
rect 464494 429019 467434 451080
rect 468214 429019 471154 451080
rect 471934 429019 474874 451080
rect 475654 429019 477714 451080
rect 478494 429019 481434 451080
rect 482214 429019 485154 451080
rect 485934 429019 488874 451080
rect 489654 429019 491714 451080
rect 492494 429019 495434 451080
rect 496214 429019 499154 451080
rect 499934 429019 502874 451080
rect 503654 429019 505714 451080
rect 506494 429019 509434 451080
rect 510214 429019 513154 451080
rect 447654 362080 513154 429019
rect 447654 252228 449714 362080
rect 450494 252228 453434 362080
rect 454214 252228 457154 362080
rect 457934 328920 460874 362080
rect 461654 328920 463714 362080
rect 464494 328920 467434 362080
rect 468214 328920 471154 362080
rect 471934 328920 474874 362080
rect 475654 328920 477714 362080
rect 478494 328920 481434 362080
rect 482214 328920 485154 362080
rect 485934 328920 488874 362080
rect 489654 328920 491714 362080
rect 492494 328920 495434 362080
rect 496214 328920 499154 362080
rect 499934 328920 502874 362080
rect 503654 328920 505714 362080
rect 506494 328920 509434 362080
rect 510214 328920 513154 362080
rect 457934 275080 513154 328920
rect 457934 252228 460874 275080
rect 461654 252228 463714 275080
rect 464494 252228 467434 275080
rect 468214 252228 471154 275080
rect 471934 252228 474874 275080
rect 475654 252228 477714 275080
rect 478494 252228 481434 275080
rect 482214 252228 485154 275080
rect 485934 252228 488874 275080
rect 489654 252228 491714 275080
rect 492494 252228 495434 275080
rect 496214 252228 499154 275080
rect 499934 252228 502874 275080
rect 503654 252228 505714 275080
rect 506494 252228 509434 275080
rect 510214 252228 513154 275080
rect 513934 252228 516496 451080
rect 377654 165080 516496 252228
rect 377654 145228 379714 165080
rect 380494 145228 383434 165080
rect 384214 145228 387154 165080
rect 387934 145228 390874 165080
rect 391654 145228 393714 165080
rect 394494 145228 397434 165080
rect 398214 145228 401154 165080
rect 401934 145228 404874 165080
rect 405654 145228 407714 165080
rect 408494 145228 411434 165080
rect 412214 145228 415154 165080
rect 415934 145228 418874 165080
rect 419654 145228 421714 165080
rect 422494 145228 425434 165080
rect 426214 145228 429154 165080
rect 429934 145228 432874 165080
rect 433654 145228 435714 165080
rect 436494 145228 439434 165080
rect 440214 145228 443154 165080
rect 443934 145228 446874 165080
rect 447654 145228 449714 165080
rect 450494 145228 453434 165080
rect 454214 145228 457154 165080
rect 457934 145228 460874 165080
rect 461654 145228 463714 165080
rect 464494 145228 467434 165080
rect 468214 145228 471154 165080
rect 471934 145228 474874 165080
rect 475654 145228 477714 165080
rect 478494 145228 481434 165080
rect 482214 145228 485154 165080
rect 485934 145228 488874 165080
rect 489654 145228 491714 165080
rect 492494 145228 495434 165080
rect 496214 145228 499154 165080
rect 499934 145228 502874 165080
rect 503654 145228 505714 165080
rect 506494 145228 509434 165080
rect 510214 145228 513154 165080
rect 513934 145228 516496 165080
rect 377654 58080 516496 145228
rect 377654 11595 379714 58080
rect 380494 11595 383434 58080
rect 384214 11595 387154 58080
rect 387934 11595 390874 58080
rect 391654 11595 393714 58080
rect 394494 11595 397434 58080
rect 398214 11595 401154 58080
rect 401934 11595 404874 58080
rect 405654 11595 407714 58080
rect 408494 11595 411434 58080
rect 412214 11595 415154 58080
rect 415934 11595 418874 58080
rect 419654 11595 421714 58080
rect 422494 11595 425434 58080
rect 426214 11595 429154 58080
rect 429934 11595 432874 58080
rect 433654 11595 435714 58080
rect 436494 11595 439434 58080
rect 440214 11595 443154 58080
rect 443934 11595 446874 58080
rect 447654 11595 449714 58080
rect 450494 11595 453434 58080
rect 454214 11595 457154 58080
rect 457934 11595 460874 58080
rect 461654 11595 463714 58080
rect 464494 11595 467434 58080
rect 468214 11595 471154 58080
rect 471934 11595 474874 58080
rect 475654 11595 477714 58080
rect 478494 11595 481434 58080
rect 482214 11595 485154 58080
rect 485934 11595 488874 58080
rect 489654 11595 491714 58080
rect 492494 11595 495434 58080
rect 496214 11595 499154 58080
rect 499934 11595 502874 58080
rect 503654 11595 505714 58080
rect 506494 11595 509434 58080
rect 510214 11595 513154 58080
rect 513934 11595 516496 58080
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 700026 592650 700646
rect -6806 696306 590730 696926
rect -4886 692586 588810 693206
rect -2966 688866 586890 689486
rect -8726 686026 592650 686646
rect -6806 682306 590730 682926
rect -4886 678586 588810 679206
rect -2966 674866 586890 675486
rect -8726 672026 592650 672646
rect -6806 668306 590730 668926
rect -4886 664586 588810 665206
rect -2966 660866 586890 661486
rect -8726 658026 592650 658646
rect -6806 654306 590730 654926
rect -4886 650586 588810 651206
rect -2966 646866 586890 647486
rect -8726 644026 592650 644646
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -2966 632866 586890 633486
rect -8726 630026 592650 630646
rect -6806 626306 590730 626926
rect -4886 622586 588810 623206
rect -2966 618866 586890 619486
rect -8726 616026 592650 616646
rect -6806 612306 590730 612926
rect -4886 608586 588810 609206
rect -2966 604866 586890 605486
rect -8726 602026 592650 602646
rect -6806 598306 590730 598926
rect -4886 594586 588810 595206
rect -2966 590866 586890 591486
rect -8726 588026 592650 588646
rect -6806 584306 590730 584926
rect -4886 580586 588810 581206
rect -2966 576866 586890 577486
rect -8726 574026 592650 574646
rect -6806 570306 590730 570926
rect -4886 566586 588810 567206
rect -2966 562866 586890 563486
rect -8726 560026 592650 560646
rect -6806 556306 590730 556926
rect -4886 552586 588810 553206
rect -2966 548866 586890 549486
rect 57794 547926 506414 548546
rect 82954 546966 503574 547586
rect -8726 546026 592650 546646
rect -6806 542306 590730 542926
rect -4886 538586 588810 539206
rect -2966 534866 586890 535486
rect -8726 532026 592650 532646
rect -6806 528306 590730 528926
rect -4886 524586 588810 525206
rect -2966 520866 586890 521486
rect -8726 518026 592650 518646
rect -6806 514306 590730 514926
rect -4886 510586 588810 511206
rect -2966 506866 586890 507486
rect -8726 504026 592650 504646
rect -6806 500306 590730 500926
rect -4886 496586 588810 497206
rect -2966 492866 586890 493486
rect -8726 490026 592650 490646
rect -6806 486306 590730 486926
rect -4886 482586 588810 483206
rect -2966 478866 586890 479486
rect -8726 476026 592650 476646
rect -6806 472306 590730 472926
rect -4886 468586 588810 469206
rect -2966 464866 586890 465486
rect -8726 462026 592650 462646
rect -6806 458306 590730 458926
rect -4886 454586 588810 455206
rect -2966 450866 586890 451486
rect -8726 448026 592650 448646
rect -6806 444306 590730 444926
rect -4886 440586 588810 441206
rect 61514 439646 146134 440266
rect 397514 439646 510134 440266
rect 57794 437806 170414 438426
rect 197794 437806 310414 438426
rect 393794 437806 506414 438426
rect -2966 436866 586890 437486
rect -8726 434026 592650 434646
rect -6806 430306 590730 430926
rect -4886 426586 588810 427206
rect -2966 422866 586890 423486
rect -8726 420026 592650 420646
rect -6806 416306 590730 416926
rect -4886 412586 588810 413206
rect -2966 408866 586890 409486
rect -8726 406026 592650 406646
rect -6806 402306 590730 402926
rect -4886 398586 588810 399206
rect -2966 394866 586890 395486
rect -8726 392026 592650 392646
rect -6806 388306 590730 388926
rect -4886 384586 588810 385206
rect -2966 380866 586890 381486
rect -8726 378026 592650 378646
rect -6806 374306 590730 374926
rect -4886 370586 588810 371206
rect -2966 366866 586890 367486
rect -8726 364026 592650 364646
rect -6806 360306 590730 360926
rect -4886 356586 588810 357206
rect -2966 352866 586890 353486
rect 365794 351926 422414 352546
rect 362954 350966 419574 351586
rect -8726 350026 592650 350646
rect -6806 346306 590730 346926
rect -4886 342586 588810 343206
rect -2966 338866 586890 339486
rect -8726 336026 592650 336646
rect -6806 332306 590730 332926
rect -4886 328586 588810 329206
rect -2966 324866 586890 325486
rect -8726 322026 592650 322646
rect -6806 318306 590730 318926
rect -4886 314586 588810 315206
rect -2966 310866 586890 311486
rect -8726 308026 592650 308646
rect -6806 304306 590730 304926
rect -4886 300586 588810 301206
rect -2966 296866 586890 297486
rect -8726 294026 592650 294646
rect -6806 290306 590730 290926
rect -4886 286586 588810 287206
rect -2966 282866 586890 283486
rect -8726 280026 592650 280646
rect -6806 276306 590730 276926
rect -4886 272586 588810 273206
rect -2966 268866 586890 269486
rect -8726 266026 592650 266646
rect 222954 265086 307574 265706
rect 390954 265086 503574 265706
rect 219234 263246 303854 263866
rect 387234 263246 499854 263866
rect -6806 262306 590730 262926
rect -4886 258586 588810 259206
rect -2966 254866 586890 255486
rect -8726 252026 592650 252646
rect -6806 248306 590730 248926
rect -4886 244586 588810 245206
rect -2966 240866 586890 241486
rect -8726 238026 592650 238646
rect -6806 234306 590730 234926
rect -4886 230586 588810 231206
rect -2966 226866 586890 227486
rect -8726 224026 592650 224646
rect -6806 220306 590730 220926
rect -4886 216586 588810 217206
rect -2966 212866 586890 213486
rect -8726 210026 592650 210646
rect -6806 206306 590730 206926
rect -4886 202586 588810 203206
rect -2966 198866 586890 199486
rect -8726 196026 592650 196646
rect -6806 192306 590730 192926
rect -4886 188586 588810 189206
rect -2966 184866 586890 185486
rect -8726 182026 592650 182646
rect -6806 178306 590730 178926
rect -4886 174586 588810 175206
rect -2966 170866 586890 171486
rect -8726 168026 592650 168646
rect -6806 164306 590730 164926
rect -4886 160586 588810 161206
rect -2966 156866 586890 157486
rect 57794 155926 506414 156546
rect 82954 154966 503574 155586
rect -8726 154026 592650 154646
rect -6806 150306 590730 150926
rect -4886 146586 588810 147206
rect -2966 142866 586890 143486
rect -8726 140026 592650 140646
rect -6806 136306 590730 136926
rect -4886 132586 588810 133206
rect -2966 128866 586890 129486
rect -8726 126026 592650 126646
rect -6806 122306 590730 122926
rect -4886 118586 588810 119206
rect -2966 114866 586890 115486
rect -8726 112026 592650 112646
rect -6806 108306 590730 108926
rect -4886 104586 588810 105206
rect -2966 100866 586890 101486
rect -8726 98026 592650 98646
rect -6806 94306 590730 94926
rect -4886 90586 588810 91206
rect -2966 86866 586890 87486
rect -8726 84026 592650 84646
rect -6806 80306 590730 80926
rect -4886 76586 588810 77206
rect -2966 72866 586890 73486
rect -8726 70026 592650 70646
rect -6806 66306 590730 66926
rect -4886 62586 588810 63206
rect -2966 58866 586890 59486
rect -8726 56026 592650 56646
rect -6806 52306 590730 52926
rect -4886 48586 588810 49206
rect -2966 44866 586890 45486
rect -8726 42026 592650 42646
rect -6806 38306 590730 38926
rect -4886 34586 588810 35206
rect -2966 30866 586890 31486
rect -8726 28026 592650 28646
rect -6806 24306 590730 24926
rect -4886 20586 588810 21206
rect -2966 16866 586890 17486
rect -8726 14026 592650 14646
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 30866 586890 31486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 58866 586890 59486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 86866 586890 87486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 114866 586890 115486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 142866 586890 143486 6 vccd1
port 532 nsew power input
rlabel metal5 s 57794 155926 506414 156546 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 170866 586890 171486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 198866 586890 199486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 226866 586890 227486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 282866 586890 283486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 310866 586890 311486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 338866 586890 339486 6 vccd1
port 532 nsew power input
rlabel metal5 s 365794 351926 422414 352546 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 366866 586890 367486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 394866 586890 395486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 422866 586890 423486 6 vccd1
port 532 nsew power input
rlabel metal5 s 57794 437806 170414 438426 6 vccd1
port 532 nsew power input
rlabel metal5 s 197794 437806 310414 438426 6 vccd1
port 532 nsew power input
rlabel metal5 s 393794 437806 506414 438426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 450866 586890 451486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 478866 586890 479486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 534866 586890 535486 6 vccd1
port 532 nsew power input
rlabel metal5 s 57794 547926 506414 548546 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 562866 586890 563486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 590866 586890 591486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 618866 586890 619486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 646866 586890 647486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 674866 586890 675486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 57794 -1894 58414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 -1894 86414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 113794 -1894 114414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 -1894 142414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 -1894 170414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 197794 -1894 198414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 225794 -1894 226414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 -1894 282414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 309794 -1894 310414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 -1894 338414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 393794 -1894 394414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 -1894 422414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 449794 -1894 450414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 477794 -1894 478414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 57794 145308 58414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 145308 86414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 113794 145308 114414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 145308 142414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 145308 170414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 197794 145308 198414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 225794 145308 226414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 145308 254414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 145308 282414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 309794 145308 310414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 145308 338414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 393794 145308 394414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 145308 422414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 449794 145308 450414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 477794 145308 478414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 145308 506414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 197794 252308 198414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 225794 252308 226414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 252308 254414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 252308 282414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 309794 252308 310414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 365794 -1894 366414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 393794 252308 394414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 252308 422414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 477794 252308 478414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 252308 506414 275000 6 vccd1
port 532 nsew power input
rlabel metal4 s 57794 252308 58414 312000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 252308 86414 312000 6 vccd1
port 532 nsew power input
rlabel metal4 s 113794 252308 114414 312000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 252308 142414 312000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 252308 170414 312000 6 vccd1
port 532 nsew power input
rlabel metal4 s 365794 342099 366414 362000 6 vccd1
port 532 nsew power input
rlabel metal4 s 393794 342099 394414 362000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 342099 422414 362000 6 vccd1
port 532 nsew power input
rlabel metal4 s 449794 252308 450414 362000 6 vccd1
port 532 nsew power input
rlabel metal4 s 477794 329000 478414 362000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 329000 506414 362000 6 vccd1
port 532 nsew power input
rlabel metal4 s 57794 427033 58414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 427033 86414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 113794 427033 114414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 427033 142414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 427033 170414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 197794 426000 198414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 225794 426000 226414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 426000 254414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 426000 282414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 309794 426000 310414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 252308 338414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 393794 429099 394414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 429099 422414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 449794 429099 450414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 477794 429099 478414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 429099 506414 451000 6 vccd1
port 532 nsew power input
rlabel metal4 s 57794 538308 58414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 538308 86414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 113794 538308 114414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 538308 142414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 538308 170414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 197794 538308 198414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 225794 538308 226414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 538308 254414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 538308 282414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 309794 538308 310414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 538308 338414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 393794 538308 394414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 538308 422414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 449794 538308 450414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 477794 538308 478414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 538308 506414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 29794 -1894 30414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 57794 645308 58414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 85794 645308 86414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 113794 645308 114414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 645308 142414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 169794 645308 170414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 197794 645308 198414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 225794 645308 226414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 645308 254414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 645308 282414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 309794 645308 310414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 337794 645308 338414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 365794 429099 366414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 393794 645308 394414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 645308 422414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 449794 645308 450414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 477794 645308 478414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 645308 506414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 533794 -1894 534414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 561794 -1894 562414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 34586 588810 35206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 62586 588810 63206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 90586 588810 91206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 118586 588810 119206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 146586 588810 147206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 174586 588810 175206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 202586 588810 203206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 230586 588810 231206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 286586 588810 287206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 314586 588810 315206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 342586 588810 343206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 370586 588810 371206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 398586 588810 399206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 426586 588810 427206 6 vccd2
port 533 nsew power input
rlabel metal5 s 61514 439646 146134 440266 6 vccd2
port 533 nsew power input
rlabel metal5 s 397514 439646 510134 440266 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 454586 588810 455206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 482586 588810 483206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 538586 588810 539206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 566586 588810 567206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 594586 588810 595206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 622586 588810 623206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 650586 588810 651206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 678586 588810 679206 6 vccd2
port 533 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 61514 -3814 62134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 -3814 90134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 117514 -3814 118134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 -3814 146134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 -3814 174134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 229514 -3814 230134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 -3814 286134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 313514 -3814 314134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 -3814 342134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 397514 -3814 398134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 -3814 426134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 453514 -3814 454134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 481514 -3814 482134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 61514 145308 62134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 145308 90134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 117514 145308 118134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 145308 146134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 145308 174134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 229514 145308 230134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 145308 258134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 145308 286134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 313514 145308 314134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 145308 342134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 397514 145308 398134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 145308 426134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 453514 145308 454134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 481514 145308 482134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 145308 510134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 201514 -3814 202134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 229514 252308 230134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 252308 258134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 252308 286134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 313514 252308 314134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 369514 -3814 370134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 397514 252308 398134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 481514 252308 482134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 252308 510134 275000 6 vccd2
port 533 nsew power input
rlabel metal4 s 61514 252308 62134 312000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 252308 90134 312000 6 vccd2
port 533 nsew power input
rlabel metal4 s 117514 252308 118134 312000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 252308 146134 312000 6 vccd2
port 533 nsew power input
rlabel metal4 s 369514 342099 370134 362000 6 vccd2
port 533 nsew power input
rlabel metal4 s 397514 342099 398134 362000 6 vccd2
port 533 nsew power input
rlabel metal4 s 453514 252308 454134 362000 6 vccd2
port 533 nsew power input
rlabel metal4 s 481514 329000 482134 362000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 329000 510134 362000 6 vccd2
port 533 nsew power input
rlabel metal4 s 61514 427033 62134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 427033 90134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 117514 427033 118134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 427033 146134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 252308 174134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 229514 426000 230134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 426000 258134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 426000 286134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 313514 426000 314134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 252308 342134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 397514 429099 398134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 252308 426134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 453514 429099 454134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 481514 429099 482134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 429099 510134 451000 6 vccd2
port 533 nsew power input
rlabel metal4 s 61514 538308 62134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 538308 90134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 117514 538308 118134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 538308 146134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 538308 174134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 229514 538308 230134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 538308 258134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 538308 286134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 313514 538308 314134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 538308 342134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 397514 538308 398134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 538308 426134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 453514 538308 454134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 481514 538308 482134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 538308 510134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 33514 -3814 34134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 61514 645308 62134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 89514 645308 90134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 117514 645308 118134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 645308 146134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 173514 645308 174134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 201514 426000 202134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 229514 645308 230134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 645308 258134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 645308 286134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 313514 645308 314134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 341514 645308 342134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 369514 429099 370134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 397514 645308 398134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 645308 426134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 453514 645308 454134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 481514 645308 482134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 645308 510134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 537514 -3814 538134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 565514 -3814 566134 707750 6 vccd2
port 533 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 38306 590730 38926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 66306 590730 66926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 94306 590730 94926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 122306 590730 122926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 150306 590730 150926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 178306 590730 178926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 206306 590730 206926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 234306 590730 234926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 290306 590730 290926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 318306 590730 318926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 346306 590730 346926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 374306 590730 374926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 402306 590730 402926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 430306 590730 430926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 458306 590730 458926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 486306 590730 486926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 542306 590730 542926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 570306 590730 570926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 598306 590730 598926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 626306 590730 626926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 654306 590730 654926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 682306 590730 682926 6 vdda1
port 534 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 65234 -5734 65854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 -5734 93854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 121234 -5734 121854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 -5734 149854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 -5734 177854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 233234 -5734 233854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 -5734 289854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 317234 -5734 317854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 -5734 345854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 401234 -5734 401854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 -5734 429854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 457234 -5734 457854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 485234 -5734 485854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 65234 145308 65854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 145308 93854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 121234 145308 121854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 145308 149854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 145308 177854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 233234 145308 233854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 145308 261854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 145308 289854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 317234 145308 317854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 145308 345854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 401234 145308 401854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 145308 429854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 457234 145308 457854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 485234 145308 485854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 145308 513854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 205234 -5734 205854 275000 6 vdda1
port 534 nsew power input
rlabel metal4 s 233234 252308 233854 275000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 252308 261854 275000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 252308 289854 275000 6 vdda1
port 534 nsew power input
rlabel metal4 s 317234 252308 317854 275000 6 vdda1
port 534 nsew power input
rlabel metal4 s 373234 -5734 373854 275000 6 vdda1
port 534 nsew power input
rlabel metal4 s 401234 252308 401854 275000 6 vdda1
port 534 nsew power input
rlabel metal4 s 485234 252308 485854 275000 6 vdda1
port 534 nsew power input
rlabel metal4 s 65234 252308 65854 312000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 252308 93854 312000 6 vdda1
port 534 nsew power input
rlabel metal4 s 121234 252308 121854 312000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 252308 149854 312000 6 vdda1
port 534 nsew power input
rlabel metal4 s 373234 342099 373854 362000 6 vdda1
port 534 nsew power input
rlabel metal4 s 401234 342099 401854 362000 6 vdda1
port 534 nsew power input
rlabel metal4 s 457234 252308 457854 362000 6 vdda1
port 534 nsew power input
rlabel metal4 s 485234 329000 485854 362000 6 vdda1
port 534 nsew power input
rlabel metal4 s 65234 427033 65854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 427033 93854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 121234 427033 121854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 427033 149854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 252308 177854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 233234 426000 233854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 426000 261854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 426000 289854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 317234 426000 317854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 252308 345854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 401234 429099 401854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 252308 429854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 457234 429099 457854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 485234 429099 485854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 252308 513854 451000 6 vdda1
port 534 nsew power input
rlabel metal4 s 65234 538308 65854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 538308 93854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 121234 538308 121854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 538308 149854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 538308 177854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 233234 538308 233854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 538308 261854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 538308 289854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 317234 538308 317854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 538308 345854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 401234 538308 401854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 538308 429854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 457234 538308 457854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 485234 538308 485854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 538308 513854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 37234 -5734 37854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 65234 645308 65854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 93234 645308 93854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 121234 645308 121854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 645308 149854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 177234 645308 177854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 205234 426000 205854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 233234 645308 233854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 645308 261854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 645308 289854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 317234 645308 317854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 345234 645308 345854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 373234 429099 373854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 401234 645308 401854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 645308 429854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 457234 645308 457854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 485234 645308 485854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 645308 513854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 541234 -5734 541854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 569234 -5734 569854 709670 6 vdda1
port 534 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 42026 592650 42646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 70026 592650 70646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 98026 592650 98646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 126026 592650 126646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 154026 592650 154646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 182026 592650 182646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 210026 592650 210646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 238026 592650 238646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 294026 592650 294646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 322026 592650 322646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 350026 592650 350646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 378026 592650 378646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 406026 592650 406646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 434026 592650 434646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 462026 592650 462646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 490026 592650 490646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 546026 592650 546646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 574026 592650 574646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 602026 592650 602646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 630026 592650 630646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 658026 592650 658646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 686026 592650 686646 6 vdda2
port 535 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 68954 -7654 69574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 -7654 97574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 124954 -7654 125574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 -7654 153574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 -7654 181574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 236954 -7654 237574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 -7654 293574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 320954 -7654 321574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 -7654 349574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 404954 -7654 405574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 -7654 433574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 460954 -7654 461574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 488954 -7654 489574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 68954 145308 69574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 145308 97574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 124954 145308 125574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 145308 153574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 145308 181574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 236954 145308 237574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 145308 265574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 145308 293574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 320954 145308 321574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 145308 349574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 404954 145308 405574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 145308 433574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 460954 145308 461574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 488954 145308 489574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 145308 517574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 208954 -7654 209574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 236954 252308 237574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 252308 265574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 252308 293574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 320954 252308 321574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 376954 -7654 377574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 404954 252308 405574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 460954 252308 461574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 488954 252308 489574 275000 6 vdda2
port 535 nsew power input
rlabel metal4 s 68954 252308 69574 312000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 252308 97574 312000 6 vdda2
port 535 nsew power input
rlabel metal4 s 124954 252308 125574 312000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 252308 153574 312000 6 vdda2
port 535 nsew power input
rlabel metal4 s 376954 342099 377574 362000 6 vdda2
port 535 nsew power input
rlabel metal4 s 404954 342099 405574 362000 6 vdda2
port 535 nsew power input
rlabel metal4 s 460954 329000 461574 362000 6 vdda2
port 535 nsew power input
rlabel metal4 s 488954 329000 489574 362000 6 vdda2
port 535 nsew power input
rlabel metal4 s 68954 427033 69574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 427033 97574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 124954 427033 125574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 427033 153574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 252308 181574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 236954 426000 237574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 426000 265574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 426000 293574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 320954 426000 321574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 252308 349574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 404954 429099 405574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 252308 433574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 460954 429099 461574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 488954 429099 489574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 252308 517574 451000 6 vdda2
port 535 nsew power input
rlabel metal4 s 68954 538308 69574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 538308 97574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 124954 538308 125574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 538308 153574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 538308 181574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 236954 538308 237574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 538308 265574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 538308 293574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 320954 538308 321574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 538308 349574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 404954 538308 405574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 538308 433574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 460954 538308 461574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 488954 538308 489574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 538308 517574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 40954 -7654 41574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 68954 645308 69574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 96954 645308 97574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 124954 645308 125574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 645308 153574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 180954 645308 181574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 208954 426000 209574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 236954 645308 237574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 645308 265574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 645308 293574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 320954 645308 321574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 348954 645308 349574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 376954 429099 377574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 404954 645308 405574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 645308 433574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 460954 645308 461574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 488954 645308 489574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 645308 517574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 544954 -7654 545574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 572954 -7654 573574 711590 6 vdda2
port 535 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 24306 590730 24926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 52306 590730 52926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 80306 590730 80926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 108306 590730 108926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 164306 590730 164926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 192306 590730 192926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 220306 590730 220926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 248306 590730 248926 6 vssa1
port 536 nsew ground input
rlabel metal5 s 219234 263246 303854 263866 6 vssa1
port 536 nsew ground input
rlabel metal5 s 387234 263246 499854 263866 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 276306 590730 276926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 304306 590730 304926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 332306 590730 332926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 360306 590730 360926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 416306 590730 416926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 444306 590730 444926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 472306 590730 472926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 500306 590730 500926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 528306 590730 528926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 556306 590730 556926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 584306 590730 584926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 612306 590730 612926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 668306 590730 668926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 696306 590730 696926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 -5734 79854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 107234 -5734 107854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 163234 -5734 163854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 191234 -5734 191854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 -5734 219854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 247234 -5734 247854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 275234 -5734 275854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 303234 -5734 303854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 331234 -5734 331854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 415234 -5734 415854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 443234 -5734 443854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 471234 -5734 471854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 -5734 499854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 145308 79854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 107234 145308 107854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 145308 135854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 163234 145308 163854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 191234 145308 191854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 145308 219854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 247234 145308 247854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 275234 145308 275854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 303234 145308 303854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 331234 145308 331854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 145308 387854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 415234 145308 415854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 443234 145308 443854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 471234 145308 471854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 145308 499854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 252308 219854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 247234 252308 247854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 275234 252308 275854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 303234 252308 303854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 359234 -5734 359854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 252308 387854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 415234 252308 415854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 471234 252308 471854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 252308 499854 275000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 252308 79854 312000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 107234 252308 107854 312000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 252308 135854 312000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 163234 252308 163854 312000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 359234 342099 359854 362000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 342099 387854 362000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 415234 342099 415854 362000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 471234 329000 471854 362000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 329000 499854 362000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 427033 79854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 107234 427033 107854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 427033 135854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 163234 427033 163854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 191234 252308 191854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 426000 219854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 247234 426000 247854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 275234 426000 275854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 303234 426000 303854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 331234 252308 331854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 429099 387854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 415234 429099 415854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 443234 252308 443854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 471234 429099 471854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 429099 499854 451000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 538308 79854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 107234 538308 107854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 538308 135854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 163234 538308 163854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 191234 538308 191854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 538308 219854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 247234 538308 247854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 275234 538308 275854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 303234 538308 303854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 331234 538308 331854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 538308 387854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 415234 538308 415854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 443234 538308 443854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 471234 538308 471854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 538308 499854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground input
rlabel metal4 s 23234 -5734 23854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 51234 -5734 51854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 645308 79854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 107234 645308 107854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 645308 135854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 163234 645308 163854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 191234 645308 191854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 645308 219854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 247234 645308 247854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 275234 645308 275854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 303234 645308 303854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 331234 645308 331854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 359234 429099 359854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 645308 387854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 415234 645308 415854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 443234 645308 443854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 471234 645308 471854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 645308 499854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 527234 -5734 527854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 555234 -5734 555854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 28026 592650 28646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 56026 592650 56646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 84026 592650 84646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 112026 592650 112646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 537 nsew ground input
rlabel metal5 s 82954 154966 503574 155586 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 168026 592650 168646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 196026 592650 196646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 224026 592650 224646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 252026 592650 252646 6 vssa2
port 537 nsew ground input
rlabel metal5 s 222954 265086 307574 265706 6 vssa2
port 537 nsew ground input
rlabel metal5 s 390954 265086 503574 265706 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 280026 592650 280646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 308026 592650 308646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 336026 592650 336646 6 vssa2
port 537 nsew ground input
rlabel metal5 s 362954 350966 419574 351586 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 364026 592650 364646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 420026 592650 420646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 448026 592650 448646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 476026 592650 476646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 504026 592650 504646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 532026 592650 532646 6 vssa2
port 537 nsew ground input
rlabel metal5 s 82954 546966 503574 547586 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 560026 592650 560646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 588026 592650 588646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 616026 592650 616646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 672026 592650 672646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 700026 592650 700646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 -7654 83574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 110954 -7654 111574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 166954 -7654 167574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 194954 -7654 195574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 -7654 223574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 250954 -7654 251574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 278954 -7654 279574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 306954 -7654 307574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 334954 -7654 335574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 418954 -7654 419574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 446954 -7654 447574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 474954 -7654 475574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 -7654 503574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 145308 83574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 110954 145308 111574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 145308 139574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 166954 145308 167574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 194954 145308 195574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 145308 223574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 250954 145308 251574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 278954 145308 279574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 306954 145308 307574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 334954 145308 335574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 145308 391574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 418954 145308 419574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 446954 145308 447574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 474954 145308 475574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 145308 503574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 252308 223574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 250954 252308 251574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 278954 252308 279574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 306954 252308 307574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 362954 -7654 363574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 252308 391574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 418954 252308 419574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 474954 252308 475574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 252308 503574 275000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 252308 83574 312000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 110954 252308 111574 312000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 252308 139574 312000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 166954 252308 167574 312000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 362954 342099 363574 362000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 342099 391574 362000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 418954 342099 419574 362000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 474954 329000 475574 362000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 329000 503574 362000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 427033 83574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 110954 427033 111574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 427033 139574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 166954 427033 167574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 194954 252308 195574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 426000 223574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 250954 426000 251574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 278954 426000 279574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 306954 426000 307574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 334954 252308 335574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 429099 391574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 418954 429099 419574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 446954 252308 447574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 474954 429099 475574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 429099 503574 451000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 538308 83574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 110954 538308 111574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 538308 139574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 166954 538308 167574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 194954 538308 195574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 538308 223574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 250954 538308 251574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 278954 538308 279574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 306954 538308 307574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 334954 538308 335574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 538308 391574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 418954 538308 419574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 446954 538308 447574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 474954 538308 475574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 538308 503574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground input
rlabel metal4 s 26954 -7654 27574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 54954 -7654 55574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 645308 83574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 110954 645308 111574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 645308 139574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 166954 645308 167574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 194954 645308 195574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 645308 223574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 250954 645308 251574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 278954 645308 279574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 306954 645308 307574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 334954 645308 335574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 362954 429099 363574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 645308 391574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 418954 645308 419574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 446954 645308 447574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 474954 645308 475574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 645308 503574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 530954 -7654 531574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 558954 -7654 559574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 16866 586890 17486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 44866 586890 45486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 72866 586890 73486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 100866 586890 101486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 156866 586890 157486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 184866 586890 185486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 212866 586890 213486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 240866 586890 241486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 268866 586890 269486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 296866 586890 297486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 324866 586890 325486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 352866 586890 353486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 408866 586890 409486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 436866 586890 437486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 464866 586890 465486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 492866 586890 493486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 520866 586890 521486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 548866 586890 549486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 576866 586890 577486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 604866 586890 605486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 660866 586890 661486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 688866 586890 689486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 -1894 72414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99794 -1894 100414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 155794 -1894 156414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 183794 -1894 184414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 239794 -1894 240414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 267794 -1894 268414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 295794 -1894 296414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 323794 -1894 324414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 -1894 352414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 407794 -1894 408414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 435794 -1894 436414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 463794 -1894 464414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 -1894 492414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 145308 72414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99794 145308 100414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 145308 128414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 155794 145308 156414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 183794 145308 184414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 239794 145308 240414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 267794 145308 268414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 295794 145308 296414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 323794 145308 324414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 145308 352414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 145308 380414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 407794 145308 408414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 435794 145308 436414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 463794 145308 464414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 145308 492414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211794 -1894 212414 275000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 239794 252308 240414 275000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 267794 252308 268414 275000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 295794 252308 296414 275000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 252308 380414 275000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 407794 252308 408414 275000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 463794 252308 464414 275000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 252308 492414 275000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 252308 72414 312000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99794 252308 100414 312000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 252308 128414 312000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 155794 252308 156414 312000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 342099 380414 362000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 407794 342099 408414 362000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 463794 329000 464414 362000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 329000 492414 362000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 427033 72414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99794 427033 100414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 427033 128414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 155794 427033 156414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 183794 252308 184414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 239794 426000 240414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 267794 426000 268414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 295794 426000 296414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 323794 252308 324414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 252308 352414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 429099 380414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 407794 429099 408414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 435794 252308 436414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 463794 429099 464414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 429099 492414 451000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 538308 72414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99794 538308 100414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 538308 128414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 155794 538308 156414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 183794 538308 184414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 239794 538308 240414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 267794 538308 268414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 295794 538308 296414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 323794 538308 324414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 538308 352414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 538308 380414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 407794 538308 408414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 435794 538308 436414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 463794 538308 464414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 538308 492414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground input
rlabel metal4 s 15794 -1894 16414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 43794 -1894 44414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 645308 72414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99794 645308 100414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 645308 128414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 155794 645308 156414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 183794 645308 184414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211794 426000 212414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 239794 645308 240414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 267794 645308 268414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 295794 645308 296414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 323794 645308 324414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 645308 352414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 645308 380414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 407794 645308 408414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 435794 645308 436414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 463794 645308 464414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 645308 492414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 519794 -1894 520414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 547794 -1894 548414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 575794 -1894 576414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 20586 588810 21206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 48586 588810 49206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 76586 588810 77206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 104586 588810 105206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 160586 588810 161206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 188586 588810 189206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 216586 588810 217206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 244586 588810 245206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 272586 588810 273206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 300586 588810 301206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 328586 588810 329206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 356586 588810 357206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 412586 588810 413206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 440586 588810 441206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 468586 588810 469206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 496586 588810 497206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 524586 588810 525206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 552586 588810 553206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 580586 588810 581206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 608586 588810 609206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 664586 588810 665206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 692586 588810 693206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 -3814 76134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 103514 -3814 104134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 159514 -3814 160134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 187514 -3814 188134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 243514 -3814 244134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 271514 -3814 272134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 299514 -3814 300134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 327514 -3814 328134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 -3814 356134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 411514 -3814 412134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 439514 -3814 440134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 467514 -3814 468134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 -3814 496134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 145308 76134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 103514 145308 104134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 145308 132134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 159514 145308 160134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 187514 145308 188134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 243514 145308 244134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 271514 145308 272134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 299514 145308 300134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 327514 145308 328134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 145308 356134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 145308 384134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 411514 145308 412134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 439514 145308 440134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 467514 145308 468134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 145308 496134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215514 -3814 216134 275000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 243514 252308 244134 275000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 271514 252308 272134 275000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 299514 252308 300134 275000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 252308 384134 275000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 411514 252308 412134 275000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 467514 252308 468134 275000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 252308 496134 275000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 252308 76134 312000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 103514 252308 104134 312000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 252308 132134 312000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 159514 252308 160134 312000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 342099 384134 362000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 411514 342099 412134 362000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 467514 329000 468134 362000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 329000 496134 362000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 427033 76134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 103514 427033 104134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 427033 132134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 159514 427033 160134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 187514 252308 188134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 243514 426000 244134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 271514 426000 272134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 299514 426000 300134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 327514 252308 328134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 252308 356134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 429099 384134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 411514 429099 412134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 439514 252308 440134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 467514 429099 468134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 429099 496134 451000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 538308 76134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 103514 538308 104134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 538308 132134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 159514 538308 160134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 187514 538308 188134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 243514 538308 244134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 271514 538308 272134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 299514 538308 300134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 327514 538308 328134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 538308 356134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 538308 384134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 411514 538308 412134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 439514 538308 440134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 467514 538308 468134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 538308 496134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground input
rlabel metal4 s 19514 -3814 20134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 47514 -3814 48134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 645308 76134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 103514 645308 104134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 645308 132134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 159514 645308 160134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 187514 645308 188134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215514 426000 216134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 243514 645308 244134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 271514 645308 272134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 299514 645308 300134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 327514 645308 328134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 645308 356134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 645308 384134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 411514 645308 412134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 439514 645308 440134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 467514 645308 468134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 645308 496134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 523514 -3814 524134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 551514 -3814 552134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 579514 -3814 580134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 93398180
string GDS_FILE /home/burak/asic_tools/caravel_vscpu3x/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 89537968
<< end >>

