magic
tech sky130A
magscale 1 2
timestamp 1655291147
<< metal1 >>
rect 38378 700952 38384 701004
rect 38436 700992 38442 701004
rect 99834 700992 99840 701004
rect 38436 700964 99840 700992
rect 38436 700952 38442 700964
rect 99834 700952 99840 700964
rect 99892 700992 99898 701004
rect 161290 700992 161296 701004
rect 99892 700964 161296 700992
rect 99892 700952 99898 700964
rect 161290 700952 161296 700964
rect 161348 700992 161354 701004
rect 222746 700992 222752 701004
rect 161348 700964 222752 700992
rect 161348 700952 161354 700964
rect 222746 700952 222752 700964
rect 222804 700992 222810 701004
rect 284202 700992 284208 701004
rect 222804 700964 284208 700992
rect 222804 700952 222810 700964
rect 284202 700952 284208 700964
rect 284260 700992 284266 701004
rect 345750 700992 345756 701004
rect 284260 700964 345756 700992
rect 284260 700952 284266 700964
rect 345750 700952 345756 700964
rect 345808 700992 345814 701004
rect 407206 700992 407212 701004
rect 345808 700964 407212 700992
rect 345808 700952 345814 700964
rect 407206 700952 407212 700964
rect 407264 700992 407270 701004
rect 468662 700992 468668 701004
rect 407264 700964 468668 700992
rect 407264 700952 407270 700964
rect 468662 700952 468668 700964
rect 468720 700992 468726 701004
rect 530118 700992 530124 701004
rect 468720 700964 530124 700992
rect 468720 700952 468726 700964
rect 530118 700952 530124 700964
rect 530176 700992 530182 701004
rect 531222 700992 531228 701004
rect 530176 700964 531228 700992
rect 530176 700952 530182 700964
rect 531222 700952 531228 700964
rect 531280 700952 531286 701004
rect 253474 700340 253480 700392
rect 253532 700380 253538 700392
rect 305638 700380 305644 700392
rect 253532 700352 305644 700380
rect 253532 700340 253538 700352
rect 305638 700340 305644 700352
rect 305696 700340 305702 700392
rect 69106 700272 69112 700324
rect 69164 700312 69170 700324
rect 304258 700312 304264 700324
rect 69164 700284 304264 700312
rect 69164 700272 69170 700284
rect 304258 700272 304264 700284
rect 304316 700272 304322 700324
rect 531222 700272 531228 700324
rect 531280 700312 531286 700324
rect 580258 700312 580264 700324
rect 531280 700284 580264 700312
rect 531280 700272 531286 700284
rect 580258 700272 580264 700284
rect 580316 700272 580322 700324
rect 37918 699660 37924 699712
rect 37976 699700 37982 699712
rect 38378 699700 38384 699712
rect 37976 699672 38384 699700
rect 37976 699660 37982 699672
rect 38378 699660 38384 699672
rect 38436 699660 38442 699712
rect 436738 699660 436744 699712
rect 436796 699700 436802 699712
rect 437934 699700 437940 699712
rect 436796 699672 437940 699700
rect 436796 699660 436802 699672
rect 437934 699660 437940 699672
rect 437992 699660 437998 699712
rect 315022 698912 315028 698964
rect 315080 698952 315086 698964
rect 400214 698952 400220 698964
rect 315080 698924 400220 698952
rect 315080 698912 315086 698924
rect 400214 698912 400220 698924
rect 400272 698912 400278 698964
rect 59262 697552 59268 697604
rect 59320 697592 59326 697604
rect 545482 697592 545488 697604
rect 59320 697564 545488 697592
rect 59320 697552 59326 697564
rect 545482 697552 545488 697564
rect 545540 697552 545546 697604
rect 3418 684496 3424 684548
rect 3476 684536 3482 684548
rect 316678 684536 316684 684548
rect 3476 684508 316684 684536
rect 3476 684496 3482 684508
rect 316678 684496 316684 684508
rect 316736 684496 316742 684548
rect 2774 660288 2780 660340
rect 2832 660328 2838 660340
rect 37918 660328 37924 660340
rect 2832 660300 37924 660328
rect 2832 660288 2838 660300
rect 37918 660288 37924 660300
rect 37976 660288 37982 660340
rect 137554 658248 137560 658300
rect 137612 658288 137618 658300
rect 579890 658288 579896 658300
rect 137612 658260 579896 658288
rect 137612 658248 137618 658260
rect 579890 658248 579896 658260
rect 579948 658248 579954 658300
rect 318794 651992 318800 652044
rect 318852 652032 318858 652044
rect 498194 652032 498200 652044
rect 318852 652004 498200 652032
rect 318852 651992 318858 652004
rect 498194 651992 498200 652004
rect 498252 651992 498258 652044
rect 129734 650632 129740 650684
rect 129792 650672 129798 650684
rect 429286 650672 429292 650684
rect 129792 650644 429292 650672
rect 129792 650632 129798 650644
rect 429286 650632 429292 650644
rect 429344 650632 429350 650684
rect 291194 650020 291200 650072
rect 291252 650060 291258 650072
rect 457438 650060 457444 650072
rect 291252 650032 457444 650060
rect 291252 650020 291258 650032
rect 457438 650020 457444 650032
rect 457496 650020 457502 650072
rect 191834 649272 191840 649324
rect 191892 649312 191898 649324
rect 430574 649312 430580 649324
rect 191892 649284 430580 649312
rect 191892 649272 191898 649284
rect 430574 649272 430580 649284
rect 430632 649272 430638 649324
rect 280982 648728 280988 648780
rect 281040 648768 281046 648780
rect 430666 648768 430672 648780
rect 281040 648740 430672 648768
rect 281040 648728 281046 648740
rect 430666 648728 430672 648740
rect 430724 648728 430730 648780
rect 289814 648660 289820 648712
rect 289872 648700 289878 648712
rect 489914 648700 489920 648712
rect 289872 648672 489920 648700
rect 289872 648660 289878 648672
rect 489914 648660 489920 648672
rect 489972 648660 489978 648712
rect 217778 648592 217784 648644
rect 217836 648632 217842 648644
rect 580258 648632 580264 648644
rect 217836 648604 580264 648632
rect 217836 648592 217842 648604
rect 580258 648592 580264 648604
rect 580316 648592 580322 648644
rect 318242 648116 318248 648168
rect 318300 648156 318306 648168
rect 427814 648156 427820 648168
rect 318300 648128 427820 648156
rect 318300 648116 318306 648128
rect 427814 648116 427820 648128
rect 427872 648116 427878 648168
rect 312538 648048 312544 648100
rect 312596 648088 312602 648100
rect 332594 648088 332600 648100
rect 312596 648060 332600 648088
rect 312596 648048 312602 648060
rect 332594 648048 332600 648060
rect 332652 648048 332658 648100
rect 298738 647980 298744 648032
rect 298796 648020 298802 648032
rect 378318 648020 378324 648032
rect 298796 647992 378324 648020
rect 298796 647980 298802 647992
rect 378318 647980 378324 647992
rect 378376 647980 378382 648032
rect 319714 647912 319720 647964
rect 319772 647952 319778 647964
rect 355134 647952 355140 647964
rect 319772 647924 355140 647952
rect 319772 647912 319778 647924
rect 355134 647912 355140 647924
rect 355192 647912 355198 647964
rect 313918 647844 313924 647896
rect 313976 647884 313982 647896
rect 359550 647884 359556 647896
rect 313976 647856 359556 647884
rect 313976 647844 313982 647856
rect 359550 647844 359556 647856
rect 359608 647844 359614 647896
rect 375374 647844 375380 647896
rect 375432 647884 375438 647896
rect 423858 647884 423864 647896
rect 375432 647856 423864 647884
rect 375432 647844 375438 647856
rect 423858 647844 423864 647856
rect 423916 647844 423922 647896
rect 316862 647776 316868 647828
rect 316920 647816 316926 647828
rect 364334 647816 364340 647828
rect 316920 647788 364340 647816
rect 316920 647776 316926 647788
rect 364334 647776 364340 647788
rect 364392 647776 364398 647828
rect 319806 647708 319812 647760
rect 319864 647748 319870 647760
rect 373166 647748 373172 647760
rect 319864 647720 373172 647748
rect 319864 647708 319870 647720
rect 373166 647708 373172 647720
rect 373224 647708 373230 647760
rect 315298 647640 315304 647692
rect 315356 647680 315362 647692
rect 368566 647680 368572 647692
rect 315356 647652 368572 647680
rect 315356 647640 315362 647652
rect 368566 647640 368572 647652
rect 368624 647640 368630 647692
rect 284938 647572 284944 647624
rect 284996 647612 285002 647624
rect 350534 647612 350540 647624
rect 284996 647584 350540 647612
rect 284996 647572 285002 647584
rect 350534 647572 350540 647584
rect 350592 647572 350598 647624
rect 314010 647504 314016 647556
rect 314068 647544 314074 647556
rect 382734 647544 382740 647556
rect 314068 647516 382740 647544
rect 314068 647504 314074 647516
rect 382734 647504 382740 647516
rect 382792 647504 382798 647556
rect 318150 647436 318156 647488
rect 318208 647476 318214 647488
rect 387334 647476 387340 647488
rect 318208 647448 387340 647476
rect 318208 647436 318214 647448
rect 387334 647436 387340 647448
rect 387392 647436 387398 647488
rect 316770 647368 316776 647420
rect 316828 647408 316834 647420
rect 396350 647408 396356 647420
rect 316828 647380 396356 647408
rect 316828 647368 316834 647380
rect 396350 647368 396356 647380
rect 396408 647368 396414 647420
rect 318058 647300 318064 647352
rect 318116 647340 318122 647352
rect 337102 647340 337108 647352
rect 318116 647312 337108 647340
rect 318116 647300 318122 647312
rect 337102 647300 337108 647312
rect 337160 647300 337166 647352
rect 319622 647232 319628 647284
rect 319680 647272 319686 647284
rect 323486 647272 323492 647284
rect 319680 647244 323492 647272
rect 319680 647232 319686 647244
rect 323486 647232 323492 647244
rect 323544 647232 323550 647284
rect 280706 646620 280712 646672
rect 280764 646660 280770 646672
rect 341518 646660 341524 646672
rect 280764 646632 341524 646660
rect 280764 646620 280770 646632
rect 341518 646620 341524 646632
rect 341576 646620 341582 646672
rect 296714 646552 296720 646604
rect 296772 646592 296778 646604
rect 429930 646592 429936 646604
rect 296772 646564 429936 646592
rect 296772 646552 296778 646564
rect 429930 646552 429936 646564
rect 429988 646552 429994 646604
rect 298094 646484 298100 646536
rect 298152 646524 298158 646536
rect 432598 646524 432604 646536
rect 298152 646496 432604 646524
rect 298152 646484 298158 646496
rect 432598 646484 432604 646496
rect 432656 646484 432662 646536
rect 291286 646416 291292 646468
rect 291344 646456 291350 646468
rect 428458 646456 428464 646468
rect 291344 646428 428464 646456
rect 291344 646416 291350 646428
rect 428458 646416 428464 646428
rect 428516 646416 428522 646468
rect 288526 646348 288532 646400
rect 288584 646388 288590 646400
rect 429838 646388 429844 646400
rect 288584 646360 429844 646388
rect 288584 646348 288590 646360
rect 429838 646348 429844 646360
rect 429896 646348 429902 646400
rect 319438 646280 319444 646332
rect 319496 646320 319502 646332
rect 466730 646320 466736 646332
rect 319496 646292 466736 646320
rect 319496 646280 319502 646292
rect 466730 646280 466736 646292
rect 466788 646280 466794 646332
rect 282178 646212 282184 646264
rect 282236 646252 282242 646264
rect 430758 646252 430764 646264
rect 282236 646224 430764 646252
rect 282236 646212 282242 646224
rect 430758 646212 430764 646224
rect 430816 646212 430822 646264
rect 293954 646144 293960 646196
rect 294012 646184 294018 646196
rect 497642 646184 497648 646196
rect 294012 646156 497648 646184
rect 294012 646144 294018 646156
rect 497642 646144 497648 646156
rect 497700 646144 497706 646196
rect 296806 646076 296812 646128
rect 296864 646116 296870 646128
rect 511994 646116 512000 646128
rect 296864 646088 512000 646116
rect 296864 646076 296870 646088
rect 511994 646076 512000 646088
rect 512052 646076 512058 646128
rect 288434 646008 288440 646060
rect 288492 646048 288498 646060
rect 510614 646048 510620 646060
rect 288492 646020 510620 646048
rect 288492 646008 288498 646020
rect 510614 646008 510620 646020
rect 510672 646008 510678 646060
rect 40678 645940 40684 645992
rect 40736 645980 40742 645992
rect 409874 645980 409880 645992
rect 40736 645952 409880 645980
rect 40736 645940 40742 645952
rect 409874 645940 409880 645952
rect 409932 645940 409938 645992
rect 218698 645872 218704 645924
rect 218756 645912 218762 645924
rect 414382 645912 414388 645924
rect 218756 645884 414388 645912
rect 218756 645872 218762 645884
rect 414382 645872 414388 645884
rect 414440 645872 414446 645924
rect 302878 644444 302884 644496
rect 302936 644484 302942 644496
rect 317598 644484 317604 644496
rect 302936 644456 317604 644484
rect 302936 644444 302942 644456
rect 317598 644444 317604 644456
rect 317656 644444 317662 644496
rect 136542 640840 136548 640892
rect 136600 640880 136606 640892
rect 149054 640880 149060 640892
rect 136600 640852 149060 640880
rect 136600 640840 136606 640852
rect 149054 640840 149060 640852
rect 149112 640840 149118 640892
rect 134886 640772 134892 640824
rect 134944 640812 134950 640824
rect 140314 640812 140320 640824
rect 134944 640784 140320 640812
rect 134944 640772 134950 640784
rect 140314 640772 140320 640784
rect 140372 640772 140378 640824
rect 213914 640772 213920 640824
rect 213972 640812 213978 640824
rect 225782 640812 225788 640824
rect 213972 640784 225788 640812
rect 213972 640772 213978 640784
rect 225782 640772 225788 640784
rect 225840 640772 225846 640824
rect 100570 640704 100576 640756
rect 100628 640744 100634 640756
rect 124490 640744 124496 640756
rect 100628 640716 124496 640744
rect 100628 640704 100634 640716
rect 124490 640704 124496 640716
rect 124548 640704 124554 640756
rect 139854 640704 139860 640756
rect 139912 640744 139918 640756
rect 157426 640744 157432 640756
rect 139912 640716 157432 640744
rect 139912 640704 139918 640716
rect 157426 640704 157432 640716
rect 157484 640704 157490 640756
rect 212534 640704 212540 640756
rect 212592 640744 212598 640756
rect 272150 640744 272156 640756
rect 212592 640716 272156 640744
rect 212592 640704 212598 640716
rect 272150 640704 272156 640716
rect 272208 640704 272214 640756
rect 115382 640636 115388 640688
rect 115440 640676 115446 640688
rect 124582 640676 124588 640688
rect 115440 640648 124588 640676
rect 115440 640636 115446 640648
rect 124582 640636 124588 640648
rect 124640 640636 124646 640688
rect 137830 640636 137836 640688
rect 137888 640676 137894 640688
rect 160646 640676 160652 640688
rect 137888 640648 160652 640676
rect 137888 640636 137894 640648
rect 160646 640636 160652 640648
rect 160704 640636 160710 640688
rect 217870 640636 217876 640688
rect 217928 640676 217934 640688
rect 243170 640676 243176 640688
rect 217928 640648 243176 640676
rect 217928 640636 217934 640648
rect 243170 640636 243176 640648
rect 243228 640636 243234 640688
rect 56502 640568 56508 640620
rect 56560 640608 56566 640620
rect 77386 640608 77392 640620
rect 56560 640580 77392 640608
rect 56560 640568 56566 640580
rect 77386 640568 77392 640580
rect 77444 640568 77450 640620
rect 112162 640568 112168 640620
rect 112220 640608 112226 640620
rect 124674 640608 124680 640620
rect 112220 640580 124680 640608
rect 112220 640568 112226 640580
rect 124674 640568 124680 640580
rect 124732 640568 124738 640620
rect 134978 640568 134984 640620
rect 135036 640608 135042 640620
rect 140222 640608 140228 640620
rect 135036 640580 140228 640608
rect 135036 640568 135042 640580
rect 140222 640568 140228 640580
rect 140280 640568 140286 640620
rect 140314 640568 140320 640620
rect 140372 640608 140378 640620
rect 166442 640608 166448 640620
rect 140372 640580 166448 640608
rect 140372 640568 140378 640580
rect 166442 640568 166448 640580
rect 166500 640568 166506 640620
rect 218882 640568 218888 640620
rect 218940 640608 218946 640620
rect 252186 640608 252192 640620
rect 218940 640580 252192 640608
rect 218940 640568 218946 640580
rect 252186 640568 252192 640580
rect 252244 640568 252250 640620
rect 54938 640500 54944 640552
rect 54996 640540 55002 640552
rect 80606 640540 80612 640552
rect 54996 640512 80612 640540
rect 54996 640500 55002 640512
rect 80606 640500 80612 640512
rect 80664 640500 80670 640552
rect 109586 640500 109592 640552
rect 109644 640540 109650 640552
rect 122834 640540 122840 640552
rect 109644 640512 122840 640540
rect 109644 640500 109650 640512
rect 122834 640500 122840 640512
rect 122892 640500 122898 640552
rect 139210 640500 139216 640552
rect 139268 640540 139274 640552
rect 174814 640540 174820 640552
rect 139268 640512 174820 640540
rect 139268 640500 139274 640512
rect 174814 640500 174820 640512
rect 174872 640500 174878 640552
rect 189626 640500 189632 640552
rect 189684 640540 189690 640552
rect 205634 640540 205640 640552
rect 189684 640512 205640 640540
rect 189684 640500 189690 640512
rect 205634 640500 205640 640512
rect 205692 640500 205698 640552
rect 218790 640500 218796 640552
rect 218848 640540 218854 640552
rect 263778 640540 263784 640552
rect 218848 640512 263784 640540
rect 218848 640500 218854 640512
rect 263778 640500 263784 640512
rect 263836 640500 263842 640552
rect 54846 640432 54852 640484
rect 54904 640472 54910 640484
rect 88978 640472 88984 640484
rect 54904 640444 88984 640472
rect 54904 640432 54910 640444
rect 88978 640432 88984 640444
rect 89036 640432 89042 640484
rect 106366 640432 106372 640484
rect 106424 640472 106430 640484
rect 121454 640472 121460 640484
rect 106424 640444 121460 640472
rect 106424 640432 106430 640444
rect 121454 640432 121460 640444
rect 121512 640432 121518 640484
rect 137646 640432 137652 640484
rect 137704 640472 137710 640484
rect 140130 640472 140136 640484
rect 137704 640444 140136 640472
rect 137704 640432 137710 640444
rect 140130 640432 140136 640444
rect 140188 640432 140194 640484
rect 140222 640432 140228 640484
rect 140280 640472 140286 640484
rect 180610 640472 180616 640484
rect 140280 640444 180616 640472
rect 140280 640432 140286 640444
rect 180610 640432 180616 640444
rect 180668 640432 180674 640484
rect 214006 640432 214012 640484
rect 214064 640472 214070 640484
rect 269574 640472 269580 640484
rect 214064 640444 269580 640472
rect 214064 640432 214070 640444
rect 269574 640432 269580 640444
rect 269632 640432 269638 640484
rect 55122 640364 55128 640416
rect 55180 640404 55186 640416
rect 92198 640404 92204 640416
rect 55180 640376 92204 640404
rect 55180 640364 55186 640376
rect 92198 640364 92204 640376
rect 92256 640364 92262 640416
rect 103790 640364 103796 640416
rect 103848 640404 103854 640416
rect 120810 640404 120816 640416
rect 103848 640376 120816 640404
rect 103848 640364 103854 640376
rect 120810 640364 120816 640376
rect 120868 640364 120874 640416
rect 124214 640364 124220 640416
rect 124272 640404 124278 640416
rect 172238 640404 172244 640416
rect 124272 640376 172244 640404
rect 124272 640364 124278 640376
rect 172238 640364 172244 640376
rect 172296 640364 172302 640416
rect 192202 640364 192208 640416
rect 192260 640404 192266 640416
rect 204346 640404 204352 640416
rect 192260 640376 204352 640404
rect 192260 640364 192266 640376
rect 204346 640364 204352 640376
rect 204404 640364 204410 640416
rect 219342 640364 219348 640416
rect 219400 640404 219406 640416
rect 275370 640404 275376 640416
rect 219400 640376 275376 640404
rect 219400 640364 219406 640376
rect 275370 640364 275376 640376
rect 275428 640364 275434 640416
rect 55030 640296 55036 640348
rect 55088 640336 55094 640348
rect 94774 640336 94780 640348
rect 55088 640308 94780 640336
rect 55088 640296 55094 640308
rect 94774 640296 94780 640308
rect 94832 640296 94838 640348
rect 133874 640296 133880 640348
rect 133932 640336 133938 640348
rect 140038 640336 140044 640348
rect 133932 640308 140044 640336
rect 133932 640296 133938 640308
rect 140038 640296 140044 640308
rect 140096 640296 140102 640348
rect 140130 640296 140136 640348
rect 140188 640336 140194 640348
rect 186406 640336 186412 640348
rect 140188 640308 186412 640336
rect 140188 640296 140194 640308
rect 186406 640296 186412 640308
rect 186464 640296 186470 640348
rect 195422 640296 195428 640348
rect 195480 640336 195486 640348
rect 200850 640336 200856 640348
rect 195480 640308 200856 640336
rect 195480 640296 195486 640308
rect 200850 640296 200856 640308
rect 200908 640296 200914 640348
rect 217318 640296 217324 640348
rect 217376 640336 217382 640348
rect 231578 640336 231584 640348
rect 217376 640308 231584 640336
rect 217376 640296 217382 640308
rect 231578 640296 231584 640308
rect 231636 640296 231642 640348
rect 287698 640296 287704 640348
rect 287756 640336 287762 640348
rect 317690 640336 317696 640348
rect 287756 640308 317696 640336
rect 287756 640296 287762 640308
rect 317690 640296 317696 640308
rect 317748 640296 317754 640348
rect 215294 639208 215300 639260
rect 215352 639248 215358 639260
rect 234798 639248 234804 639260
rect 215352 639220 234804 639248
rect 215352 639208 215358 639220
rect 234798 639208 234804 639220
rect 234856 639208 234862 639260
rect 219618 639140 219624 639192
rect 219676 639180 219682 639192
rect 246390 639180 246396 639192
rect 219676 639152 246396 639180
rect 219676 639140 219682 639152
rect 246390 639140 246396 639152
rect 246448 639140 246454 639192
rect 210418 639072 210424 639124
rect 210476 639112 210482 639124
rect 237374 639112 237380 639124
rect 210476 639084 237380 639112
rect 210476 639072 210482 639084
rect 237374 639072 237380 639084
rect 237432 639072 237438 639124
rect 133138 639004 133144 639056
rect 133196 639044 133202 639056
rect 151630 639044 151636 639056
rect 133196 639016 151636 639044
rect 133196 639004 133202 639016
rect 151630 639004 151636 639016
rect 151688 639004 151694 639056
rect 206278 639004 206284 639056
rect 206336 639044 206342 639056
rect 254762 639044 254768 639056
rect 206336 639016 254768 639044
rect 206336 639004 206342 639016
rect 254762 639004 254768 639016
rect 254820 639004 254826 639056
rect 69014 638936 69020 638988
rect 69072 638976 69078 638988
rect 124306 638976 124312 638988
rect 69072 638948 124312 638976
rect 69072 638936 69078 638948
rect 124306 638936 124312 638948
rect 124364 638936 124370 638988
rect 135254 638936 135260 638988
rect 135312 638976 135318 638988
rect 183830 638976 183836 638988
rect 135312 638948 183836 638976
rect 135312 638936 135318 638948
rect 183830 638936 183836 638948
rect 183888 638936 183894 638988
rect 204254 638936 204260 638988
rect 204312 638976 204318 638988
rect 277946 638976 277952 638988
rect 204312 638948 277952 638976
rect 204312 638936 204318 638948
rect 277946 638936 277952 638948
rect 278004 638936 278010 638988
rect 223758 638188 223764 638240
rect 223816 638228 223822 638240
rect 223816 638200 229094 638228
rect 223816 638188 223822 638200
rect 215938 638120 215944 638172
rect 215996 638160 216002 638172
rect 215996 638132 228956 638160
rect 215996 638120 216002 638132
rect 217962 638052 217968 638104
rect 218020 638092 218026 638104
rect 228726 638092 228732 638104
rect 218020 638064 228732 638092
rect 218020 638052 218026 638064
rect 228726 638052 228732 638064
rect 228784 638052 228790 638104
rect 126238 637984 126244 638036
rect 126296 638024 126302 638036
rect 177850 638024 177856 638036
rect 126296 637996 177856 638024
rect 126296 637984 126302 637996
rect 177850 637984 177856 637996
rect 177908 637984 177914 638036
rect 204898 637984 204904 638036
rect 204956 638024 204962 638036
rect 223758 638024 223764 638036
rect 204956 637996 223764 638024
rect 204956 637984 204962 637996
rect 223758 637984 223764 637996
rect 223816 637984 223822 638036
rect 135162 637916 135168 637968
rect 135220 637956 135226 637968
rect 145558 637956 145564 637968
rect 135220 637928 145564 637956
rect 135220 637916 135226 637928
rect 145558 637916 145564 637928
rect 145616 637916 145622 637968
rect 213178 637916 213184 637968
rect 213236 637956 213242 637968
rect 222838 637956 222844 637968
rect 213236 637928 222844 637956
rect 213236 637916 213242 637928
rect 222838 637916 222844 637928
rect 222896 637916 222902 637968
rect 228928 637956 228956 638132
rect 229066 638024 229094 638200
rect 266262 638024 266268 638036
rect 229066 637996 266268 638024
rect 266262 637984 266268 637996
rect 266320 637984 266326 638036
rect 260190 637956 260196 637968
rect 228928 637928 260196 637956
rect 260190 637916 260196 637928
rect 260248 637916 260254 637968
rect 57790 637848 57796 637900
rect 57848 637888 57854 637900
rect 71222 637888 71228 637900
rect 57848 637860 71228 637888
rect 57848 637848 57854 637860
rect 71222 637848 71228 637860
rect 71280 637848 71286 637900
rect 136450 637848 136456 637900
rect 136508 637888 136514 637900
rect 154574 637888 154580 637900
rect 136508 637860 154580 637888
rect 136508 637848 136514 637860
rect 154574 637848 154580 637860
rect 154632 637848 154638 637900
rect 208394 637848 208400 637900
rect 208452 637888 208458 637900
rect 240318 637888 240324 637900
rect 208452 637860 240324 637888
rect 208452 637848 208458 637860
rect 240318 637848 240324 637860
rect 240376 637848 240382 637900
rect 56318 637780 56324 637832
rect 56376 637820 56382 637832
rect 65518 637820 65524 637832
rect 56376 637792 65524 637820
rect 56376 637780 56382 637792
rect 65518 637780 65524 637792
rect 65576 637780 65582 637832
rect 135070 637780 135076 637832
rect 135128 637820 135134 637832
rect 162854 637820 162860 637832
rect 135128 637792 162860 637820
rect 135128 637780 135134 637792
rect 162854 637780 162860 637792
rect 162912 637780 162918 637832
rect 206370 637780 206376 637832
rect 206428 637820 206434 637832
rect 248690 637820 248696 637832
rect 206428 637792 248696 637820
rect 206428 637780 206434 637792
rect 248690 637780 248696 637792
rect 248748 637780 248754 637832
rect 59354 637712 59360 637764
rect 59412 637752 59418 637764
rect 97902 637752 97908 637764
rect 59412 637724 97908 637752
rect 59412 637712 59418 637724
rect 97902 637712 97908 637724
rect 97960 637712 97966 637764
rect 124398 637752 124404 637764
rect 103486 637724 124404 637752
rect 56410 637644 56416 637696
rect 56468 637684 56474 637696
rect 62942 637684 62948 637696
rect 56468 637656 62948 637684
rect 56468 637644 56474 637656
rect 62942 637644 62948 637656
rect 63000 637644 63006 637696
rect 86770 637644 86776 637696
rect 86828 637684 86834 637696
rect 103486 637684 103514 637724
rect 124398 637712 124404 637724
rect 124456 637712 124462 637764
rect 138658 637712 138664 637764
rect 138716 637752 138722 637764
rect 168742 637752 168748 637764
rect 138716 637724 168748 637752
rect 138716 637712 138722 637724
rect 168742 637712 168748 637724
rect 168800 637712 168806 637764
rect 210510 637712 210516 637764
rect 210568 637752 210574 637764
rect 257614 637752 257620 637764
rect 210568 637724 257620 637752
rect 210568 637712 210574 637724
rect 257614 637712 257620 637724
rect 257672 637712 257678 637764
rect 121638 637684 121644 637696
rect 86828 637656 103514 637684
rect 117424 637656 121644 637684
rect 86828 637644 86834 637656
rect 59170 637576 59176 637628
rect 59228 637616 59234 637628
rect 74626 637616 74632 637628
rect 59228 637588 74632 637616
rect 59228 637576 59234 637588
rect 74626 637576 74632 637588
rect 74684 637576 74690 637628
rect 83458 637576 83464 637628
rect 83516 637616 83522 637628
rect 117424 637616 117452 637656
rect 121638 637644 121644 637656
rect 121696 637644 121702 637696
rect 138750 637644 138756 637696
rect 138808 637684 138814 637696
rect 142982 637684 142988 637696
rect 138808 637656 142988 637684
rect 138808 637644 138814 637656
rect 142982 637644 142988 637656
rect 143040 637644 143046 637696
rect 198274 637644 198280 637696
rect 198332 637684 198338 637696
rect 201494 637684 201500 637696
rect 198332 637656 201500 637684
rect 198332 637644 198338 637656
rect 201494 637644 201500 637656
rect 201552 637644 201558 637696
rect 216030 637644 216036 637696
rect 216088 637684 216094 637696
rect 219710 637684 219716 637696
rect 216088 637656 219716 637684
rect 216088 637644 216094 637656
rect 219710 637644 219716 637656
rect 219768 637644 219774 637696
rect 83516 637588 117452 637616
rect 83516 637576 83522 637588
rect 118234 637576 118240 637628
rect 118292 637616 118298 637628
rect 120902 637616 120908 637628
rect 118292 637588 120908 637616
rect 118292 637576 118298 637588
rect 120902 637576 120908 637588
rect 120960 637576 120966 637628
rect 137922 637576 137928 637628
rect 137980 637616 137986 637628
rect 218698 637616 218704 637628
rect 137980 637588 218704 637616
rect 137980 637576 137986 637588
rect 218698 637576 218704 637588
rect 218756 637576 218762 637628
rect 280706 637440 280712 637492
rect 280764 637440 280770 637492
rect 280724 637288 280752 637440
rect 280706 637236 280712 637288
rect 280764 637236 280770 637288
rect 429930 636896 429936 636948
rect 429988 636936 429994 636948
rect 474734 636936 474740 636948
rect 429988 636908 474740 636936
rect 429988 636896 429994 636908
rect 474734 636896 474740 636908
rect 474792 636896 474798 636948
rect 432598 636828 432604 636880
rect 432656 636868 432662 636880
rect 505462 636868 505468 636880
rect 432656 636840 505468 636868
rect 432656 636828 432662 636840
rect 505462 636828 505468 636840
rect 505520 636828 505526 636880
rect 482922 636216 482928 636268
rect 482980 636256 482986 636268
rect 511350 636256 511356 636268
rect 482980 636228 511356 636256
rect 482980 636216 482986 636228
rect 511350 636216 511356 636228
rect 511408 636216 511414 636268
rect 206462 634788 206468 634840
rect 206520 634828 206526 634840
rect 216674 634828 216680 634840
rect 206520 634800 216680 634828
rect 206520 634788 206526 634800
rect 216674 634788 216680 634800
rect 216732 634788 216738 634840
rect 289078 634788 289084 634840
rect 289136 634828 289142 634840
rect 317966 634828 317972 634840
rect 289136 634800 317972 634828
rect 289136 634788 289142 634800
rect 317966 634788 317972 634800
rect 318024 634788 318030 634840
rect 428458 634720 428464 634772
rect 428516 634760 428522 634772
rect 456794 634760 456800 634772
rect 428516 634732 456800 634760
rect 428516 634720 428522 634732
rect 456794 634720 456800 634732
rect 456852 634720 456858 634772
rect 208486 632068 208492 632120
rect 208544 632108 208550 632120
rect 216674 632108 216680 632120
rect 208544 632080 216680 632108
rect 208544 632068 208550 632080
rect 216674 632068 216680 632080
rect 216732 632068 216738 632120
rect 307018 630640 307024 630692
rect 307076 630680 307082 630692
rect 317414 630680 317420 630692
rect 307076 630652 317420 630680
rect 307076 630640 307082 630652
rect 317414 630640 317420 630652
rect 317472 630640 317478 630692
rect 211798 626560 211804 626612
rect 211856 626600 211862 626612
rect 216674 626600 216680 626612
rect 211856 626572 216680 626600
rect 211856 626560 211862 626572
rect 216674 626560 216680 626572
rect 216732 626560 216738 626612
rect 429838 626492 429844 626544
rect 429896 626532 429902 626544
rect 456794 626532 456800 626544
rect 429896 626504 456800 626532
rect 429896 626492 429902 626504
rect 456794 626492 456800 626504
rect 456852 626492 456858 626544
rect 311158 625132 311164 625184
rect 311216 625172 311222 625184
rect 317966 625172 317972 625184
rect 311216 625144 317972 625172
rect 311216 625132 311222 625144
rect 317966 625132 317972 625144
rect 318024 625132 318030 625184
rect 132494 622412 132500 622464
rect 132552 622452 132558 622464
rect 136634 622452 136640 622464
rect 132552 622424 136640 622452
rect 132552 622412 132558 622424
rect 136634 622412 136640 622424
rect 136692 622412 136698 622464
rect 204990 622412 204996 622464
rect 205048 622452 205054 622464
rect 216674 622452 216680 622464
rect 205048 622424 216680 622452
rect 205048 622412 205054 622424
rect 216674 622412 216680 622424
rect 216732 622412 216738 622464
rect 287790 620984 287796 621036
rect 287848 621024 287854 621036
rect 317966 621024 317972 621036
rect 287848 620996 317972 621024
rect 287848 620984 287854 620996
rect 317966 620984 317972 620996
rect 318024 620984 318030 621036
rect 135346 618196 135352 618248
rect 135404 618236 135410 618248
rect 137278 618236 137284 618248
rect 135404 618208 137284 618236
rect 135404 618196 135410 618208
rect 137278 618196 137284 618208
rect 137336 618196 137342 618248
rect 295978 615476 295984 615528
rect 296036 615516 296042 615528
rect 317414 615516 317420 615528
rect 296036 615488 317420 615516
rect 296036 615476 296042 615488
rect 317414 615476 317420 615488
rect 317472 615476 317478 615528
rect 286318 611328 286324 611380
rect 286376 611368 286382 611380
rect 317966 611368 317972 611380
rect 286376 611340 317972 611368
rect 286376 611328 286382 611340
rect 317966 611328 317972 611340
rect 318024 611328 318030 611380
rect 134518 604460 134524 604512
rect 134576 604500 134582 604512
rect 137370 604500 137376 604512
rect 134576 604472 137376 604500
rect 134576 604460 134582 604472
rect 137370 604460 137376 604472
rect 137428 604460 137434 604512
rect 213270 604460 213276 604512
rect 213328 604500 213334 604512
rect 216674 604500 216680 604512
rect 213328 604472 216680 604500
rect 213328 604460 213334 604472
rect 216674 604460 216680 604472
rect 216732 604460 216738 604512
rect 124122 603100 124128 603152
rect 124180 603140 124186 603152
rect 134610 603140 134616 603152
rect 124180 603112 134616 603140
rect 124180 603100 124186 603112
rect 134610 603100 134616 603112
rect 134668 603100 134674 603152
rect 203886 603100 203892 603152
rect 203944 603140 203950 603152
rect 216766 603140 216772 603152
rect 203944 603112 216772 603140
rect 203944 603100 203950 603112
rect 216766 603100 216772 603112
rect 216824 603100 216830 603152
rect 283650 603100 283656 603152
rect 283708 603140 283714 603152
rect 300210 603140 300216 603152
rect 283708 603112 300216 603140
rect 283708 603100 283714 603112
rect 300210 603100 300216 603112
rect 300268 603100 300274 603152
rect 211154 601672 211160 601724
rect 211212 601712 211218 601724
rect 216674 601712 216680 601724
rect 211212 601684 216680 601712
rect 211212 601672 211218 601684
rect 216674 601672 216680 601684
rect 216732 601672 216738 601724
rect 296070 601672 296076 601724
rect 296128 601712 296134 601724
rect 317966 601712 317972 601724
rect 296128 601684 317972 601712
rect 296128 601672 296134 601684
rect 317966 601672 317972 601684
rect 318024 601672 318030 601724
rect 57422 600244 57428 600296
rect 57480 600284 57486 600296
rect 58618 600284 58624 600296
rect 57480 600256 58624 600284
rect 57480 600244 57486 600256
rect 58618 600244 58624 600256
rect 58676 600244 58682 600296
rect 214558 597524 214564 597576
rect 214616 597564 214622 597576
rect 217042 597564 217048 597576
rect 214616 597536 217048 597564
rect 214616 597524 214622 597536
rect 217042 597524 217048 597536
rect 217100 597524 217106 597576
rect 286410 597524 286416 597576
rect 286468 597564 286474 597576
rect 317966 597564 317972 597576
rect 286468 597536 317972 597564
rect 286468 597524 286474 597536
rect 317966 597524 317972 597536
rect 318024 597524 318030 597576
rect 217686 595960 217692 596012
rect 217744 596000 217750 596012
rect 218698 596000 218704 596012
rect 217744 595972 218704 596000
rect 217744 595960 217750 595972
rect 218698 595960 218704 595972
rect 218756 595960 218762 596012
rect 125594 592016 125600 592068
rect 125652 592056 125658 592068
rect 136634 592056 136640 592068
rect 125652 592028 136640 592056
rect 125652 592016 125658 592028
rect 136634 592016 136640 592028
rect 136692 592016 136698 592068
rect 210602 592016 210608 592068
rect 210660 592056 210666 592068
rect 216674 592056 216680 592068
rect 210660 592028 216680 592056
rect 210660 592016 210666 592028
rect 216674 592016 216680 592028
rect 216732 592016 216738 592068
rect 300118 592016 300124 592068
rect 300176 592056 300182 592068
rect 317966 592056 317972 592068
rect 300176 592028 317972 592056
rect 300176 592016 300182 592028
rect 317966 592016 317972 592028
rect 318024 592016 318030 592068
rect 130378 589296 130384 589348
rect 130436 589336 130442 589348
rect 136634 589336 136640 589348
rect 130436 589308 136640 589336
rect 130436 589296 130442 589308
rect 136634 589296 136640 589308
rect 136692 589296 136698 589348
rect 209038 589296 209044 589348
rect 209096 589336 209102 589348
rect 216674 589336 216680 589348
rect 209096 589308 216680 589336
rect 209096 589296 209102 589308
rect 216674 589296 216680 589308
rect 216732 589296 216738 589348
rect 210694 586508 210700 586560
rect 210752 586548 210758 586560
rect 216674 586548 216680 586560
rect 210752 586520 216680 586548
rect 210752 586508 210758 586520
rect 216674 586508 216680 586520
rect 216732 586508 216738 586560
rect 289170 586508 289176 586560
rect 289228 586548 289234 586560
rect 317414 586548 317420 586560
rect 289228 586520 317420 586548
rect 289228 586508 289234 586520
rect 317414 586508 317420 586520
rect 317472 586508 317478 586560
rect 300210 584128 300216 584180
rect 300268 584168 300274 584180
rect 302234 584168 302240 584180
rect 300268 584140 302240 584168
rect 300268 584128 300274 584140
rect 302234 584128 302240 584140
rect 302292 584128 302298 584180
rect 281626 583312 281632 583364
rect 281684 583352 281690 583364
rect 282270 583352 282276 583364
rect 281684 583324 282276 583352
rect 281684 583312 281690 583324
rect 282270 583312 282276 583324
rect 282328 583312 282334 583364
rect 207014 577464 207020 577516
rect 207072 577504 207078 577516
rect 217410 577504 217416 577516
rect 207072 577476 217416 577504
rect 207072 577464 207078 577476
rect 217410 577464 217416 577476
rect 217468 577464 217474 577516
rect 57882 576172 57888 576224
rect 57940 576212 57946 576224
rect 137278 576212 137284 576224
rect 57940 576184 137284 576212
rect 57940 576172 57946 576184
rect 137278 576172 137284 576184
rect 137336 576172 137342 576224
rect 217686 576172 217692 576224
rect 217744 576212 217750 576224
rect 219894 576212 219900 576224
rect 217744 576184 219900 576212
rect 217744 576172 217750 576184
rect 219894 576172 219900 576184
rect 219952 576172 219958 576224
rect 57238 575492 57244 575544
rect 57296 575532 57302 575544
rect 60366 575532 60372 575544
rect 57296 575504 60372 575532
rect 57296 575492 57302 575504
rect 60366 575492 60372 575504
rect 60424 575492 60430 575544
rect 137370 575492 137376 575544
rect 137428 575532 137434 575544
rect 140130 575532 140136 575544
rect 137428 575504 140136 575532
rect 137428 575492 137434 575504
rect 140130 575492 140136 575504
rect 140188 575492 140194 575544
rect 200942 575492 200948 575544
rect 201000 575532 201006 575544
rect 203334 575532 203340 575544
rect 201000 575504 203340 575532
rect 201000 575492 201006 575504
rect 203334 575492 203340 575504
rect 203392 575492 203398 575544
rect 3510 575424 3516 575476
rect 3568 575464 3574 575476
rect 286410 575464 286416 575476
rect 3568 575436 286416 575464
rect 3568 575424 3574 575436
rect 286410 575424 286416 575436
rect 286468 575424 286474 575476
rect 134610 575356 134616 575408
rect 134668 575396 134674 575408
rect 216766 575396 216772 575408
rect 134668 575368 216772 575396
rect 134668 575356 134674 575368
rect 216766 575356 216772 575368
rect 216824 575396 216830 575408
rect 302234 575396 302240 575408
rect 216824 575368 302240 575396
rect 216824 575356 216830 575368
rect 302234 575356 302240 575368
rect 302292 575356 302298 575408
rect 58434 575220 58440 575272
rect 58492 575260 58498 575272
rect 62390 575260 62396 575272
rect 58492 575232 62396 575260
rect 58492 575220 58498 575232
rect 62390 575220 62396 575232
rect 62448 575220 62454 575272
rect 139210 575220 139216 575272
rect 139268 575260 139274 575272
rect 142154 575260 142160 575272
rect 139268 575232 142160 575260
rect 139268 575220 139274 575232
rect 142154 575220 142160 575232
rect 142212 575220 142218 575272
rect 139854 575152 139860 575204
rect 139912 575192 139918 575204
rect 140774 575192 140780 575204
rect 139912 575164 140780 575192
rect 139912 575152 139918 575164
rect 140774 575152 140780 575164
rect 140832 575152 140838 575204
rect 164326 575152 164332 575204
rect 164384 575192 164390 575204
rect 200850 575192 200856 575204
rect 164384 575164 200856 575192
rect 164384 575152 164390 575164
rect 200850 575152 200856 575164
rect 200908 575152 200914 575204
rect 106274 575084 106280 575136
rect 106332 575124 106338 575136
rect 124582 575124 124588 575136
rect 106332 575096 124588 575124
rect 106332 575084 106338 575096
rect 124582 575084 124588 575096
rect 124640 575084 124646 575136
rect 137646 575084 137652 575136
rect 137704 575124 137710 575136
rect 145466 575124 145472 575136
rect 137704 575096 145472 575124
rect 137704 575084 137710 575096
rect 145466 575084 145472 575096
rect 145524 575084 145530 575136
rect 183462 575084 183468 575136
rect 183520 575124 183526 575136
rect 218882 575124 218888 575136
rect 183520 575096 218888 575124
rect 183520 575084 183526 575096
rect 218882 575084 218888 575096
rect 218940 575084 218946 575136
rect 100386 575016 100392 575068
rect 100444 575056 100450 575068
rect 121546 575056 121552 575068
rect 100444 575028 121552 575056
rect 100444 575016 100450 575028
rect 121546 575016 121552 575028
rect 121604 575016 121610 575068
rect 156230 575016 156236 575068
rect 156288 575056 156294 575068
rect 205634 575056 205640 575068
rect 156288 575028 205640 575056
rect 156288 575016 156294 575028
rect 205634 575016 205640 575028
rect 205692 575016 205698 575068
rect 98178 574948 98184 575000
rect 98236 574988 98242 575000
rect 122834 574988 122840 575000
rect 98236 574960 122840 574988
rect 98236 574948 98242 574960
rect 122834 574948 122840 574960
rect 122892 574948 122898 575000
rect 138842 574948 138848 575000
rect 138900 574988 138906 575000
rect 149146 574988 149152 575000
rect 138900 574960 149152 574988
rect 138900 574948 138906 574960
rect 149146 574948 149152 574960
rect 149204 574948 149210 575000
rect 154574 574948 154580 575000
rect 154632 574988 154638 575000
rect 204346 574988 204352 575000
rect 154632 574960 204352 574988
rect 154632 574948 154638 574960
rect 204346 574948 204352 574960
rect 204404 574948 204410 575000
rect 219342 574948 219348 575000
rect 219400 574988 219406 575000
rect 223574 574988 223580 575000
rect 219400 574960 223580 574988
rect 219400 574948 219406 574960
rect 223574 574948 223580 574960
rect 223632 574948 223638 575000
rect 273254 574948 273260 575000
rect 273312 574988 273318 575000
rect 318242 574988 318248 575000
rect 273312 574960 318248 574988
rect 273312 574948 273318 574960
rect 318242 574948 318248 574960
rect 318300 574948 318306 575000
rect 54846 574880 54852 574932
rect 54904 574920 54910 574932
rect 78674 574920 78680 574932
rect 54904 574892 78680 574920
rect 54904 574880 54910 574892
rect 78674 574880 78680 574892
rect 78732 574880 78738 574932
rect 97442 574880 97448 574932
rect 97500 574920 97506 574932
rect 124674 574920 124680 574932
rect 97500 574892 124680 574920
rect 97500 574880 97506 574892
rect 124674 574880 124680 574892
rect 124732 574880 124738 574932
rect 129734 574880 129740 574932
rect 129792 574920 129798 574932
rect 202966 574920 202972 574932
rect 129792 574892 202972 574920
rect 129792 574880 129798 574892
rect 202966 574880 202972 574892
rect 203024 574880 203030 574932
rect 217870 574880 217876 574932
rect 217928 574920 217934 574932
rect 222194 574920 222200 574932
rect 217928 574892 222200 574920
rect 217928 574880 217934 574892
rect 222194 574880 222200 574892
rect 222252 574880 222258 574932
rect 229278 574880 229284 574932
rect 229336 574920 229342 574932
rect 281258 574920 281264 574932
rect 229336 574892 281264 574920
rect 229336 574880 229342 574892
rect 281258 574880 281264 574892
rect 281316 574880 281322 574932
rect 57606 574812 57612 574864
rect 57664 574852 57670 574864
rect 83182 574852 83188 574864
rect 57664 574824 83188 574852
rect 57664 574812 57670 574824
rect 83182 574812 83188 574824
rect 83240 574812 83246 574864
rect 93854 574812 93860 574864
rect 93912 574852 93918 574864
rect 124490 574852 124496 574864
rect 93912 574824 124496 574852
rect 93912 574812 93918 574824
rect 124490 574812 124496 574824
rect 124548 574812 124554 574864
rect 134978 574812 134984 574864
rect 135036 574852 135042 574864
rect 151906 574852 151912 574864
rect 135036 574824 151912 574852
rect 135036 574812 135042 574824
rect 151906 574812 151912 574824
rect 151964 574812 151970 574864
rect 197078 574812 197084 574864
rect 197136 574852 197142 574864
rect 281994 574852 282000 574864
rect 197136 574824 282000 574852
rect 197136 574812 197142 574824
rect 281994 574812 282000 574824
rect 282052 574812 282058 574864
rect 63494 574744 63500 574796
rect 63552 574784 63558 574796
rect 123570 574784 123576 574796
rect 63552 574756 123576 574784
rect 63552 574744 63558 574756
rect 123570 574744 123576 574756
rect 123628 574744 123634 574796
rect 134886 574744 134892 574796
rect 134944 574784 134950 574796
rect 161934 574784 161940 574796
rect 134944 574756 161940 574784
rect 134944 574744 134950 574756
rect 161934 574744 161940 574756
rect 161992 574744 161998 574796
rect 179414 574744 179420 574796
rect 179472 574784 179478 574796
rect 281626 574784 281632 574796
rect 179472 574756 281632 574784
rect 179472 574744 179478 574756
rect 281626 574744 281632 574756
rect 281684 574744 281690 574796
rect 58802 574268 58808 574320
rect 58860 574308 58866 574320
rect 60918 574308 60924 574320
rect 58860 574280 60924 574308
rect 58860 574268 58866 574280
rect 60918 574268 60924 574280
rect 60976 574268 60982 574320
rect 139026 574200 139032 574252
rect 139084 574240 139090 574252
rect 141234 574240 141240 574252
rect 139084 574212 141240 574240
rect 139084 574200 139090 574212
rect 141234 574200 141240 574212
rect 141292 574200 141298 574252
rect 302234 574064 302240 574116
rect 302292 574104 302298 574116
rect 302970 574104 302976 574116
rect 302292 574076 302976 574104
rect 302292 574064 302298 574076
rect 302970 574064 302976 574076
rect 303028 574064 303034 574116
rect 59446 573860 59452 573912
rect 59504 573900 59510 573912
rect 63218 573900 63224 573912
rect 59504 573872 63224 573900
rect 59504 573860 59510 573872
rect 63218 573860 63224 573872
rect 63276 573860 63282 573912
rect 112530 573656 112536 573708
rect 112588 573696 112594 573708
rect 123018 573696 123024 573708
rect 112588 573668 123024 573696
rect 112588 573656 112594 573668
rect 123018 573656 123024 573668
rect 123076 573656 123082 573708
rect 88150 573588 88156 573640
rect 88208 573628 88214 573640
rect 120902 573628 120908 573640
rect 88208 573600 120908 573628
rect 88208 573588 88214 573600
rect 120902 573588 120908 573600
rect 120960 573588 120966 573640
rect 128998 573588 129004 573640
rect 129056 573628 129062 573640
rect 203150 573628 203156 573640
rect 129056 573600 203156 573628
rect 129056 573588 129062 573600
rect 203150 573588 203156 573600
rect 203208 573588 203214 573640
rect 57146 573520 57152 573572
rect 57204 573560 57210 573572
rect 81710 573560 81716 573572
rect 57204 573532 81716 573560
rect 57204 573520 57210 573532
rect 81710 573520 81716 573532
rect 81768 573520 81774 573572
rect 86954 573520 86960 573572
rect 87012 573560 87018 573572
rect 121454 573560 121460 573572
rect 87012 573532 121460 573560
rect 87012 573520 87018 573532
rect 121454 573520 121460 573532
rect 121512 573520 121518 573572
rect 126146 573520 126152 573572
rect 126204 573560 126210 573572
rect 201954 573560 201960 573572
rect 126204 573532 201960 573560
rect 126204 573520 126210 573532
rect 201954 573520 201960 573532
rect 202012 573520 202018 573572
rect 219250 573520 219256 573572
rect 219308 573560 219314 573572
rect 224310 573560 224316 573572
rect 219308 573532 224316 573560
rect 219308 573520 219314 573532
rect 224310 573520 224316 573532
rect 224368 573520 224374 573572
rect 240778 573520 240784 573572
rect 240836 573560 240842 573572
rect 315298 573560 315304 573572
rect 240836 573532 315304 573560
rect 240836 573520 240842 573532
rect 315298 573520 315304 573532
rect 315356 573520 315362 573572
rect 59262 573452 59268 573504
rect 59320 573492 59326 573504
rect 68830 573492 68836 573504
rect 59320 573464 68836 573492
rect 59320 573452 59326 573464
rect 68830 573452 68836 573464
rect 68888 573452 68894 573504
rect 78858 573452 78864 573504
rect 78916 573492 78922 573504
rect 122282 573492 122288 573504
rect 78916 573464 122288 573492
rect 78916 573452 78922 573464
rect 122282 573452 122288 573464
rect 122340 573452 122346 573504
rect 186314 573452 186320 573504
rect 186372 573492 186378 573504
rect 282914 573492 282920 573504
rect 186372 573464 282920 573492
rect 186372 573452 186378 573464
rect 282914 573452 282920 573464
rect 282972 573452 282978 573504
rect 67634 573384 67640 573436
rect 67692 573424 67698 573436
rect 121822 573424 121828 573436
rect 67692 573396 121828 573424
rect 67692 573384 67698 573396
rect 121822 573384 121828 573396
rect 121880 573384 121886 573436
rect 139118 573384 139124 573436
rect 139176 573424 139182 573436
rect 150618 573424 150624 573436
rect 139176 573396 150624 573424
rect 139176 573384 139182 573396
rect 150618 573384 150624 573396
rect 150676 573384 150682 573436
rect 182266 573384 182272 573436
rect 182324 573424 182330 573436
rect 281534 573424 281540 573436
rect 182324 573396 281540 573424
rect 182324 573384 182330 573396
rect 281534 573384 281540 573396
rect 281592 573384 281598 573436
rect 64506 573316 64512 573368
rect 64564 573356 64570 573368
rect 122926 573356 122932 573368
rect 64564 573328 122932 573356
rect 64564 573316 64570 573328
rect 122926 573316 122932 573328
rect 122984 573316 122990 573368
rect 137002 573316 137008 573368
rect 137060 573356 137066 573368
rect 160554 573356 160560 573368
rect 137060 573328 160560 573356
rect 137060 573316 137066 573328
rect 160554 573316 160560 573328
rect 160612 573316 160618 573368
rect 180794 573316 180800 573368
rect 180852 573356 180858 573368
rect 283374 573356 283380 573368
rect 180852 573328 283380 573356
rect 180852 573316 180858 573328
rect 283374 573316 283380 573328
rect 283432 573316 283438 573368
rect 268010 572704 268016 572756
rect 268068 572744 268074 572756
rect 317966 572744 317972 572756
rect 268068 572716 317972 572744
rect 268068 572704 268074 572716
rect 317966 572704 317972 572716
rect 318024 572704 318030 572756
rect 150986 572500 150992 572552
rect 151044 572540 151050 572552
rect 160738 572540 160744 572552
rect 151044 572512 160744 572540
rect 151044 572500 151050 572512
rect 160738 572500 160744 572512
rect 160796 572500 160802 572552
rect 197998 572500 198004 572552
rect 198056 572540 198062 572552
rect 200574 572540 200580 572552
rect 198056 572512 200580 572540
rect 198056 572500 198062 572512
rect 200574 572500 200580 572512
rect 200632 572500 200638 572552
rect 266998 572500 267004 572552
rect 267056 572540 267062 572552
rect 268930 572540 268936 572552
rect 267056 572512 268936 572540
rect 267056 572500 267062 572512
rect 268930 572500 268936 572512
rect 268988 572500 268994 572552
rect 148410 572432 148416 572484
rect 148468 572472 148474 572484
rect 159358 572472 159364 572484
rect 148468 572444 159364 572472
rect 148468 572432 148474 572444
rect 159358 572432 159364 572444
rect 159416 572432 159422 572484
rect 143534 572364 143540 572416
rect 143592 572404 143598 572416
rect 156782 572404 156788 572416
rect 143592 572376 156788 572404
rect 143592 572364 143598 572376
rect 156782 572364 156788 572376
rect 156840 572364 156846 572416
rect 160002 572364 160008 572416
rect 160060 572404 160066 572416
rect 164878 572404 164884 572416
rect 160060 572376 164884 572404
rect 160060 572364 160066 572376
rect 164878 572364 164884 572376
rect 164936 572364 164942 572416
rect 82538 572296 82544 572348
rect 82596 572336 82602 572348
rect 88978 572336 88984 572348
rect 82596 572308 88984 572336
rect 82596 572296 82602 572308
rect 88978 572296 88984 572308
rect 89036 572296 89042 572348
rect 147674 572296 147680 572348
rect 147732 572336 147738 572348
rect 162578 572336 162584 572348
rect 147732 572308 162584 572336
rect 147732 572296 147738 572308
rect 162578 572296 162584 572308
rect 162636 572296 162642 572348
rect 74534 572228 74540 572280
rect 74592 572268 74598 572280
rect 97350 572268 97356 572280
rect 74592 572240 97356 572268
rect 74592 572228 74598 572240
rect 97350 572228 97356 572240
rect 97408 572228 97414 572280
rect 99926 572228 99932 572280
rect 99984 572268 99990 572280
rect 115474 572268 115480 572280
rect 99984 572240 115480 572268
rect 99984 572228 99990 572240
rect 115474 572228 115480 572240
rect 115532 572228 115538 572280
rect 154850 572228 154856 572280
rect 154908 572268 154914 572280
rect 171594 572268 171600 572280
rect 154908 572240 171600 572268
rect 154908 572228 154914 572240
rect 171594 572228 171600 572240
rect 171652 572228 171658 572280
rect 232222 572228 232228 572280
rect 232280 572268 232286 572280
rect 259914 572268 259920 572280
rect 232280 572240 259920 572268
rect 232280 572228 232286 572240
rect 259914 572228 259920 572240
rect 259972 572228 259978 572280
rect 62574 572160 62580 572212
rect 62632 572200 62638 572212
rect 71038 572200 71044 572212
rect 62632 572172 71044 572200
rect 62632 572160 62638 572172
rect 71038 572160 71044 572172
rect 71096 572160 71102 572212
rect 85758 572160 85764 572212
rect 85816 572200 85822 572212
rect 108298 572200 108304 572212
rect 85816 572172 108304 572200
rect 85816 572160 85822 572172
rect 108298 572160 108304 572172
rect 108356 572160 108362 572212
rect 129826 572160 129832 572212
rect 129884 572200 129890 572212
rect 154206 572200 154212 572212
rect 129884 572172 154212 572200
rect 129884 572160 129890 572172
rect 154206 572160 154212 572172
rect 154264 572160 154270 572212
rect 158714 572160 158720 572212
rect 158772 572200 158778 572212
rect 183186 572200 183192 572212
rect 158772 572172 183192 572200
rect 158772 572160 158778 572172
rect 183186 572160 183192 572172
rect 183244 572160 183250 572212
rect 188338 572160 188344 572212
rect 188396 572200 188402 572212
rect 203426 572200 203432 572212
rect 188396 572172 203432 572200
rect 188396 572160 188402 572172
rect 203426 572160 203432 572172
rect 203484 572160 203490 572212
rect 222286 572160 222292 572212
rect 222344 572200 222350 572212
rect 254118 572200 254124 572212
rect 222344 572172 254124 572200
rect 222344 572160 222350 572172
rect 254118 572160 254124 572172
rect 254176 572160 254182 572212
rect 269666 572160 269672 572212
rect 269724 572200 269730 572212
rect 286318 572200 286324 572212
rect 269724 572172 286324 572200
rect 269724 572160 269730 572172
rect 286318 572160 286324 572172
rect 286376 572160 286382 572212
rect 68370 572092 68376 572144
rect 68428 572132 68434 572144
rect 105538 572132 105544 572144
rect 68428 572104 105544 572132
rect 68428 572092 68434 572104
rect 105538 572092 105544 572104
rect 105596 572092 105602 572144
rect 119706 572092 119712 572144
rect 119764 572132 119770 572144
rect 145190 572132 145196 572144
rect 119764 572104 145196 572132
rect 119764 572092 119770 572104
rect 145190 572092 145196 572104
rect 145248 572092 145254 572144
rect 147766 572092 147772 572144
rect 147824 572132 147830 572144
rect 185762 572132 185768 572144
rect 147824 572104 185768 572132
rect 147824 572092 147830 572104
rect 185762 572092 185768 572104
rect 185820 572092 185826 572144
rect 190454 572092 190460 572144
rect 190512 572132 190518 572144
rect 257338 572132 257344 572144
rect 190512 572104 257344 572132
rect 190512 572092 190518 572104
rect 257338 572092 257344 572104
rect 257396 572092 257402 572144
rect 263686 572092 263692 572144
rect 263744 572132 263750 572144
rect 312538 572132 312544 572144
rect 263744 572104 312544 572132
rect 263744 572092 263750 572104
rect 312538 572092 312544 572104
rect 312596 572092 312602 572144
rect 70946 572024 70952 572076
rect 71004 572064 71010 572076
rect 108390 572064 108396 572076
rect 71004 572036 108396 572064
rect 71004 572024 71010 572036
rect 108390 572024 108396 572036
rect 108448 572024 108454 572076
rect 110414 572024 110420 572076
rect 110472 572064 110478 572076
rect 120718 572064 120724 572076
rect 110472 572036 120724 572064
rect 110472 572024 110478 572036
rect 120718 572024 120724 572036
rect 120776 572024 120782 572076
rect 134150 572024 134156 572076
rect 134208 572064 134214 572076
rect 197354 572064 197360 572076
rect 134208 572036 197360 572064
rect 134208 572024 134214 572036
rect 197354 572024 197360 572036
rect 197412 572024 197418 572076
rect 227898 572024 227904 572076
rect 227956 572064 227962 572076
rect 245746 572064 245752 572076
rect 227956 572036 245752 572064
rect 227956 572024 227962 572036
rect 245746 572024 245752 572036
rect 245804 572024 245810 572076
rect 247034 572024 247040 572076
rect 247092 572064 247098 572076
rect 319806 572064 319812 572076
rect 247092 572036 319812 572064
rect 247092 572024 247098 572036
rect 319806 572024 319812 572036
rect 319864 572024 319870 572076
rect 58894 571956 58900 572008
rect 58952 571996 58958 572008
rect 74626 571996 74632 572008
rect 58952 571968 74632 571996
rect 58952 571956 58958 571968
rect 74626 571956 74632 571968
rect 74684 571956 74690 572008
rect 76834 571956 76840 572008
rect 76892 571996 76898 572008
rect 117314 571996 117320 572008
rect 76892 571968 117320 571996
rect 76892 571956 76898 571968
rect 117314 571956 117320 571968
rect 117372 571956 117378 572008
rect 132678 571956 132684 572008
rect 132736 571996 132742 572008
rect 177390 571996 177396 572008
rect 132736 571968 177396 571996
rect 132736 571956 132742 571968
rect 177390 571956 177396 571968
rect 177448 571956 177454 572008
rect 192754 571956 192760 572008
rect 192812 571996 192818 572008
rect 277302 571996 277308 572008
rect 192812 571968 277308 571996
rect 192812 571956 192818 571968
rect 277302 571956 277308 571968
rect 277360 571956 277366 572008
rect 113266 571616 113272 571668
rect 113324 571656 113330 571668
rect 121086 571656 121092 571668
rect 113324 571628 121092 571656
rect 113324 571616 113330 571628
rect 121086 571616 121092 571628
rect 121144 571616 121150 571668
rect 94130 571412 94136 571464
rect 94188 571452 94194 571464
rect 101398 571452 101404 571464
rect 94188 571424 101404 571452
rect 94188 571412 94194 571424
rect 101398 571412 101404 571424
rect 101456 571412 101462 571464
rect 262858 571412 262864 571464
rect 262916 571452 262922 571464
rect 265710 571452 265716 571464
rect 262916 571424 265716 571452
rect 262916 571412 262922 571424
rect 265710 571412 265716 571424
rect 265768 571412 265774 571464
rect 59998 571344 60004 571396
rect 60056 571384 60062 571396
rect 61378 571384 61384 571396
rect 60056 571356 61384 571384
rect 60056 571344 60062 571356
rect 61378 571344 61384 571356
rect 61436 571344 61442 571396
rect 72418 571344 72424 571396
rect 72476 571384 72482 571396
rect 74166 571384 74172 571396
rect 72476 571356 74172 571384
rect 72476 571344 72482 571356
rect 74166 571344 74172 571356
rect 74224 571344 74230 571396
rect 76742 571344 76748 571396
rect 76800 571384 76806 571396
rect 83458 571384 83464 571396
rect 76800 571356 83464 571384
rect 76800 571344 76806 571356
rect 83458 571344 83464 571356
rect 83516 571344 83522 571396
rect 91554 571344 91560 571396
rect 91612 571384 91618 571396
rect 93118 571384 93124 571396
rect 91612 571356 93124 571384
rect 91612 571344 91618 571356
rect 93118 571344 93124 571356
rect 93176 571344 93182 571396
rect 100754 571344 100760 571396
rect 100812 571384 100818 571396
rect 103146 571384 103152 571396
rect 100812 571356 103152 571384
rect 100812 571344 100818 571356
rect 103146 571344 103152 571356
rect 103204 571344 103210 571396
rect 106918 571344 106924 571396
rect 106976 571384 106982 571396
rect 108942 571384 108948 571396
rect 106976 571356 108948 571384
rect 106976 571344 106982 571356
rect 108942 571344 108948 571356
rect 109000 571344 109006 571396
rect 116578 571344 116584 571396
rect 116636 571384 116642 571396
rect 120534 571384 120540 571396
rect 116636 571356 120540 571384
rect 116636 571344 116642 571356
rect 120534 571344 120540 571356
rect 120592 571344 120598 571396
rect 165798 571344 165804 571396
rect 165856 571384 165862 571396
rect 167822 571384 167828 571396
rect 165856 571356 167828 571384
rect 165856 571344 165862 571356
rect 167822 571344 167828 571356
rect 167880 571344 167886 571396
rect 171778 571344 171784 571396
rect 171836 571384 171842 571396
rect 174170 571384 174176 571396
rect 171836 571356 174176 571384
rect 171836 571344 171842 571356
rect 174170 571344 174176 571356
rect 174228 571344 174234 571396
rect 184198 571344 184204 571396
rect 184256 571384 184262 571396
rect 188982 571384 188988 571396
rect 184256 571356 188988 571384
rect 184256 571344 184262 571356
rect 188982 571344 188988 571356
rect 189040 571344 189046 571396
rect 219986 571344 219992 571396
rect 220044 571384 220050 571396
rect 221458 571384 221464 571396
rect 220044 571356 221464 571384
rect 220044 571344 220050 571356
rect 221458 571344 221464 571356
rect 221516 571344 221522 571396
rect 222562 571344 222568 571396
rect 222620 571384 222626 571396
rect 224954 571384 224960 571396
rect 222620 571356 224960 571384
rect 222620 571344 222626 571356
rect 224954 571344 224960 571356
rect 225012 571344 225018 571396
rect 225046 571344 225052 571396
rect 225104 571384 225110 571396
rect 228358 571384 228364 571396
rect 225104 571356 228364 571384
rect 225104 571344 225110 571356
rect 228358 571344 228364 571356
rect 228416 571344 228422 571396
rect 260098 571344 260104 571396
rect 260156 571384 260162 571396
rect 263134 571384 263140 571396
rect 260156 571356 263140 571384
rect 260156 571344 260162 571356
rect 263134 571344 263140 571356
rect 263192 571344 263198 571396
rect 269758 571344 269764 571396
rect 269816 571384 269822 571396
rect 271506 571384 271512 571396
rect 269816 571356 271512 571384
rect 269816 571344 269822 571356
rect 271506 571344 271512 571356
rect 271564 571344 271570 571396
rect 278038 571344 278044 571396
rect 278096 571384 278102 571396
rect 280522 571384 280528 571396
rect 278096 571356 280528 571384
rect 278096 571344 278102 571356
rect 280522 571344 280528 571356
rect 280580 571344 280586 571396
rect 193214 570868 193220 570920
rect 193272 570908 193278 570920
rect 218790 570908 218796 570920
rect 193272 570880 218796 570908
rect 193272 570868 193278 570880
rect 218790 570868 218796 570880
rect 218848 570868 218854 570920
rect 94590 570800 94596 570852
rect 94648 570840 94654 570852
rect 123294 570840 123300 570852
rect 94648 570812 123300 570840
rect 94648 570800 94654 570812
rect 123294 570800 123300 570812
rect 123352 570800 123358 570852
rect 168466 570800 168472 570852
rect 168524 570840 168530 570852
rect 200666 570840 200672 570852
rect 168524 570812 200672 570840
rect 168524 570800 168530 570812
rect 200666 570800 200672 570812
rect 200724 570800 200730 570852
rect 57330 570732 57336 570784
rect 57388 570772 57394 570784
rect 89806 570772 89812 570784
rect 57388 570744 89812 570772
rect 57388 570732 57394 570744
rect 89806 570732 89812 570744
rect 89864 570732 89870 570784
rect 122834 570732 122840 570784
rect 122892 570772 122898 570784
rect 202138 570772 202144 570784
rect 122892 570744 202144 570772
rect 122892 570732 122898 570744
rect 202138 570732 202144 570744
rect 202196 570732 202202 570784
rect 215846 570732 215852 570784
rect 215904 570772 215910 570784
rect 281166 570772 281172 570784
rect 215904 570744 281172 570772
rect 215904 570732 215910 570744
rect 281166 570732 281172 570744
rect 281224 570732 281230 570784
rect 65978 570664 65984 570716
rect 66036 570704 66042 570716
rect 121914 570704 121920 570716
rect 66036 570676 121920 570704
rect 66036 570664 66042 570676
rect 121914 570664 121920 570676
rect 121972 570664 121978 570716
rect 137922 570664 137928 570716
rect 137980 570704 137986 570716
rect 169110 570704 169116 570716
rect 137980 570676 169116 570704
rect 137980 570664 137986 570676
rect 169110 570664 169116 570676
rect 169168 570664 169174 570716
rect 180610 570664 180616 570716
rect 180668 570704 180674 570716
rect 282270 570704 282276 570716
rect 180668 570676 282276 570704
rect 180668 570664 180674 570676
rect 282270 570664 282276 570676
rect 282328 570664 282334 570716
rect 7558 570596 7564 570648
rect 7616 570636 7622 570648
rect 317506 570636 317512 570648
rect 7616 570608 317512 570636
rect 7616 570596 7622 570608
rect 317506 570596 317512 570608
rect 317564 570596 317570 570648
rect 266630 569440 266636 569492
rect 266688 569480 266694 569492
rect 298738 569480 298744 569492
rect 266688 569452 298744 569480
rect 266688 569440 266694 569452
rect 298738 569440 298744 569452
rect 298796 569440 298802 569492
rect 59078 569372 59084 569424
rect 59136 569412 59142 569424
rect 92566 569412 92572 569424
rect 59136 569384 92572 569412
rect 59136 569372 59142 569384
rect 92566 569372 92572 569384
rect 92624 569372 92630 569424
rect 138290 569372 138296 569424
rect 138348 569412 138354 569424
rect 200758 569412 200764 569424
rect 138348 569384 200764 569412
rect 138348 569372 138354 569384
rect 200758 569372 200764 569384
rect 200816 569372 200822 569424
rect 250070 569372 250076 569424
rect 250128 569412 250134 569424
rect 295978 569412 295984 569424
rect 250128 569384 295984 569412
rect 250128 569372 250134 569384
rect 295978 569372 295984 569384
rect 296036 569372 296042 569424
rect 79962 569304 79968 569356
rect 80020 569344 80026 569356
rect 114738 569344 114744 569356
rect 80020 569316 114744 569344
rect 80020 569304 80026 569316
rect 114738 569304 114744 569316
rect 114796 569304 114802 569356
rect 195238 569304 195244 569356
rect 195296 569344 195302 569356
rect 283006 569344 283012 569356
rect 195296 569316 283012 569344
rect 195296 569304 195302 569316
rect 283006 569304 283012 569316
rect 283064 569304 283070 569356
rect 69014 569236 69020 569288
rect 69072 569276 69078 569288
rect 123478 569276 123484 569288
rect 69072 569248 123484 569276
rect 69072 569236 69078 569248
rect 123478 569236 123484 569248
rect 123536 569236 123542 569288
rect 138474 569236 138480 569288
rect 138532 569276 138538 569288
rect 159082 569276 159088 569288
rect 138532 569248 159088 569276
rect 138532 569236 138538 569248
rect 159082 569236 159088 569248
rect 159140 569236 159146 569288
rect 181346 569236 181352 569288
rect 181404 569276 181410 569288
rect 281902 569276 281908 569288
rect 181404 569248 281908 569276
rect 181404 569236 181410 569248
rect 281902 569236 281908 569248
rect 281960 569236 281966 569288
rect 3418 569168 3424 569220
rect 3476 569208 3482 569220
rect 319806 569208 319812 569220
rect 3476 569180 319812 569208
rect 3476 569168 3482 569180
rect 319806 569168 319812 569180
rect 319864 569168 319870 569220
rect 193490 568012 193496 568064
rect 193548 568052 193554 568064
rect 206462 568052 206468 568064
rect 193548 568024 206468 568052
rect 193548 568012 193554 568024
rect 206462 568012 206468 568024
rect 206520 568012 206526 568064
rect 259454 568012 259460 568064
rect 259512 568052 259518 568064
rect 302878 568052 302884 568064
rect 259512 568024 302884 568052
rect 259512 568012 259518 568024
rect 302878 568012 302884 568024
rect 302936 568012 302942 568064
rect 170582 567944 170588 567996
rect 170640 567984 170646 567996
rect 201770 567984 201776 567996
rect 170640 567956 201776 567984
rect 170640 567944 170646 567956
rect 201770 567944 201776 567956
rect 201828 567944 201834 567996
rect 255314 567944 255320 567996
rect 255372 567984 255378 567996
rect 309778 567984 309784 567996
rect 255372 567956 309784 567984
rect 255372 567944 255378 567956
rect 309778 567944 309784 567956
rect 309836 567944 309842 567996
rect 57054 567876 57060 567928
rect 57112 567916 57118 567928
rect 101490 567916 101496 567928
rect 57112 567888 101496 567916
rect 57112 567876 57118 567888
rect 101490 567876 101496 567888
rect 101548 567876 101554 567928
rect 187050 567876 187056 567928
rect 187108 567916 187114 567928
rect 283282 567916 283288 567928
rect 187108 567888 283288 567916
rect 187108 567876 187114 567888
rect 283282 567876 283288 567888
rect 283340 567876 283346 567928
rect 70946 567808 70952 567860
rect 71004 567848 71010 567860
rect 123202 567848 123208 567860
rect 71004 567820 123208 567848
rect 71004 567808 71010 567820
rect 123202 567808 123208 567820
rect 123260 567808 123266 567860
rect 137094 567808 137100 567860
rect 137152 567848 137158 567860
rect 166258 567848 166264 567860
rect 137152 567820 166264 567848
rect 137152 567808 137158 567820
rect 166258 567808 166264 567820
rect 166316 567808 166322 567860
rect 183554 567808 183560 567860
rect 183612 567848 183618 567860
rect 281718 567848 281724 567860
rect 183612 567820 281724 567848
rect 183612 567808 183618 567820
rect 281718 567808 281724 567820
rect 281776 567808 281782 567860
rect 11698 567196 11704 567248
rect 11756 567236 11762 567248
rect 317966 567236 317972 567248
rect 11756 567208 317972 567236
rect 11756 567196 11762 567208
rect 317966 567196 317972 567208
rect 318024 567196 318030 567248
rect 266538 566720 266544 566772
rect 266596 566760 266602 566772
rect 284938 566760 284944 566772
rect 266596 566732 284944 566760
rect 266596 566720 266602 566732
rect 284938 566720 284944 566732
rect 284996 566720 285002 566772
rect 84562 566652 84568 566704
rect 84620 566692 84626 566704
rect 122098 566692 122104 566704
rect 84620 566664 122104 566692
rect 84620 566652 84626 566664
rect 122098 566652 122104 566664
rect 122156 566652 122162 566704
rect 157978 566652 157984 566704
rect 158036 566692 158042 566704
rect 203058 566692 203064 566704
rect 158036 566664 203064 566692
rect 158036 566652 158042 566664
rect 203058 566652 203064 566664
rect 203116 566652 203122 566704
rect 226426 566652 226432 566704
rect 226484 566692 226490 566704
rect 280798 566692 280804 566704
rect 226484 566664 280804 566692
rect 226484 566652 226490 566664
rect 280798 566652 280804 566664
rect 280856 566652 280862 566704
rect 188062 566584 188068 566636
rect 188120 566624 188126 566636
rect 233234 566624 233240 566636
rect 188120 566596 233240 566624
rect 188120 566584 188126 566596
rect 233234 566584 233240 566596
rect 233292 566584 233298 566636
rect 257982 566584 257988 566636
rect 258040 566624 258046 566636
rect 314010 566624 314016 566636
rect 258040 566596 314016 566624
rect 258040 566584 258046 566596
rect 314010 566584 314016 566596
rect 314068 566584 314074 566636
rect 58986 566516 58992 566568
rect 59044 566556 59050 566568
rect 108206 566556 108212 566568
rect 59044 566528 108212 566556
rect 59044 566516 59050 566528
rect 108206 566516 108212 566528
rect 108264 566516 108270 566568
rect 122558 566516 122564 566568
rect 122616 566556 122622 566568
rect 201586 566556 201592 566568
rect 122616 566528 201592 566556
rect 122616 566516 122622 566528
rect 201586 566516 201592 566528
rect 201644 566516 201650 566568
rect 213914 566516 213920 566568
rect 213972 566556 213978 566568
rect 215018 566556 215024 566568
rect 213972 566528 215024 566556
rect 213972 566516 213978 566528
rect 215018 566516 215024 566528
rect 215076 566516 215082 566568
rect 245102 566516 245108 566568
rect 245160 566556 245166 566568
rect 313918 566556 313924 566568
rect 245160 566528 313924 566556
rect 245160 566516 245166 566528
rect 313918 566516 313924 566528
rect 313976 566516 313982 566568
rect 65242 566448 65248 566500
rect 65300 566488 65306 566500
rect 123386 566488 123392 566500
rect 65300 566460 123392 566488
rect 65300 566448 65306 566460
rect 123386 566448 123392 566460
rect 123444 566448 123450 566500
rect 138566 566448 138572 566500
rect 138624 566488 138630 566500
rect 160646 566488 160652 566500
rect 138624 566460 160652 566488
rect 138624 566448 138630 566460
rect 160646 566448 160652 566460
rect 160704 566448 160710 566500
rect 194962 566448 194968 566500
rect 195020 566488 195026 566500
rect 283558 566488 283564 566500
rect 195020 566460 283564 566488
rect 195020 566448 195026 566460
rect 283558 566448 283564 566460
rect 283616 566448 283622 566500
rect 220722 565360 220728 565412
rect 220780 565400 220786 565412
rect 247126 565400 247132 565412
rect 220780 565372 247132 565400
rect 220780 565360 220786 565372
rect 247126 565360 247132 565372
rect 247184 565360 247190 565412
rect 190638 565292 190644 565344
rect 190696 565332 190702 565344
rect 204990 565332 204996 565344
rect 190696 565304 204996 565332
rect 190696 565292 190702 565304
rect 204990 565292 204996 565304
rect 205048 565292 205054 565344
rect 228634 565292 228640 565344
rect 228692 565332 228698 565344
rect 282086 565332 282092 565344
rect 228692 565304 282092 565332
rect 228692 565292 228698 565304
rect 282086 565292 282092 565304
rect 282144 565292 282150 565344
rect 88334 565224 88340 565276
rect 88392 565264 88398 565276
rect 104618 565264 104624 565276
rect 88392 565236 104624 565264
rect 88392 565224 88398 565236
rect 104618 565224 104624 565236
rect 104676 565224 104682 565276
rect 177022 565224 177028 565276
rect 177080 565264 177086 565276
rect 213270 565264 213276 565276
rect 177080 565236 213276 565264
rect 177080 565224 177086 565236
rect 213270 565224 213276 565236
rect 213328 565224 213334 565276
rect 246482 565224 246488 565276
rect 246540 565264 246546 565276
rect 311158 565264 311164 565276
rect 246540 565236 311164 565264
rect 246540 565224 246546 565236
rect 311158 565224 311164 565236
rect 311216 565224 311222 565276
rect 71038 565156 71044 565208
rect 71096 565196 71102 565208
rect 109678 565196 109684 565208
rect 71096 565168 109684 565196
rect 71096 565156 71102 565168
rect 109678 565156 109684 565168
rect 109736 565156 109742 565208
rect 142614 565156 142620 565208
rect 142672 565196 142678 565208
rect 202046 565196 202052 565208
rect 142672 565168 202052 565196
rect 142672 565156 142678 565168
rect 202046 565156 202052 565168
rect 202104 565156 202110 565208
rect 206370 565156 206376 565208
rect 206428 565196 206434 565208
rect 241514 565196 241520 565208
rect 206428 565168 241520 565196
rect 206428 565156 206434 565168
rect 241514 565156 241520 565168
rect 241572 565156 241578 565208
rect 242894 565156 242900 565208
rect 242952 565196 242958 565208
rect 318150 565196 318156 565208
rect 242952 565168 318156 565196
rect 242952 565156 242958 565168
rect 318150 565156 318156 565168
rect 318208 565156 318214 565208
rect 57698 565088 57704 565140
rect 57756 565128 57762 565140
rect 76834 565128 76840 565140
rect 57756 565100 76840 565128
rect 57756 565088 57762 565100
rect 76834 565088 76840 565100
rect 76892 565088 76898 565140
rect 80330 565088 80336 565140
rect 80388 565128 80394 565140
rect 122006 565128 122012 565140
rect 80388 565100 122012 565128
rect 80388 565088 80394 565100
rect 122006 565088 122012 565100
rect 122064 565088 122070 565140
rect 122098 565088 122104 565140
rect 122156 565128 122162 565140
rect 190546 565128 190552 565140
rect 122156 565100 190552 565128
rect 122156 565088 122162 565100
rect 190546 565088 190552 565100
rect 190604 565088 190610 565140
rect 196342 565088 196348 565140
rect 196400 565128 196406 565140
rect 283098 565128 283104 565140
rect 196400 565100 283104 565128
rect 196400 565088 196406 565100
rect 283098 565088 283104 565100
rect 283156 565088 283162 565140
rect 135254 564884 135260 564936
rect 135312 564924 135318 564936
rect 136174 564924 136180 564936
rect 135312 564896 136180 564924
rect 135312 564884 135318 564896
rect 136174 564884 136180 564896
rect 136232 564884 136238 564936
rect 304258 564340 304264 564392
rect 304316 564380 304322 564392
rect 317966 564380 317972 564392
rect 304316 564352 317972 564380
rect 304316 564340 304322 564352
rect 317966 564340 317972 564352
rect 318024 564340 318030 564392
rect 197814 564000 197820 564052
rect 197872 564040 197878 564052
rect 210694 564040 210700 564052
rect 197872 564012 210700 564040
rect 197872 564000 197878 564012
rect 210694 564000 210700 564012
rect 210752 564000 210758 564052
rect 177758 563932 177764 563984
rect 177816 563972 177822 563984
rect 225138 563972 225144 563984
rect 177816 563944 225144 563972
rect 177816 563932 177822 563944
rect 225138 563932 225144 563944
rect 225196 563932 225202 563984
rect 89622 563864 89628 563916
rect 89680 563904 89686 563916
rect 104894 563904 104900 563916
rect 89680 563876 104900 563904
rect 89680 563864 89686 563876
rect 104894 563864 104900 563876
rect 104952 563864 104958 563916
rect 144086 563864 144092 563916
rect 144144 563904 144150 563916
rect 201678 563904 201684 563916
rect 144144 563876 201684 563904
rect 144144 563864 144150 563876
rect 201678 563864 201684 563876
rect 201736 563864 201742 563916
rect 260190 563864 260196 563916
rect 260248 563904 260254 563916
rect 289170 563904 289176 563916
rect 260248 563876 289176 563904
rect 260248 563864 260254 563876
rect 289170 563864 289176 563876
rect 289228 563864 289234 563916
rect 80974 563796 80980 563848
rect 81032 563836 81038 563848
rect 120994 563836 121000 563848
rect 81032 563808 121000 563836
rect 81032 563796 81038 563808
rect 120994 563796 121000 563808
rect 121052 563796 121058 563848
rect 189166 563796 189172 563848
rect 189224 563836 189230 563848
rect 266998 563836 267004 563848
rect 189224 563808 267004 563836
rect 189224 563796 189230 563808
rect 266998 563796 267004 563808
rect 267056 563796 267062 563848
rect 59538 563728 59544 563780
rect 59596 563768 59602 563780
rect 101030 563768 101036 563780
rect 59596 563740 101036 563768
rect 59596 563728 59602 563740
rect 101030 563728 101036 563740
rect 101088 563728 101094 563780
rect 142246 563728 142252 563780
rect 142304 563768 142310 563780
rect 167730 563768 167736 563780
rect 142304 563740 167736 563768
rect 142304 563728 142310 563740
rect 167730 563728 167736 563740
rect 167788 563728 167794 563780
rect 200666 563728 200672 563780
rect 200724 563768 200730 563780
rect 281810 563768 281816 563780
rect 200724 563740 281816 563768
rect 200724 563728 200730 563740
rect 281810 563728 281816 563740
rect 281868 563728 281874 563780
rect 66714 563660 66720 563712
rect 66772 563700 66778 563712
rect 121178 563700 121184 563712
rect 66772 563672 121184 563700
rect 66772 563660 66778 563672
rect 121178 563660 121184 563672
rect 121236 563660 121242 563712
rect 121546 563660 121552 563712
rect 121604 563700 121610 563712
rect 201126 563700 201132 563712
rect 121604 563672 201132 563700
rect 121604 563660 121610 563672
rect 201126 563660 201132 563672
rect 201184 563660 201190 563712
rect 234338 563660 234344 563712
rect 234396 563700 234402 563712
rect 319714 563700 319720 563712
rect 234396 563672 319720 563700
rect 234396 563660 234402 563672
rect 319714 563660 319720 563672
rect 319772 563660 319778 563712
rect 158714 563388 158720 563440
rect 158772 563428 158778 563440
rect 159818 563428 159824 563440
rect 158772 563400 159824 563428
rect 158772 563388 158778 563400
rect 159818 563388 159824 563400
rect 159876 563388 159882 563440
rect 189902 562572 189908 562624
rect 189960 562612 189966 562624
rect 217318 562612 217324 562624
rect 189960 562584 217324 562612
rect 189960 562572 189966 562584
rect 217318 562572 217324 562584
rect 217376 562572 217382 562624
rect 205726 562504 205732 562556
rect 205784 562544 205790 562556
rect 262858 562544 262864 562556
rect 205784 562516 262864 562544
rect 205784 562504 205790 562516
rect 262858 562504 262864 562516
rect 262916 562504 262922 562556
rect 86034 562436 86040 562488
rect 86092 562476 86098 562488
rect 122190 562476 122196 562488
rect 86092 562448 122196 562476
rect 86092 562436 86098 562448
rect 122190 562436 122196 562448
rect 122248 562436 122254 562488
rect 138474 562436 138480 562488
rect 138532 562476 138538 562488
rect 203242 562476 203248 562488
rect 138532 562448 203248 562476
rect 138532 562436 138538 562448
rect 203242 562436 203248 562448
rect 203300 562436 203306 562488
rect 212166 562436 212172 562488
rect 212224 562476 212230 562488
rect 280890 562476 280896 562488
rect 212224 562448 280896 562476
rect 212224 562436 212230 562448
rect 280890 562436 280896 562448
rect 280948 562436 280954 562488
rect 58526 562368 58532 562420
rect 58584 562408 58590 562420
rect 58584 562380 98316 562408
rect 58584 562368 58590 562380
rect 63126 562300 63132 562352
rect 63184 562340 63190 562352
rect 63184 562312 84194 562340
rect 63184 562300 63190 562312
rect 69014 562232 69020 562284
rect 69072 562272 69078 562284
rect 70302 562272 70308 562284
rect 69072 562244 70308 562272
rect 69072 562232 69078 562244
rect 70302 562232 70308 562244
rect 70360 562232 70366 562284
rect 74534 562232 74540 562284
rect 74592 562272 74598 562284
rect 75270 562272 75276 562284
rect 74592 562244 75276 562272
rect 74592 562232 74598 562244
rect 75270 562232 75276 562244
rect 75328 562232 75334 562284
rect 78674 562232 78680 562284
rect 78732 562272 78738 562284
rect 79594 562272 79600 562284
rect 78732 562244 79600 562272
rect 78732 562232 78738 562244
rect 79594 562232 79600 562244
rect 79652 562232 79658 562284
rect 84166 562204 84194 562312
rect 89806 562300 89812 562352
rect 89864 562340 89870 562352
rect 91002 562340 91008 562352
rect 89864 562312 91008 562340
rect 89864 562300 89870 562312
rect 91002 562300 91008 562312
rect 91060 562300 91066 562352
rect 98288 562340 98316 562380
rect 100754 562368 100760 562420
rect 100812 562408 100818 562420
rect 101766 562408 101772 562420
rect 100812 562380 101772 562408
rect 100812 562368 100818 562380
rect 101766 562368 101772 562380
rect 101824 562368 101830 562420
rect 127618 562368 127624 562420
rect 127676 562408 127682 562420
rect 194594 562408 194600 562420
rect 127676 562380 194600 562408
rect 127676 562368 127682 562380
rect 194594 562368 194600 562380
rect 194652 562368 194658 562420
rect 199194 562368 199200 562420
rect 199252 562408 199258 562420
rect 211798 562408 211804 562420
rect 199252 562380 211804 562408
rect 199252 562368 199258 562380
rect 211798 562368 211804 562380
rect 211856 562368 211862 562420
rect 218146 562368 218152 562420
rect 218204 562408 218210 562420
rect 219250 562408 219256 562420
rect 218204 562380 219256 562408
rect 218204 562368 218210 562380
rect 219250 562368 219256 562380
rect 219308 562368 219314 562420
rect 222194 562368 222200 562420
rect 222252 562408 222258 562420
rect 222838 562408 222844 562420
rect 222252 562380 222844 562408
rect 222252 562368 222258 562380
rect 222838 562368 222844 562380
rect 222896 562368 222902 562420
rect 224954 562368 224960 562420
rect 225012 562408 225018 562420
rect 225782 562408 225788 562420
rect 225012 562380 225788 562408
rect 225012 562368 225018 562380
rect 225782 562368 225788 562380
rect 225840 562368 225846 562420
rect 255314 562368 255320 562420
rect 255372 562408 255378 562420
rect 256510 562408 256516 562420
rect 255372 562380 256516 562408
rect 255372 562368 255378 562380
rect 256510 562368 256516 562380
rect 256568 562368 256574 562420
rect 319622 562408 319628 562420
rect 256712 562380 319628 562408
rect 102502 562340 102508 562352
rect 98288 562312 102508 562340
rect 102502 562300 102508 562312
rect 102560 562300 102566 562352
rect 106274 562300 106280 562352
rect 106332 562340 106338 562352
rect 107562 562340 107568 562352
rect 106332 562312 107568 562340
rect 106332 562300 106338 562312
rect 107562 562300 107568 562312
rect 107620 562300 107626 562352
rect 124214 562300 124220 562352
rect 124272 562340 124278 562352
rect 125410 562340 125416 562352
rect 124272 562312 125416 562340
rect 124272 562300 124278 562312
rect 125410 562300 125416 562312
rect 125468 562300 125474 562352
rect 125594 562300 125600 562352
rect 125652 562340 125658 562352
rect 126882 562340 126888 562352
rect 125652 562312 126888 562340
rect 125652 562300 125658 562312
rect 126882 562300 126888 562312
rect 126940 562300 126946 562352
rect 140774 562300 140780 562352
rect 140832 562340 140838 562352
rect 141878 562340 141884 562352
rect 140832 562312 141884 562340
rect 140832 562300 140838 562312
rect 141878 562300 141884 562312
rect 141936 562300 141942 562352
rect 173158 562340 173164 562352
rect 142126 562312 173164 562340
rect 137462 562232 137468 562284
rect 137520 562272 137526 562284
rect 142126 562272 142154 562312
rect 173158 562300 173164 562312
rect 173216 562300 173222 562352
rect 180794 562300 180800 562352
rect 180852 562340 180858 562352
rect 181990 562340 181996 562352
rect 180852 562312 181996 562340
rect 180852 562300 180858 562312
rect 181990 562300 181996 562312
rect 182048 562300 182054 562352
rect 185578 562300 185584 562352
rect 185636 562340 185642 562352
rect 185636 562312 238754 562340
rect 185636 562300 185642 562312
rect 137520 562244 142154 562272
rect 137520 562232 137526 562244
rect 143534 562232 143540 562284
rect 143592 562272 143598 562284
rect 144730 562272 144736 562284
rect 143592 562244 144736 562272
rect 143592 562232 143598 562244
rect 144730 562232 144736 562244
rect 144788 562232 144794 562284
rect 147674 562232 147680 562284
rect 147732 562272 147738 562284
rect 148318 562272 148324 562284
rect 147732 562244 148324 562272
rect 147732 562232 147738 562244
rect 148318 562232 148324 562244
rect 148376 562232 148382 562284
rect 154574 562232 154580 562284
rect 154632 562272 154638 562284
rect 155494 562272 155500 562284
rect 154632 562244 155500 562272
rect 154632 562232 154638 562244
rect 155494 562232 155500 562244
rect 155552 562232 155558 562284
rect 164326 562232 164332 562284
rect 164384 562272 164390 562284
rect 165522 562272 165528 562284
rect 164384 562244 165528 562272
rect 164384 562232 164390 562244
rect 165522 562232 165528 562244
rect 165580 562232 165586 562284
rect 208394 562232 208400 562284
rect 208452 562272 208458 562284
rect 209222 562272 209228 562284
rect 208452 562244 209228 562272
rect 208452 562232 208458 562244
rect 209222 562232 209228 562244
rect 209280 562232 209286 562284
rect 110506 562204 110512 562216
rect 84166 562176 110512 562204
rect 110506 562164 110512 562176
rect 110564 562164 110570 562216
rect 142154 562164 142160 562216
rect 142212 562204 142218 562216
rect 143350 562204 143356 562216
rect 142212 562176 143356 562204
rect 142212 562164 142218 562176
rect 143350 562164 143356 562176
rect 143408 562164 143414 562216
rect 238726 562204 238754 562312
rect 250806 562232 250812 562284
rect 250864 562272 250870 562284
rect 256712 562272 256740 562380
rect 319622 562368 319628 562380
rect 319680 562368 319686 562420
rect 273254 562300 273260 562352
rect 273312 562340 273318 562352
rect 274450 562340 274456 562352
rect 273312 562312 274456 562340
rect 273312 562300 273318 562312
rect 274450 562300 274456 562312
rect 274508 562300 274514 562352
rect 275186 562300 275192 562352
rect 275244 562340 275250 562352
rect 318058 562340 318064 562352
rect 275244 562312 318064 562340
rect 275244 562300 275250 562312
rect 318058 562300 318064 562312
rect 318116 562300 318122 562352
rect 274634 562272 274640 562284
rect 250864 562244 256740 562272
rect 258046 562244 274640 562272
rect 250864 562232 250870 562244
rect 258046 562204 258074 562244
rect 274634 562232 274640 562244
rect 274692 562232 274698 562284
rect 238726 562176 258074 562204
rect 283742 561824 283748 561876
rect 283800 561864 283806 561876
rect 287790 561864 287796 561876
rect 283800 561836 287796 561864
rect 283800 561824 283806 561836
rect 287790 561824 287796 561836
rect 287848 561824 287854 561876
rect 192110 561212 192116 561264
rect 192168 561252 192174 561264
rect 216030 561252 216036 561264
rect 192168 561224 216036 561252
rect 192168 561212 192174 561224
rect 216030 561212 216036 561224
rect 216088 561212 216094 561264
rect 178494 561144 178500 561196
rect 178552 561184 178558 561196
rect 209038 561184 209044 561196
rect 178552 561156 209044 561184
rect 178552 561144 178558 561156
rect 209038 561144 209044 561156
rect 209096 561144 209102 561196
rect 217870 561144 217876 561196
rect 217928 561184 217934 561196
rect 260098 561184 260104 561196
rect 217928 561156 260104 561184
rect 217928 561144 217934 561156
rect 260098 561144 260104 561156
rect 260156 561144 260162 561196
rect 61378 561076 61384 561128
rect 61436 561116 61442 561128
rect 105354 561116 105360 561128
rect 61436 561088 105360 561116
rect 61436 561076 61442 561088
rect 105354 561076 105360 561088
rect 105412 561076 105418 561128
rect 140498 561076 140504 561128
rect 140556 561116 140562 561128
rect 197998 561116 198004 561128
rect 140556 561088 198004 561116
rect 140556 561076 140562 561088
rect 197998 561076 198004 561088
rect 198056 561076 198062 561128
rect 209130 561076 209136 561128
rect 209188 561116 209194 561128
rect 235994 561116 236000 561128
rect 209188 561088 236000 561116
rect 209188 561076 209194 561088
rect 235994 561076 236000 561088
rect 236052 561076 236058 561128
rect 251542 561076 251548 561128
rect 251600 561116 251606 561128
rect 316862 561116 316868 561128
rect 251600 561088 316868 561116
rect 251600 561076 251606 561088
rect 316862 561076 316868 561088
rect 316920 561076 316926 561128
rect 69566 561008 69572 561060
rect 69624 561048 69630 561060
rect 114646 561048 114652 561060
rect 69624 561020 114652 561048
rect 69624 561008 69630 561020
rect 114646 561008 114652 561020
rect 114704 561008 114710 561060
rect 139486 561008 139492 561060
rect 139544 561048 139550 561060
rect 163406 561048 163412 561060
rect 139544 561020 163412 561048
rect 139544 561008 139550 561020
rect 163406 561008 163412 561020
rect 163464 561008 163470 561060
rect 198550 561008 198556 561060
rect 198608 561048 198614 561060
rect 278038 561048 278044 561060
rect 198608 561020 278044 561048
rect 198608 561008 198614 561020
rect 278038 561008 278044 561020
rect 278096 561008 278102 561060
rect 279510 561008 279516 561060
rect 279568 561048 279574 561060
rect 289078 561048 289084 561060
rect 279568 561020 289084 561048
rect 279568 561008 279574 561020
rect 289078 561008 289084 561020
rect 289136 561008 289142 561060
rect 71682 560940 71688 560992
rect 71740 560980 71746 560992
rect 121730 560980 121736 560992
rect 71740 560952 121736 560980
rect 71740 560940 71746 560952
rect 121730 560940 121736 560952
rect 121788 560940 121794 560992
rect 124030 560940 124036 560992
rect 124088 560980 124094 560992
rect 201862 560980 201868 560992
rect 124088 560952 201868 560980
rect 124088 560940 124094 560952
rect 201862 560940 201868 560952
rect 201920 560940 201926 560992
rect 207106 560940 207112 560992
rect 207164 560980 207170 560992
rect 214558 560980 214564 560992
rect 207164 560952 214564 560980
rect 207164 560940 207170 560952
rect 214558 560940 214564 560952
rect 214616 560940 214622 560992
rect 235074 560940 235080 560992
rect 235132 560980 235138 560992
rect 319530 560980 319536 560992
rect 235132 560952 319536 560980
rect 235132 560940 235138 560952
rect 319530 560940 319536 560952
rect 319588 560940 319594 560992
rect 190454 560804 190460 560856
rect 190512 560844 190518 560856
rect 191374 560844 191380 560856
rect 190512 560816 191380 560844
rect 190512 560804 190518 560816
rect 191374 560804 191380 560816
rect 191432 560804 191438 560856
rect 237926 559852 237932 559904
rect 237984 559892 237990 559904
rect 315482 559892 315488 559904
rect 237984 559864 315488 559892
rect 237984 559852 237990 559864
rect 315482 559852 315488 559864
rect 315540 559852 315546 559904
rect 269482 559784 269488 559836
rect 269540 559824 269546 559836
rect 300118 559824 300124 559836
rect 269540 559796 300124 559824
rect 269540 559784 269546 559796
rect 300118 559784 300124 559796
rect 300176 559784 300182 559836
rect 57514 559716 57520 559768
rect 57572 559756 57578 559768
rect 88242 559756 88248 559768
rect 57572 559728 88248 559756
rect 57572 559716 57578 559728
rect 88242 559716 88248 559728
rect 88300 559716 88306 559768
rect 184934 559716 184940 559768
rect 184992 559756 184998 559768
rect 210602 559756 210608 559768
rect 184992 559728 210608 559756
rect 184992 559716 184998 559728
rect 210602 559716 210608 559728
rect 210660 559716 210666 559768
rect 253658 559716 253664 559768
rect 253716 559756 253722 559768
rect 316770 559756 316776 559768
rect 253716 559728 316776 559756
rect 253716 559716 253722 559728
rect 316770 559716 316776 559728
rect 316828 559716 316834 559768
rect 73154 559648 73160 559700
rect 73212 559688 73218 559700
rect 106918 559688 106924 559700
rect 73212 559660 106924 559688
rect 73212 559648 73218 559660
rect 106918 559648 106924 559660
rect 106976 559648 106982 559700
rect 136910 559648 136916 559700
rect 136968 559688 136974 559700
rect 202230 559688 202236 559700
rect 136968 559660 202236 559688
rect 136968 559648 136974 559660
rect 202230 559648 202236 559660
rect 202288 559648 202294 559700
rect 210694 559648 210700 559700
rect 210752 559688 210758 559700
rect 283190 559688 283196 559700
rect 210752 559660 283196 559688
rect 210752 559648 210758 559660
rect 283190 559648 283196 559660
rect 283248 559648 283254 559700
rect 82446 559580 82452 559632
rect 82504 559620 82510 559632
rect 116578 559620 116584 559632
rect 82504 559592 116584 559620
rect 82504 559580 82510 559592
rect 116578 559580 116584 559592
rect 116636 559580 116642 559632
rect 124674 559580 124680 559632
rect 124732 559620 124738 559632
rect 201218 559620 201224 559632
rect 124732 559592 201224 559620
rect 124732 559580 124738 559592
rect 201218 559580 201224 559592
rect 201276 559580 201282 559632
rect 202138 559580 202144 559632
rect 202196 559620 202202 559632
rect 283466 559620 283472 559632
rect 202196 559592 283472 559620
rect 202196 559580 202202 559592
rect 283466 559580 283472 559592
rect 283524 559580 283530 559632
rect 58710 559512 58716 559564
rect 58768 559552 58774 559564
rect 111058 559552 111064 559564
rect 58768 559524 111064 559552
rect 58768 559512 58774 559524
rect 111058 559512 111064 559524
rect 111116 559512 111122 559564
rect 120442 559512 120448 559564
rect 120500 559552 120506 559564
rect 130378 559552 130384 559564
rect 120500 559524 130384 559552
rect 120500 559512 120506 559524
rect 130378 559512 130384 559524
rect 130436 559512 130442 559564
rect 179138 559512 179144 559564
rect 179196 559552 179202 559564
rect 269758 559552 269764 559564
rect 179196 559524 269764 559552
rect 179196 559512 179202 559524
rect 269758 559512 269764 559524
rect 269816 559512 269822 559564
rect 282362 559512 282368 559564
rect 282420 559552 282426 559564
rect 296070 559552 296076 559564
rect 282420 559524 296076 559552
rect 282420 559512 282426 559524
rect 296070 559512 296076 559524
rect 296128 559512 296134 559564
rect 293770 559444 293776 559496
rect 293828 559484 293834 559496
rect 312722 559484 312728 559496
rect 293828 559456 312728 559484
rect 293828 559444 293834 559456
rect 312722 559444 312728 559456
rect 312780 559444 312786 559496
rect 286686 559376 286692 559428
rect 286744 559416 286750 559428
rect 309778 559416 309784 559428
rect 286744 559388 309784 559416
rect 286744 559376 286750 559388
rect 309778 559376 309784 559388
rect 309836 559376 309842 559428
rect 288066 559308 288072 559360
rect 288124 559348 288130 559360
rect 312538 559348 312544 559360
rect 288124 559320 312544 559348
rect 288124 559308 288130 559320
rect 312538 559308 312544 559320
rect 312596 559308 312602 559360
rect 285214 559240 285220 559292
rect 285272 559280 285278 559292
rect 312814 559280 312820 559292
rect 285272 559252 312820 559280
rect 285272 559240 285278 559252
rect 312814 559240 312820 559252
rect 312872 559240 312878 559292
rect 284938 559172 284944 559224
rect 284996 559212 285002 559224
rect 315298 559212 315304 559224
rect 284996 559184 315304 559212
rect 284996 559172 285002 559184
rect 315298 559172 315304 559184
rect 315356 559172 315362 559224
rect 284478 559104 284484 559156
rect 284536 559144 284542 559156
rect 315574 559144 315580 559156
rect 284536 559116 315580 559144
rect 284536 559104 284542 559116
rect 315574 559104 315580 559116
rect 315632 559104 315638 559156
rect 284202 559036 284208 559088
rect 284260 559076 284266 559088
rect 315390 559076 315396 559088
rect 284260 559048 315396 559076
rect 284260 559036 284266 559048
rect 315390 559036 315396 559048
rect 315448 559036 315454 559088
rect 193214 558968 193220 559020
rect 193272 559008 193278 559020
rect 194226 559008 194232 559020
rect 193272 558980 194232 559008
rect 193272 558968 193278 558980
rect 194226 558968 194232 558980
rect 194284 558968 194290 559020
rect 242250 558968 242256 559020
rect 242308 559008 242314 559020
rect 318242 559008 318248 559020
rect 242308 558980 318248 559008
rect 242308 558968 242314 558980
rect 318242 558968 318248 558980
rect 318300 558968 318306 559020
rect 293126 558900 293132 558952
rect 293184 558940 293190 558952
rect 312906 558940 312912 558952
rect 293184 558912 312912 558940
rect 293184 558900 293190 558912
rect 312906 558900 312912 558912
rect 312964 558900 312970 558952
rect 138934 558288 138940 558340
rect 138992 558328 138998 558340
rect 149790 558328 149796 558340
rect 138992 558300 149796 558328
rect 138992 558288 138998 558300
rect 149790 558288 149796 558300
rect 149848 558288 149854 558340
rect 152642 558288 152648 558340
rect 152700 558328 152706 558340
rect 202874 558328 202880 558340
rect 152700 558300 202880 558328
rect 152700 558288 152706 558300
rect 202874 558288 202880 558300
rect 202932 558288 202938 558340
rect 244366 558288 244372 558340
rect 244424 558328 244430 558340
rect 318058 558328 318064 558340
rect 244424 558300 318064 558328
rect 244424 558288 244430 558300
rect 318058 558288 318064 558300
rect 318116 558288 318122 558340
rect 131206 558220 131212 558272
rect 131264 558260 131270 558272
rect 184198 558260 184204 558272
rect 131264 558232 184204 558260
rect 131264 558220 131270 558232
rect 184198 558220 184204 558232
rect 184256 558220 184262 558272
rect 219158 558220 219164 558272
rect 219216 558260 219222 558272
rect 227162 558260 227168 558272
rect 219216 558232 227168 558260
rect 219216 558220 219222 558232
rect 227162 558220 227168 558232
rect 227220 558220 227226 558272
rect 271598 558220 271604 558272
rect 271656 558260 271662 558272
rect 287698 558260 287704 558272
rect 271656 558232 287704 558260
rect 271656 558220 271662 558232
rect 287698 558220 287704 558232
rect 287756 558220 287762 558272
rect 57422 558152 57428 558204
rect 57480 558192 57486 558204
rect 99190 558192 99196 558204
rect 57480 558164 99196 558192
rect 57480 558152 57486 558164
rect 99190 558152 99196 558164
rect 99248 558152 99254 558204
rect 99282 558152 99288 558204
rect 99340 558192 99346 558204
rect 123110 558192 123116 558204
rect 99340 558164 123116 558192
rect 99340 558152 99346 558164
rect 123110 558152 123116 558164
rect 123168 558152 123174 558204
rect 128262 558152 128268 558204
rect 128320 558192 128326 558204
rect 201034 558192 201040 558204
rect 128320 558164 201040 558192
rect 128320 558152 128326 558164
rect 201034 558152 201040 558164
rect 201092 558152 201098 558204
rect 251174 558192 251180 558204
rect 219406 558164 251180 558192
rect 212810 557948 212816 558000
rect 212868 557988 212874 558000
rect 219406 557988 219434 558164
rect 251174 558152 251180 558164
rect 251232 558152 251238 558204
rect 265894 558152 265900 558204
rect 265952 558192 265958 558204
rect 301498 558192 301504 558204
rect 265952 558164 301504 558192
rect 265952 558152 265958 558164
rect 301498 558152 301504 558164
rect 301556 558152 301562 558204
rect 273070 558084 273076 558136
rect 273128 558124 273134 558136
rect 311158 558124 311164 558136
rect 273128 558096 311164 558124
rect 273128 558084 273134 558096
rect 311158 558084 311164 558096
rect 311216 558084 311222 558136
rect 264422 558016 264428 558068
rect 264480 558056 264486 558068
rect 304350 558056 304356 558068
rect 264480 558028 304356 558056
rect 264480 558016 264486 558028
rect 304350 558016 304356 558028
rect 304408 558016 304414 558068
rect 212868 557960 219434 557988
rect 212868 557948 212874 557960
rect 260834 557948 260840 558000
rect 260892 557988 260898 558000
rect 304258 557988 304264 558000
rect 260892 557960 304264 557988
rect 260892 557948 260898 557960
rect 304258 557948 304264 557960
rect 304316 557948 304322 558000
rect 273714 557880 273720 557932
rect 273772 557920 273778 557932
rect 318150 557920 318156 557932
rect 273772 557892 318156 557920
rect 273772 557880 273778 557892
rect 318150 557880 318156 557892
rect 318208 557880 318214 557932
rect 272334 557812 272340 557864
rect 272392 557852 272398 557864
rect 316678 557852 316684 557864
rect 272392 557824 316684 557852
rect 272392 557812 272398 557824
rect 316678 557812 316684 557824
rect 316736 557812 316742 557864
rect 254394 557744 254400 557796
rect 254452 557784 254458 557796
rect 319622 557784 319628 557796
rect 254452 557756 319628 557784
rect 254452 557744 254458 557756
rect 319622 557744 319628 557756
rect 319680 557744 319686 557796
rect 252278 557676 252284 557728
rect 252336 557716 252342 557728
rect 317966 557716 317972 557728
rect 252336 557688 317972 557716
rect 252336 557676 252342 557688
rect 317966 557676 317972 557688
rect 318024 557676 318030 557728
rect 247218 557608 247224 557660
rect 247276 557648 247282 557660
rect 319530 557648 319536 557660
rect 247276 557620 319536 557648
rect 247276 557608 247282 557620
rect 319530 557608 319536 557620
rect 319588 557608 319594 557660
rect 287330 557540 287336 557592
rect 287388 557580 287394 557592
rect 312630 557580 312636 557592
rect 287388 557552 312636 557580
rect 287388 557540 287394 557552
rect 312630 557540 312636 557552
rect 312688 557540 312694 557592
rect 61654 557472 61660 557524
rect 61712 557512 61718 557524
rect 64874 557512 64880 557524
rect 61712 557484 64880 557512
rect 61712 557472 61718 557484
rect 64874 557472 64880 557484
rect 64932 557472 64938 557524
rect 83458 557472 83464 557524
rect 83516 557512 83522 557524
rect 86770 557512 86776 557524
rect 83516 557484 86776 557512
rect 83516 557472 83522 557484
rect 86770 557472 86776 557484
rect 86828 557472 86834 557524
rect 131850 557472 131856 557524
rect 131908 557512 131914 557524
rect 133138 557512 133144 557524
rect 131908 557484 133144 557512
rect 131908 557472 131914 557484
rect 133138 557472 133144 557484
rect 133196 557472 133202 557524
rect 187786 557472 187792 557524
rect 187844 557512 187850 557524
rect 195238 557512 195244 557524
rect 187844 557484 195244 557512
rect 187844 557472 187850 557484
rect 195238 557472 195244 557484
rect 195296 557472 195302 557524
rect 511350 557472 511356 557524
rect 511408 557512 511414 557524
rect 580166 557512 580172 557524
rect 511408 557484 580172 557512
rect 511408 557472 511414 557484
rect 580166 557472 580172 557484
rect 580224 557472 580230 557524
rect 55122 557404 55128 557456
rect 55180 557444 55186 557456
rect 67358 557444 67364 557456
rect 55180 557416 67364 557444
rect 55180 557404 55186 557416
rect 67358 557404 67364 557416
rect 67416 557404 67422 557456
rect 68370 557404 68376 557456
rect 68428 557444 68434 557456
rect 77386 557444 77392 557456
rect 68428 557416 77392 557444
rect 68428 557404 68434 557416
rect 77386 557404 77392 557416
rect 77444 557404 77450 557456
rect 101398 557404 101404 557456
rect 101456 557444 101462 557456
rect 106090 557444 106096 557456
rect 101456 557416 106096 557444
rect 101456 557404 101462 557416
rect 106090 557404 106096 557416
rect 106148 557404 106154 557456
rect 108390 557404 108396 557456
rect 108448 557444 108454 557456
rect 114646 557444 114652 557456
rect 108448 557416 114652 557444
rect 108448 557404 108454 557416
rect 114646 557404 114652 557416
rect 114704 557404 114710 557456
rect 277302 557404 277308 557456
rect 277360 557444 277366 557456
rect 301682 557444 301688 557456
rect 277360 557416 301688 557444
rect 277360 557404 277366 557416
rect 301682 557404 301688 557416
rect 301740 557404 301746 557456
rect 56502 557336 56508 557388
rect 56560 557376 56566 557388
rect 83918 557376 83924 557388
rect 56560 557348 83924 557376
rect 56560 557336 56566 557348
rect 83918 557336 83924 557348
rect 83976 557336 83982 557388
rect 138750 557336 138756 557388
rect 138808 557376 138814 557388
rect 146938 557376 146944 557388
rect 138808 557348 146944 557376
rect 138808 557336 138814 557348
rect 146938 557336 146944 557348
rect 146996 557336 147002 557388
rect 164878 557336 164884 557388
rect 164936 557376 164942 557388
rect 173434 557376 173440 557388
rect 164936 557348 173440 557376
rect 164936 557336 164942 557348
rect 173434 557336 173440 557348
rect 173492 557336 173498 557388
rect 278038 557336 278044 557388
rect 278096 557376 278102 557388
rect 318610 557376 318616 557388
rect 278096 557348 318616 557376
rect 278096 557336 278102 557348
rect 318610 557336 318616 557348
rect 318668 557336 318674 557388
rect 55030 557268 55036 557320
rect 55088 557308 55094 557320
rect 85298 557308 85304 557320
rect 55088 557280 85304 557308
rect 55088 557268 55094 557280
rect 85298 557268 85304 557280
rect 85356 557268 85362 557320
rect 137830 557268 137836 557320
rect 137888 557308 137894 557320
rect 151262 557308 151268 557320
rect 137888 557280 151268 557308
rect 137888 557268 137894 557280
rect 151262 557268 151268 557280
rect 151320 557268 151326 557320
rect 159358 557268 159364 557320
rect 159416 557308 159422 557320
rect 166994 557308 167000 557320
rect 159416 557280 167000 557308
rect 159416 557268 159422 557280
rect 166994 557268 167000 557280
rect 167052 557268 167058 557320
rect 257246 557268 257252 557320
rect 257304 557308 257310 557320
rect 303062 557308 303068 557320
rect 257304 557280 303068 557308
rect 257304 557268 257310 557280
rect 303062 557268 303068 557280
rect 303120 557268 303126 557320
rect 56410 557200 56416 557252
rect 56468 557240 56474 557252
rect 88886 557240 88892 557252
rect 56468 557212 88892 557240
rect 56468 557200 56474 557212
rect 88886 557200 88892 557212
rect 88944 557200 88950 557252
rect 95326 557240 95332 557252
rect 93826 557212 95332 557240
rect 60366 557132 60372 557184
rect 60424 557172 60430 557184
rect 93826 557172 93854 557212
rect 95326 557200 95332 557212
rect 95384 557200 95390 557252
rect 139854 557200 139860 557252
rect 139912 557240 139918 557252
rect 153378 557240 153384 557252
rect 139912 557212 153384 557240
rect 139912 557200 139918 557212
rect 153378 557200 153384 557212
rect 153436 557200 153442 557252
rect 164142 557200 164148 557252
rect 164200 557240 164206 557252
rect 171778 557240 171784 557252
rect 164200 557212 171784 557240
rect 164200 557200 164206 557212
rect 171778 557200 171784 557212
rect 171836 557200 171842 557252
rect 252922 557200 252928 557252
rect 252980 557240 252986 557252
rect 319346 557240 319352 557252
rect 252980 557212 319352 557240
rect 252980 557200 252986 557212
rect 319346 557200 319352 557212
rect 319404 557200 319410 557252
rect 60424 557144 93854 557172
rect 60424 557132 60430 557144
rect 114002 557132 114008 557184
rect 114060 557172 114066 557184
rect 124306 557172 124312 557184
rect 114060 557144 124312 557172
rect 114060 557132 114066 557144
rect 124306 557132 124312 557144
rect 124364 557132 124370 557184
rect 135162 557132 135168 557184
rect 135220 557172 135226 557184
rect 156966 557172 156972 557184
rect 135220 557144 156972 557172
rect 135220 557132 135226 557144
rect 156966 557132 156972 557144
rect 157024 557132 157030 557184
rect 160738 557132 160744 557184
rect 160796 557172 160802 557184
rect 172698 557172 172704 557184
rect 160796 557144 172704 557172
rect 160796 557132 160802 557144
rect 172698 557132 172704 557144
rect 172756 557132 172762 557184
rect 255866 557132 255872 557184
rect 255924 557172 255930 557184
rect 301774 557172 301780 557184
rect 255924 557144 301780 557172
rect 255924 557132 255930 557144
rect 301774 557132 301780 557144
rect 301832 557132 301838 557184
rect 54938 557064 54944 557116
rect 54996 557104 55002 557116
rect 93026 557104 93032 557116
rect 54996 557076 93032 557104
rect 54996 557064 55002 557076
rect 93026 557064 93032 557076
rect 93084 557064 93090 557116
rect 93118 557064 93124 557116
rect 93176 557104 93182 557116
rect 96798 557104 96804 557116
rect 93176 557076 96804 557104
rect 93176 557064 93182 557076
rect 96798 557064 96804 557076
rect 96856 557064 96862 557116
rect 99190 557064 99196 557116
rect 99248 557104 99254 557116
rect 116854 557104 116860 557116
rect 99248 557076 116860 557104
rect 99248 557064 99254 557076
rect 116854 557064 116860 557076
rect 116912 557064 116918 557116
rect 118234 557064 118240 557116
rect 118292 557104 118298 557116
rect 126238 557104 126244 557116
rect 118292 557076 126244 557104
rect 118292 557064 118298 557076
rect 126238 557064 126244 557076
rect 126296 557064 126302 557116
rect 135070 557064 135076 557116
rect 135128 557104 135134 557116
rect 164878 557104 164884 557116
rect 135128 557076 164884 557104
rect 135128 557064 135134 557076
rect 164878 557064 164884 557076
rect 164936 557064 164942 557116
rect 171962 557104 171968 557116
rect 171106 557076 171968 557104
rect 58618 556996 58624 557048
rect 58676 557036 58682 557048
rect 68370 557036 68376 557048
rect 58676 557008 68376 557036
rect 58676 556996 58682 557008
rect 68370 556996 68376 557008
rect 68428 556996 68434 557048
rect 68462 556996 68468 557048
rect 68520 557036 68526 557048
rect 99650 557036 99656 557048
rect 68520 557008 99656 557036
rect 68520 556996 68526 557008
rect 99650 556996 99656 557008
rect 99708 556996 99714 557048
rect 106826 556996 106832 557048
rect 106884 557036 106890 557048
rect 121638 557036 121644 557048
rect 106884 557008 121644 557036
rect 106884 556996 106890 557008
rect 121638 556996 121644 557008
rect 121696 556996 121702 557048
rect 136542 556996 136548 557048
rect 136600 557036 136606 557048
rect 171106 557036 171134 557076
rect 171962 557064 171968 557076
rect 172020 557064 172026 557116
rect 176286 557064 176292 557116
rect 176344 557104 176350 557116
rect 210510 557104 210516 557116
rect 176344 557076 210516 557104
rect 176344 557064 176350 557076
rect 210510 557064 210516 557076
rect 210568 557064 210574 557116
rect 261570 557064 261576 557116
rect 261628 557104 261634 557116
rect 282178 557104 282184 557116
rect 261628 557076 282184 557104
rect 261628 557064 261634 557076
rect 282178 557064 282184 557076
rect 282236 557064 282242 557116
rect 136600 557008 171134 557036
rect 136600 556996 136606 557008
rect 171318 556996 171324 557048
rect 171376 557036 171382 557048
rect 188338 557036 188344 557048
rect 171376 557008 188344 557036
rect 171376 556996 171382 557008
rect 188338 556996 188344 557008
rect 188396 556996 188402 557048
rect 199930 556996 199936 557048
rect 199988 557036 199994 557048
rect 210418 557036 210424 557048
rect 199988 557008 210424 557036
rect 199988 556996 199994 557008
rect 210418 556996 210424 557008
rect 210476 556996 210482 557048
rect 217962 556996 217968 557048
rect 218020 557036 218026 557048
rect 218606 557036 218612 557048
rect 218020 557008 218612 557036
rect 218020 556996 218026 557008
rect 218606 556996 218612 557008
rect 218664 556996 218670 557048
rect 245838 556996 245844 557048
rect 245896 557036 245902 557048
rect 281074 557036 281080 557048
rect 245896 557008 281080 557036
rect 245896 556996 245902 557008
rect 281074 556996 281080 557008
rect 281132 556996 281138 557048
rect 63218 556928 63224 556980
rect 63276 556968 63282 556980
rect 76006 556968 76012 556980
rect 63276 556940 76012 556968
rect 63276 556928 63282 556940
rect 76006 556928 76012 556940
rect 76064 556928 76070 556980
rect 76834 556928 76840 556980
rect 76892 556968 76898 556980
rect 117590 556968 117596 556980
rect 76892 556940 117596 556968
rect 76892 556928 76898 556940
rect 117590 556928 117596 556940
rect 117648 556928 117654 556980
rect 118970 556928 118976 556980
rect 119028 556968 119034 556980
rect 134518 556968 134524 556980
rect 119028 556940 134524 556968
rect 119028 556928 119034 556940
rect 134518 556928 134524 556940
rect 134576 556928 134582 556980
rect 137738 556928 137744 556980
rect 137796 556968 137802 556980
rect 175550 556968 175556 556980
rect 137796 556940 175556 556968
rect 137796 556928 137802 556940
rect 175550 556928 175556 556940
rect 175608 556928 175614 556980
rect 195606 556928 195612 556980
rect 195664 556968 195670 556980
rect 206462 556968 206468 556980
rect 195664 556940 206468 556968
rect 195664 556928 195670 556940
rect 206462 556928 206468 556940
rect 206520 556928 206526 556980
rect 218054 556928 218060 556980
rect 218112 556968 218118 556980
rect 230014 556968 230020 556980
rect 218112 556940 230020 556968
rect 218112 556928 218118 556940
rect 230014 556928 230020 556940
rect 230072 556928 230078 556980
rect 231486 556928 231492 556980
rect 231544 556968 231550 556980
rect 238754 556968 238760 556980
rect 231544 556940 238760 556968
rect 231544 556928 231550 556940
rect 238754 556928 238760 556940
rect 238812 556928 238818 556980
rect 239398 556928 239404 556980
rect 239456 556968 239462 556980
rect 280982 556968 280988 556980
rect 239456 556940 280988 556968
rect 239456 556928 239462 556940
rect 280982 556928 280988 556940
rect 281040 556928 281046 556980
rect 56318 556860 56324 556912
rect 56376 556900 56382 556912
rect 98914 556900 98920 556912
rect 56376 556872 98920 556900
rect 56376 556860 56382 556872
rect 98914 556860 98920 556872
rect 98972 556860 98978 556912
rect 103974 556860 103980 556912
rect 104032 556900 104038 556912
rect 124398 556900 124404 556912
rect 104032 556872 124404 556900
rect 104032 556860 104038 556872
rect 124398 556860 124404 556872
rect 124456 556860 124462 556912
rect 136450 556860 136456 556912
rect 136508 556900 136514 556912
rect 157702 556900 157708 556912
rect 136508 556872 157708 556900
rect 136508 556860 136514 556872
rect 157702 556860 157708 556872
rect 157760 556860 157766 556912
rect 158346 556860 158352 556912
rect 158404 556900 158410 556912
rect 200942 556900 200948 556912
rect 158404 556872 200948 556900
rect 158404 556860 158410 556872
rect 200942 556860 200948 556872
rect 201000 556860 201006 556912
rect 220078 556860 220084 556912
rect 220136 556900 220142 556912
rect 232866 556900 232872 556912
rect 220136 556872 232872 556900
rect 220136 556860 220142 556872
rect 232866 556860 232872 556872
rect 232924 556860 232930 556912
rect 238662 556860 238668 556912
rect 238720 556900 238726 556912
rect 284938 556900 284944 556912
rect 238720 556872 284944 556900
rect 238720 556860 238726 556872
rect 284938 556860 284944 556872
rect 284996 556860 285002 556912
rect 57790 556792 57796 556844
rect 57848 556832 57854 556844
rect 73798 556832 73804 556844
rect 57848 556804 73804 556832
rect 57848 556792 57854 556804
rect 73798 556792 73804 556804
rect 73856 556792 73862 556844
rect 78122 556792 78128 556844
rect 78180 556832 78186 556844
rect 120810 556832 120816 556844
rect 78180 556804 120816 556832
rect 78180 556792 78186 556804
rect 120810 556792 120816 556804
rect 120868 556792 120874 556844
rect 146202 556792 146208 556844
rect 146260 556832 146266 556844
rect 201494 556832 201500 556844
rect 146260 556804 201500 556832
rect 146260 556792 146266 556804
rect 201494 556792 201500 556804
rect 201552 556792 201558 556844
rect 204990 556792 204996 556844
rect 205048 556832 205054 556844
rect 213178 556832 213184 556844
rect 205048 556804 213184 556832
rect 205048 556792 205054 556804
rect 213178 556792 213184 556804
rect 213236 556792 213242 556844
rect 218698 556792 218704 556844
rect 218756 556832 218762 556844
rect 233602 556832 233608 556844
rect 218756 556804 233608 556832
rect 218756 556792 218762 556804
rect 233602 556792 233608 556804
rect 233660 556792 233666 556844
rect 237190 556792 237196 556844
rect 237248 556832 237254 556844
rect 284202 556832 284208 556844
rect 237248 556804 284208 556832
rect 237248 556792 237254 556804
rect 284202 556792 284208 556804
rect 284260 556792 284266 556844
rect 299566 556792 299572 556844
rect 299624 556832 299630 556844
rect 319438 556832 319444 556844
rect 299624 556804 319444 556832
rect 299624 556792 299630 556804
rect 319438 556792 319444 556804
rect 319496 556792 319502 556844
rect 59170 556724 59176 556776
rect 59228 556764 59234 556776
rect 68462 556764 68468 556776
rect 59228 556736 68468 556764
rect 59228 556724 59234 556736
rect 68462 556724 68468 556736
rect 68520 556724 68526 556776
rect 105538 556724 105544 556776
rect 105596 556764 105602 556776
rect 108942 556764 108948 556776
rect 105596 556736 108948 556764
rect 105596 556724 105602 556736
rect 108942 556724 108948 556736
rect 109000 556724 109006 556776
rect 275922 556724 275928 556776
rect 275980 556764 275986 556776
rect 300394 556764 300400 556776
rect 275980 556736 300400 556764
rect 275980 556724 275986 556736
rect 300394 556724 300400 556736
rect 300452 556724 300458 556776
rect 270862 556656 270868 556708
rect 270920 556696 270926 556708
rect 300210 556696 300216 556708
rect 270920 556668 300216 556696
rect 270920 556656 270926 556668
rect 300210 556656 300216 556668
rect 300268 556656 300274 556708
rect 285950 556588 285956 556640
rect 286008 556628 286014 556640
rect 319714 556628 319720 556640
rect 286008 556600 319720 556628
rect 286008 556588 286014 556600
rect 319714 556588 319720 556600
rect 319772 556588 319778 556640
rect 280154 556520 280160 556572
rect 280212 556560 280218 556572
rect 316862 556560 316868 556572
rect 280212 556532 316868 556560
rect 280212 556520 280218 556532
rect 316862 556520 316868 556532
rect 316920 556520 316926 556572
rect 88978 556452 88984 556504
rect 89036 556492 89042 556504
rect 90358 556492 90364 556504
rect 89036 556464 90364 556492
rect 89036 556452 89042 556464
rect 90358 556452 90364 556464
rect 90416 556452 90422 556504
rect 262306 556452 262312 556504
rect 262364 556492 262370 556504
rect 300302 556492 300308 556504
rect 262364 556464 300308 556492
rect 262364 556452 262370 556464
rect 300302 556452 300308 556464
rect 300360 556452 300366 556504
rect 173158 556384 173164 556436
rect 173216 556424 173222 556436
rect 174906 556424 174912 556436
rect 173216 556396 174912 556424
rect 173216 556384 173222 556396
rect 174906 556384 174912 556396
rect 174964 556384 174970 556436
rect 240042 556384 240048 556436
rect 240100 556424 240106 556436
rect 266354 556424 266360 556436
rect 240100 556396 266360 556424
rect 240100 556384 240106 556396
rect 266354 556384 266360 556396
rect 266412 556384 266418 556436
rect 281626 556384 281632 556436
rect 281684 556424 281690 556436
rect 300118 556424 300124 556436
rect 281684 556396 300124 556424
rect 281684 556384 281690 556396
rect 300118 556384 300124 556396
rect 300176 556384 300182 556436
rect 101490 556316 101496 556368
rect 101548 556356 101554 556368
rect 103238 556356 103244 556368
rect 101548 556328 103244 556356
rect 101548 556316 101554 556328
rect 103238 556316 103244 556328
rect 103296 556316 103302 556368
rect 108298 556316 108304 556368
rect 108356 556356 108362 556368
rect 111794 556356 111800 556368
rect 108356 556328 111800 556356
rect 108356 556316 108362 556328
rect 111794 556316 111800 556328
rect 111852 556316 111858 556368
rect 202782 556316 202788 556368
rect 202840 556356 202846 556368
rect 209130 556356 209136 556368
rect 202840 556328 209136 556356
rect 202840 556316 202846 556328
rect 209130 556316 209136 556328
rect 209188 556316 209194 556368
rect 283098 556316 283104 556368
rect 283156 556356 283162 556368
rect 301590 556356 301596 556368
rect 283156 556328 301596 556356
rect 283156 556316 283162 556328
rect 301590 556316 301596 556328
rect 301648 556316 301654 556368
rect 88242 556248 88248 556300
rect 88300 556288 88306 556300
rect 91738 556288 91744 556300
rect 88300 556260 91744 556288
rect 88300 556248 88306 556260
rect 91738 556248 91744 556260
rect 91796 556248 91802 556300
rect 137646 556248 137652 556300
rect 137704 556288 137710 556300
rect 138658 556288 138664 556300
rect 137704 556260 138664 556288
rect 137704 556248 137710 556260
rect 138658 556248 138664 556260
rect 138716 556248 138722 556300
rect 162670 556248 162676 556300
rect 162728 556288 162734 556300
rect 168374 556288 168380 556300
rect 162728 556260 168380 556288
rect 162728 556248 162734 556260
rect 168374 556248 168380 556260
rect 168432 556248 168438 556300
rect 174170 556248 174176 556300
rect 174228 556288 174234 556300
rect 179506 556288 179512 556300
rect 174228 556260 179512 556288
rect 174228 556248 174234 556260
rect 179506 556248 179512 556260
rect 179564 556248 179570 556300
rect 201402 556248 201408 556300
rect 201460 556288 201466 556300
rect 206278 556288 206284 556300
rect 201460 556260 206284 556288
rect 201460 556248 201466 556260
rect 206278 556248 206284 556260
rect 206336 556248 206342 556300
rect 209958 556248 209964 556300
rect 210016 556288 210022 556300
rect 215938 556288 215944 556300
rect 210016 556260 215944 556288
rect 210016 556248 210022 556260
rect 215938 556248 215944 556260
rect 215996 556248 216002 556300
rect 293954 556248 293960 556300
rect 294012 556288 294018 556300
rect 295242 556288 295248 556300
rect 294012 556260 295248 556288
rect 294012 556248 294018 556260
rect 295242 556248 295248 556260
rect 295300 556248 295306 556300
rect 296714 556248 296720 556300
rect 296772 556288 296778 556300
rect 297358 556288 297364 556300
rect 296772 556260 297364 556288
rect 296772 556248 296778 556260
rect 297358 556248 297364 556260
rect 297416 556248 297422 556300
rect 298094 556248 298100 556300
rect 298152 556288 298158 556300
rect 316770 556288 316776 556300
rect 298152 556260 316776 556288
rect 298152 556248 298158 556260
rect 316770 556248 316776 556260
rect 316828 556248 316834 556300
rect 96062 556180 96068 556232
rect 96120 556220 96126 556232
rect 99282 556220 99288 556232
rect 96120 556192 99288 556220
rect 96120 556180 96126 556192
rect 99282 556180 99288 556192
rect 99340 556180 99346 556232
rect 115474 556180 115480 556232
rect 115532 556220 115538 556232
rect 116118 556220 116124 556232
rect 115532 556192 116124 556220
rect 115532 556180 115538 556192
rect 116118 556180 116124 556192
rect 116176 556180 116182 556232
rect 121086 556180 121092 556232
rect 121144 556220 121150 556232
rect 122098 556220 122104 556232
rect 121144 556192 122104 556220
rect 121144 556180 121150 556192
rect 122098 556180 122104 556192
rect 122156 556180 122162 556232
rect 154114 556180 154120 556232
rect 154172 556220 154178 556232
rect 157978 556220 157984 556232
rect 154172 556192 157984 556220
rect 154172 556180 154178 556192
rect 157978 556180 157984 556192
rect 158036 556180 158042 556232
rect 167822 556180 167828 556232
rect 167880 556220 167886 556232
rect 169846 556220 169852 556232
rect 167880 556192 169852 556220
rect 167880 556180 167886 556192
rect 169846 556180 169852 556192
rect 169904 556180 169910 556232
rect 203518 556180 203524 556232
rect 203576 556220 203582 556232
rect 204898 556220 204904 556232
rect 203576 556192 204904 556220
rect 203576 556180 203582 556192
rect 204898 556180 204904 556192
rect 204956 556180 204962 556232
rect 276566 556180 276572 556232
rect 276624 556220 276630 556232
rect 301866 556220 301872 556232
rect 276624 556192 301872 556220
rect 276624 556180 276630 556192
rect 301866 556180 301872 556192
rect 301924 556180 301930 556232
rect 295978 555704 295984 555756
rect 296036 555744 296042 555756
rect 313090 555744 313096 555756
rect 296036 555716 313096 555744
rect 296036 555704 296042 555716
rect 313090 555704 313096 555716
rect 313148 555704 313154 555756
rect 294506 555636 294512 555688
rect 294564 555676 294570 555688
rect 315666 555676 315672 555688
rect 294564 555648 315672 555676
rect 294564 555636 294570 555648
rect 315666 555636 315672 555648
rect 315724 555636 315730 555688
rect 278774 555568 278780 555620
rect 278832 555608 278838 555620
rect 300762 555608 300768 555620
rect 278832 555580 300768 555608
rect 278832 555568 278838 555580
rect 300762 555568 300768 555580
rect 300820 555568 300826 555620
rect 268746 555500 268752 555552
rect 268804 555540 268810 555552
rect 302878 555540 302884 555552
rect 268804 555512 302884 555540
rect 268804 555500 268810 555512
rect 302878 555500 302884 555512
rect 302936 555500 302942 555552
rect 266354 555432 266360 555484
rect 266412 555472 266418 555484
rect 318702 555472 318708 555484
rect 266412 555444 318708 555472
rect 266412 555432 266418 555444
rect 318702 555432 318708 555444
rect 318760 555432 318766 555484
rect 263042 555364 263048 555416
rect 263100 555404 263106 555416
rect 301958 555404 301964 555416
rect 263100 555376 301964 555404
rect 263100 555364 263106 555376
rect 301958 555364 301964 555376
rect 302016 555364 302022 555416
rect 265158 555296 265164 555348
rect 265216 555336 265222 555348
rect 312998 555336 313004 555348
rect 265216 555308 313004 555336
rect 265216 555296 265222 555308
rect 312998 555296 313004 555308
rect 313056 555296 313062 555348
rect 243630 555228 243636 555280
rect 243688 555268 243694 555280
rect 305730 555268 305736 555280
rect 243688 555240 305736 555268
rect 243688 555228 243694 555240
rect 305730 555228 305736 555240
rect 305788 555228 305794 555280
rect 236470 555160 236476 555212
rect 236528 555200 236534 555212
rect 301406 555200 301412 555212
rect 236528 555172 301412 555200
rect 236528 555160 236534 555172
rect 301406 555160 301412 555172
rect 301464 555160 301470 555212
rect 249442 555092 249448 555144
rect 249500 555132 249506 555144
rect 318426 555132 318432 555144
rect 249500 555104 318432 555132
rect 249500 555092 249506 555104
rect 318426 555092 318432 555104
rect 318484 555092 318490 555144
rect 235902 555024 235908 555076
rect 235960 555064 235966 555076
rect 319438 555064 319444 555076
rect 235960 555036 319444 555064
rect 235960 555024 235966 555036
rect 319438 555024 319444 555036
rect 319496 555024 319502 555076
rect 300762 554684 300768 554736
rect 300820 554724 300826 554736
rect 317966 554724 317972 554736
rect 300820 554696 317972 554724
rect 300820 554684 300826 554696
rect 317966 554684 317972 554696
rect 318024 554684 318030 554736
rect 301406 550536 301412 550588
rect 301464 550576 301470 550588
rect 317414 550576 317420 550588
rect 301464 550548 317420 550576
rect 301464 550536 301470 550548
rect 317414 550536 317420 550548
rect 317472 550536 317478 550588
rect 305730 545028 305736 545080
rect 305788 545068 305794 545080
rect 317966 545068 317972 545080
rect 305788 545040 317972 545068
rect 305788 545028 305794 545040
rect 317966 545028 317972 545040
rect 318024 545028 318030 545080
rect 430942 543192 430948 543244
rect 431000 543232 431006 543244
rect 431402 543232 431408 543244
rect 431000 543204 431408 543232
rect 431000 543192 431006 543204
rect 431402 543192 431408 543204
rect 431460 543192 431466 543244
rect 430758 543056 430764 543108
rect 430816 543096 430822 543108
rect 430942 543096 430948 543108
rect 430816 543068 430948 543096
rect 430816 543056 430822 543068
rect 430942 543056 430948 543068
rect 431000 543056 431006 543108
rect 319254 542988 319260 543040
rect 319312 543028 319318 543040
rect 319438 543028 319444 543040
rect 319312 543000 319444 543028
rect 319312 542988 319318 543000
rect 319438 542988 319444 543000
rect 319496 542988 319502 543040
rect 319162 536256 319168 536308
rect 319220 536296 319226 536308
rect 319530 536296 319536 536308
rect 319220 536268 319536 536296
rect 319220 536256 319226 536268
rect 319530 536256 319536 536268
rect 319588 536256 319594 536308
rect 312906 535372 312912 535424
rect 312964 535412 312970 535424
rect 512178 535412 512184 535424
rect 312964 535384 512184 535412
rect 312964 535372 312970 535384
rect 512178 535372 512184 535384
rect 512236 535372 512242 535424
rect 313090 535304 313096 535356
rect 313148 535344 313154 535356
rect 505094 535344 505100 535356
rect 313148 535316 505100 535344
rect 313148 535304 313154 535316
rect 505094 535304 505100 535316
rect 505152 535304 505158 535356
rect 312814 535236 312820 535288
rect 312872 535276 312878 535288
rect 466454 535276 466460 535288
rect 312872 535248 466460 535276
rect 312872 535236 312878 535248
rect 466454 535236 466460 535248
rect 466512 535236 466518 535288
rect 300486 535168 300492 535220
rect 300544 535208 300550 535220
rect 430666 535208 430672 535220
rect 300544 535180 430672 535208
rect 300544 535168 300550 535180
rect 430666 535168 430672 535180
rect 430724 535168 430730 535220
rect 300670 535100 300676 535152
rect 300728 535140 300734 535152
rect 430758 535140 430764 535152
rect 300728 535112 430764 535140
rect 300728 535100 300734 535112
rect 430758 535100 430764 535112
rect 430816 535100 430822 535152
rect 303062 535032 303068 535084
rect 303120 535072 303126 535084
rect 431310 535072 431316 535084
rect 303120 535044 431316 535072
rect 303120 535032 303126 535044
rect 431310 535032 431316 535044
rect 431368 535032 431374 535084
rect 315574 534964 315580 535016
rect 315632 535004 315638 535016
rect 429470 535004 429476 535016
rect 315632 534976 429476 535004
rect 315632 534964 315638 534976
rect 429470 534964 429476 534976
rect 429528 534964 429534 535016
rect 316862 534896 316868 534948
rect 316920 534936 316926 534948
rect 430574 534936 430580 534948
rect 316920 534908 430580 534936
rect 316920 534896 316926 534908
rect 430574 534896 430580 534908
rect 430632 534896 430638 534948
rect 318610 534828 318616 534880
rect 318668 534868 318674 534880
rect 431218 534868 431224 534880
rect 318668 534840 431224 534868
rect 318668 534828 318674 534840
rect 431218 534828 431224 534840
rect 431276 534828 431282 534880
rect 319346 534760 319352 534812
rect 319404 534800 319410 534812
rect 431126 534800 431132 534812
rect 319404 534772 431132 534800
rect 319404 534760 319410 534772
rect 431126 534760 431132 534772
rect 431184 534760 431190 534812
rect 318242 534692 318248 534744
rect 318300 534732 318306 534744
rect 428458 534732 428464 534744
rect 318300 534704 428464 534732
rect 318300 534692 318306 534704
rect 428458 534692 428464 534704
rect 428516 534692 428522 534744
rect 300394 534148 300400 534200
rect 300452 534188 300458 534200
rect 351270 534188 351276 534200
rect 300452 534160 351276 534188
rect 300452 534148 300458 534160
rect 351270 534148 351276 534160
rect 351328 534148 351334 534200
rect 305638 534080 305644 534132
rect 305696 534120 305702 534132
rect 369302 534120 369308 534132
rect 305696 534092 369308 534120
rect 305696 534080 305702 534092
rect 369302 534080 369308 534092
rect 369360 534080 369366 534132
rect 309778 534012 309784 534064
rect 309836 534052 309842 534064
rect 512086 534052 512092 534064
rect 309836 534024 512092 534052
rect 309836 534012 309842 534024
rect 512086 534012 512092 534024
rect 512144 534012 512150 534064
rect 318334 533944 318340 533996
rect 318392 533984 318398 533996
rect 489914 533984 489920 533996
rect 318392 533956 489920 533984
rect 318392 533944 318398 533956
rect 489914 533944 489920 533956
rect 489972 533944 489978 533996
rect 319530 533876 319536 533928
rect 319588 533916 319594 533928
rect 483014 533916 483020 533928
rect 319588 533888 483020 533916
rect 319588 533876 319594 533888
rect 483014 533876 483020 533888
rect 483072 533876 483078 533928
rect 302970 533808 302976 533860
rect 303028 533848 303034 533860
rect 457622 533848 457628 533860
rect 303028 533820 457628 533848
rect 303028 533808 303034 533820
rect 457622 533808 457628 533820
rect 457680 533808 457686 533860
rect 312722 533740 312728 533792
rect 312780 533780 312786 533792
rect 459554 533780 459560 533792
rect 312780 533752 459560 533780
rect 312780 533740 312786 533752
rect 459554 533740 459560 533752
rect 459612 533740 459618 533792
rect 315666 533672 315672 533724
rect 315724 533712 315730 533724
rect 457530 533712 457536 533724
rect 315724 533684 457536 533712
rect 315724 533672 315730 533684
rect 457530 533672 457536 533684
rect 457588 533672 457594 533724
rect 316770 533604 316776 533656
rect 316828 533644 316834 533656
rect 457438 533644 457444 533656
rect 316828 533616 457444 533644
rect 316828 533604 316834 533616
rect 457438 533604 457444 533616
rect 457496 533604 457502 533656
rect 300118 533536 300124 533588
rect 300176 533576 300182 533588
rect 431034 533576 431040 533588
rect 300176 533548 431040 533576
rect 300176 533536 300182 533548
rect 431034 533536 431040 533548
rect 431092 533536 431098 533588
rect 300210 533468 300216 533520
rect 300268 533508 300274 533520
rect 430850 533508 430856 533520
rect 300268 533480 430856 533508
rect 300268 533468 300274 533480
rect 430850 533468 430856 533480
rect 430908 533468 430914 533520
rect 301682 533400 301688 533452
rect 301740 533440 301746 533452
rect 431402 533440 431408 533452
rect 301740 533412 431408 533440
rect 301740 533400 301746 533412
rect 431402 533400 431408 533412
rect 431460 533400 431466 533452
rect 301590 533332 301596 533384
rect 301648 533372 301654 533384
rect 430942 533372 430948 533384
rect 301648 533344 430948 533372
rect 301648 533332 301654 533344
rect 430942 533332 430948 533344
rect 431000 533332 431006 533384
rect 301866 533264 301872 533316
rect 301924 533304 301930 533316
rect 414934 533304 414940 533316
rect 301924 533276 414940 533304
rect 301924 533264 301930 533276
rect 414934 533264 414940 533276
rect 414992 533264 414998 533316
rect 301774 533196 301780 533248
rect 301832 533236 301838 533248
rect 405918 533236 405924 533248
rect 301832 533208 405924 533236
rect 301832 533196 301838 533208
rect 405918 533196 405924 533208
rect 405976 533196 405982 533248
rect 300302 533128 300308 533180
rect 300360 533168 300366 533180
rect 328638 533168 328644 533180
rect 300360 533140 328644 533168
rect 300360 533128 300366 533140
rect 328638 533128 328644 533140
rect 328696 533128 328702 533180
rect 304258 532652 304264 532704
rect 304316 532692 304322 532704
rect 342254 532692 342260 532704
rect 304316 532664 342260 532692
rect 304316 532652 304322 532664
rect 342254 532652 342260 532664
rect 342312 532652 342318 532704
rect 312998 532584 313004 532636
rect 313056 532624 313062 532636
rect 319622 532624 319628 532636
rect 313056 532596 319628 532624
rect 313056 532584 313062 532596
rect 319622 532584 319628 532596
rect 319680 532584 319686 532636
rect 346670 532624 346676 532636
rect 319732 532596 346676 532624
rect 319438 532516 319444 532568
rect 319496 532556 319502 532568
rect 319732 532556 319760 532596
rect 346670 532584 346676 532596
rect 346728 532584 346734 532636
rect 333238 532556 333244 532568
rect 319496 532528 319760 532556
rect 319824 532528 333244 532556
rect 319496 532516 319502 532528
rect 319254 532448 319260 532500
rect 319312 532488 319318 532500
rect 319824 532488 319852 532528
rect 333238 532516 333244 532528
rect 333296 532516 333302 532568
rect 319312 532460 319852 532488
rect 319312 532448 319318 532460
rect 319898 532448 319904 532500
rect 319956 532488 319962 532500
rect 410518 532488 410524 532500
rect 319956 532460 410524 532488
rect 319956 532448 319962 532460
rect 410518 532448 410524 532460
rect 410576 532448 410582 532500
rect 302878 532380 302884 532432
rect 302936 532420 302942 532432
rect 387886 532420 387892 532432
rect 302936 532392 387892 532420
rect 302936 532380 302942 532392
rect 387886 532380 387892 532392
rect 387944 532380 387950 532432
rect 301498 532312 301504 532364
rect 301556 532352 301562 532364
rect 383654 532352 383660 532364
rect 301556 532324 383660 532352
rect 301556 532312 301562 532324
rect 383654 532312 383660 532324
rect 383712 532312 383718 532364
rect 318150 532244 318156 532296
rect 318208 532284 318214 532296
rect 396902 532284 396908 532296
rect 318208 532256 396908 532284
rect 318208 532244 318214 532256
rect 396902 532244 396908 532256
rect 396960 532244 396966 532296
rect 304350 532176 304356 532228
rect 304408 532216 304414 532228
rect 374454 532216 374460 532228
rect 304408 532188 374460 532216
rect 304408 532176 304414 532188
rect 374454 532176 374460 532188
rect 374512 532176 374518 532228
rect 311158 532108 311164 532160
rect 311216 532148 311222 532160
rect 364702 532148 364708 532160
rect 311216 532120 364708 532148
rect 311216 532108 311222 532120
rect 364702 532108 364708 532120
rect 364760 532108 364766 532160
rect 319162 532040 319168 532092
rect 319220 532080 319226 532092
rect 360286 532080 360292 532092
rect 319220 532052 360292 532080
rect 319220 532040 319226 532052
rect 360286 532040 360292 532052
rect 360344 532040 360350 532092
rect 318518 531972 318524 532024
rect 318576 532012 318582 532024
rect 356238 532012 356244 532024
rect 318576 531984 356244 532012
rect 318576 531972 318582 531984
rect 356238 531972 356244 531984
rect 356296 531972 356302 532024
rect 316678 531904 316684 531956
rect 316736 531944 316742 531956
rect 319898 531944 319904 531956
rect 316736 531916 319904 531944
rect 316736 531904 316742 531916
rect 319898 531904 319904 531916
rect 319956 531904 319962 531956
rect 319990 531904 319996 531956
rect 320048 531944 320054 531956
rect 419534 531944 419540 531956
rect 320048 531916 419540 531944
rect 320048 531904 320054 531916
rect 419534 531904 419540 531916
rect 419592 531904 419598 531956
rect 318426 531836 318432 531888
rect 318484 531876 318490 531888
rect 423950 531876 423956 531888
rect 318484 531848 423956 531876
rect 318484 531836 318490 531848
rect 423950 531836 423956 531848
rect 424008 531836 424014 531888
rect 301958 531768 301964 531820
rect 302016 531808 302022 531820
rect 401594 531808 401600 531820
rect 302016 531780 401600 531808
rect 302016 531768 302022 531780
rect 401594 531768 401600 531780
rect 401652 531768 401658 531820
rect 318058 531700 318064 531752
rect 318116 531740 318122 531752
rect 319990 531740 319996 531752
rect 318116 531712 319996 531740
rect 318116 531700 318122 531712
rect 319990 531700 319996 531712
rect 320048 531700 320054 531752
rect 312630 531224 312636 531276
rect 312688 531264 312694 531276
rect 474734 531264 474740 531276
rect 312688 531236 474740 531264
rect 312688 531224 312694 531236
rect 474734 531224 474740 531236
rect 474792 531224 474798 531276
rect 315482 531156 315488 531208
rect 315540 531196 315546 531208
rect 428366 531196 428372 531208
rect 315540 531168 428372 531196
rect 315540 531156 315546 531168
rect 428366 531156 428372 531168
rect 428424 531156 428430 531208
rect 303246 530544 303252 530596
rect 303304 530584 303310 530596
rect 518158 530584 518164 530596
rect 303304 530556 518164 530584
rect 303304 530544 303310 530556
rect 518158 530544 518164 530556
rect 518216 530544 518222 530596
rect 312538 529864 312544 529916
rect 312596 529904 312602 529916
rect 511994 529904 512000 529916
rect 312596 529876 512000 529904
rect 312596 529864 312602 529876
rect 511994 529864 512000 529876
rect 512052 529864 512058 529916
rect 315298 529796 315304 529848
rect 315356 529836 315362 529848
rect 429378 529836 429384 529848
rect 315356 529808 429384 529836
rect 315356 529796 315362 529808
rect 429378 529796 429384 529808
rect 429436 529796 429442 529848
rect 315390 529728 315396 529780
rect 315448 529768 315454 529780
rect 428550 529768 428556 529780
rect 315448 529740 428556 529768
rect 315448 529728 315454 529740
rect 428550 529728 428556 529740
rect 428608 529728 428614 529780
rect 302326 529184 302332 529236
rect 302384 529224 302390 529236
rect 578878 529224 578884 529236
rect 302384 529196 578884 529224
rect 302384 529184 302390 529196
rect 578878 529184 578884 529196
rect 578936 529184 578942 529236
rect 42702 525036 42708 525088
rect 42760 525076 42766 525088
rect 57698 525076 57704 525088
rect 42760 525048 57704 525076
rect 42760 525036 42766 525048
rect 57698 525036 57704 525048
rect 57756 525036 57762 525088
rect 302878 502324 302884 502376
rect 302936 502364 302942 502376
rect 540238 502364 540244 502376
rect 302936 502336 540244 502364
rect 302936 502324 302942 502336
rect 540238 502324 540244 502336
rect 540296 502324 540302 502376
rect 82906 494912 82912 494964
rect 82964 494952 82970 494964
rect 83182 494952 83188 494964
rect 82964 494924 83188 494952
rect 82964 494912 82970 494924
rect 83182 494912 83188 494924
rect 83240 494912 83246 494964
rect 128354 494912 128360 494964
rect 128412 494952 128418 494964
rect 128538 494952 128544 494964
rect 128412 494924 128544 494952
rect 128412 494912 128418 494924
rect 128538 494912 128544 494924
rect 128596 494912 128602 494964
rect 136634 494912 136640 494964
rect 136692 494952 136698 494964
rect 136910 494952 136916 494964
rect 136692 494924 136916 494952
rect 136692 494912 136698 494924
rect 136910 494912 136916 494924
rect 136968 494912 136974 494964
rect 176746 494912 176752 494964
rect 176804 494952 176810 494964
rect 177022 494952 177028 494964
rect 176804 494924 177028 494952
rect 176804 494912 176810 494924
rect 177022 494912 177028 494924
rect 177080 494912 177086 494964
rect 229094 494912 229100 494964
rect 229152 494952 229158 494964
rect 229462 494952 229468 494964
rect 229152 494924 229468 494952
rect 229152 494912 229158 494924
rect 229462 494912 229468 494924
rect 229520 494912 229526 494964
rect 259546 494912 259552 494964
rect 259604 494952 259610 494964
rect 259822 494952 259828 494964
rect 259604 494924 259828 494952
rect 259604 494912 259610 494924
rect 259822 494912 259828 494924
rect 259880 494912 259886 494964
rect 197554 494776 197560 494828
rect 197612 494816 197618 494828
rect 198274 494816 198280 494828
rect 197612 494788 198280 494816
rect 197612 494776 197618 494788
rect 198274 494776 198280 494788
rect 198332 494776 198338 494828
rect 207214 494776 207220 494828
rect 207272 494816 207278 494828
rect 207382 494816 207388 494828
rect 207272 494788 207388 494816
rect 207272 494776 207278 494788
rect 207382 494776 207388 494788
rect 207440 494776 207446 494828
rect 242910 494776 242916 494828
rect 242968 494816 242974 494828
rect 243078 494816 243084 494828
rect 242968 494788 243084 494816
rect 242968 494776 242974 494788
rect 243078 494776 243084 494788
rect 243136 494776 243142 494828
rect 244366 494776 244372 494828
rect 244424 494816 244430 494828
rect 244550 494816 244556 494828
rect 244424 494788 244556 494816
rect 244424 494776 244430 494788
rect 244550 494776 244556 494788
rect 244608 494776 244614 494828
rect 273270 494776 273276 494828
rect 273328 494816 273334 494828
rect 273438 494816 273444 494828
rect 273328 494788 273444 494816
rect 273328 494776 273334 494788
rect 273438 494776 273444 494788
rect 273496 494776 273502 494828
rect 284310 494776 284316 494828
rect 284368 494816 284374 494828
rect 284478 494816 284484 494828
rect 284368 494788 284484 494816
rect 284368 494776 284374 494788
rect 284478 494776 284484 494788
rect 284536 494776 284542 494828
rect 498194 493960 498200 494012
rect 498252 494000 498258 494012
rect 580166 494000 580172 494012
rect 498252 493972 580172 494000
rect 498252 493960 498258 493972
rect 580166 493960 580172 493972
rect 580224 493960 580230 494012
rect 56318 493348 56324 493400
rect 56376 493388 56382 493400
rect 90542 493388 90548 493400
rect 56376 493360 90548 493388
rect 56376 493348 56382 493360
rect 90542 493348 90548 493360
rect 90600 493348 90606 493400
rect 51810 493280 51816 493332
rect 51868 493320 51874 493332
rect 99374 493320 99380 493332
rect 51868 493292 99380 493320
rect 51868 493280 51874 493292
rect 99374 493280 99380 493292
rect 99432 493280 99438 493332
rect 109770 493280 109776 493332
rect 109828 493320 109834 493332
rect 207106 493320 207112 493332
rect 109828 493292 207112 493320
rect 109828 493280 109834 493292
rect 207106 493280 207112 493292
rect 207164 493280 207170 493332
rect 161566 492736 161572 492788
rect 161624 492776 161630 492788
rect 161934 492776 161940 492788
rect 161624 492748 161940 492776
rect 161624 492736 161630 492748
rect 161934 492736 161940 492748
rect 161992 492736 161998 492788
rect 166994 492736 167000 492788
rect 167052 492776 167058 492788
rect 167730 492776 167736 492788
rect 167052 492748 167736 492776
rect 167052 492736 167058 492748
rect 167730 492736 167736 492748
rect 167788 492736 167794 492788
rect 219526 492736 219532 492788
rect 219584 492736 219590 492788
rect 220998 492736 221004 492788
rect 221056 492776 221062 492788
rect 221182 492776 221188 492788
rect 221056 492748 221188 492776
rect 221056 492736 221062 492748
rect 221182 492736 221188 492748
rect 221240 492736 221246 492788
rect 69106 492668 69112 492720
rect 69164 492708 69170 492720
rect 69934 492708 69940 492720
rect 69164 492680 69940 492708
rect 69164 492668 69170 492680
rect 69934 492668 69940 492680
rect 69992 492668 69998 492720
rect 74626 492668 74632 492720
rect 74684 492708 74690 492720
rect 75270 492708 75276 492720
rect 74684 492680 75276 492708
rect 74684 492668 74690 492680
rect 75270 492668 75276 492680
rect 75328 492668 75334 492720
rect 75914 492668 75920 492720
rect 75972 492708 75978 492720
rect 76558 492708 76564 492720
rect 75972 492680 76564 492708
rect 75972 492668 75978 492680
rect 76558 492668 76564 492680
rect 76616 492668 76622 492720
rect 78674 492668 78680 492720
rect 78732 492708 78738 492720
rect 79686 492708 79692 492720
rect 78732 492680 79692 492708
rect 78732 492668 78738 492680
rect 79686 492668 79692 492680
rect 79744 492668 79750 492720
rect 161474 492668 161480 492720
rect 161532 492708 161538 492720
rect 161750 492708 161756 492720
rect 161532 492680 161756 492708
rect 161532 492668 161538 492680
rect 161750 492668 161756 492680
rect 161808 492668 161814 492720
rect 162854 492668 162860 492720
rect 162912 492708 162918 492720
rect 163314 492708 163320 492720
rect 162912 492680 163320 492708
rect 162912 492668 162918 492680
rect 163314 492668 163320 492680
rect 163372 492668 163378 492720
rect 164234 492668 164240 492720
rect 164292 492708 164298 492720
rect 165062 492708 165068 492720
rect 164292 492680 165068 492708
rect 164292 492668 164298 492680
rect 165062 492668 165068 492680
rect 165120 492668 165126 492720
rect 167086 492668 167092 492720
rect 167144 492708 167150 492720
rect 167270 492708 167276 492720
rect 167144 492680 167276 492708
rect 167144 492668 167150 492680
rect 167270 492668 167276 492680
rect 167328 492668 167334 492720
rect 168466 492668 168472 492720
rect 168524 492708 168530 492720
rect 169110 492708 169116 492720
rect 168524 492680 169116 492708
rect 168524 492668 168530 492680
rect 169110 492668 169116 492680
rect 169168 492668 169174 492720
rect 169846 492668 169852 492720
rect 169904 492708 169910 492720
rect 170398 492708 170404 492720
rect 169904 492680 170404 492708
rect 169904 492668 169910 492680
rect 170398 492668 170404 492680
rect 170456 492668 170462 492720
rect 171226 492668 171232 492720
rect 171284 492708 171290 492720
rect 172054 492708 172060 492720
rect 171284 492680 172060 492708
rect 171284 492668 171290 492680
rect 172054 492668 172060 492680
rect 172112 492668 172118 492720
rect 172606 492668 172612 492720
rect 172664 492708 172670 492720
rect 173526 492708 173532 492720
rect 172664 492680 173532 492708
rect 172664 492668 172670 492680
rect 173526 492668 173532 492680
rect 173584 492668 173590 492720
rect 173986 492668 173992 492720
rect 174044 492708 174050 492720
rect 174814 492708 174820 492720
rect 174044 492680 174820 492708
rect 174044 492668 174050 492680
rect 174814 492668 174820 492680
rect 174872 492668 174878 492720
rect 175274 492668 175280 492720
rect 175332 492708 175338 492720
rect 176102 492708 176108 492720
rect 175332 492680 176108 492708
rect 175332 492668 175338 492680
rect 176102 492668 176108 492680
rect 176160 492668 176166 492720
rect 176654 492668 176660 492720
rect 176712 492708 176718 492720
rect 177390 492708 177396 492720
rect 176712 492680 177396 492708
rect 176712 492668 176718 492680
rect 177390 492668 177396 492680
rect 177448 492668 177454 492720
rect 178034 492668 178040 492720
rect 178092 492708 178098 492720
rect 178678 492708 178684 492720
rect 178092 492680 178684 492708
rect 178092 492668 178098 492680
rect 178678 492668 178684 492680
rect 178736 492668 178742 492720
rect 179414 492668 179420 492720
rect 179472 492708 179478 492720
rect 180058 492708 180064 492720
rect 179472 492680 180064 492708
rect 179472 492668 179478 492680
rect 180058 492668 180064 492680
rect 180116 492668 180122 492720
rect 180886 492668 180892 492720
rect 180944 492708 180950 492720
rect 181438 492708 181444 492720
rect 180944 492680 181444 492708
rect 180944 492668 180950 492680
rect 181438 492668 181444 492680
rect 181496 492668 181502 492720
rect 182174 492668 182180 492720
rect 182232 492708 182238 492720
rect 182726 492708 182732 492720
rect 182232 492680 182732 492708
rect 182232 492668 182238 492680
rect 182726 492668 182732 492680
rect 182784 492668 182790 492720
rect 184934 492668 184940 492720
rect 184992 492708 184998 492720
rect 185854 492708 185860 492720
rect 184992 492680 185860 492708
rect 184992 492668 184998 492680
rect 185854 492668 185860 492680
rect 185912 492668 185918 492720
rect 59262 492600 59268 492652
rect 59320 492640 59326 492652
rect 59320 492612 89714 492640
rect 59320 492600 59326 492612
rect 60090 492532 60096 492584
rect 60148 492572 60154 492584
rect 61930 492572 61936 492584
rect 60148 492544 61936 492572
rect 60148 492532 60154 492544
rect 61930 492532 61936 492544
rect 61988 492532 61994 492584
rect 62114 492532 62120 492584
rect 62172 492572 62178 492584
rect 62942 492572 62948 492584
rect 62172 492544 62948 492572
rect 62172 492532 62178 492544
rect 62942 492532 62948 492544
rect 63000 492532 63006 492584
rect 63034 492532 63040 492584
rect 63092 492572 63098 492584
rect 88794 492572 88800 492584
rect 63092 492544 88800 492572
rect 63092 492532 63098 492544
rect 88794 492532 88800 492544
rect 88852 492532 88858 492584
rect 89686 492572 89714 492612
rect 139394 492600 139400 492652
rect 139452 492640 139458 492652
rect 139854 492640 139860 492652
rect 139452 492612 139860 492640
rect 139452 492600 139458 492612
rect 139854 492600 139860 492612
rect 139912 492600 139918 492652
rect 150434 492600 150440 492652
rect 150492 492640 150498 492652
rect 150492 492612 151814 492640
rect 150492 492600 150498 492612
rect 91094 492572 91100 492584
rect 89686 492544 91100 492572
rect 91094 492532 91100 492544
rect 91152 492532 91158 492584
rect 92566 492532 92572 492584
rect 92624 492572 92630 492584
rect 93302 492572 93308 492584
rect 92624 492544 93308 492572
rect 92624 492532 92630 492544
rect 93302 492532 93308 492544
rect 93360 492532 93366 492584
rect 129918 492532 129924 492584
rect 129976 492572 129982 492584
rect 130102 492572 130108 492584
rect 129976 492544 130108 492572
rect 129976 492532 129982 492544
rect 130102 492532 130108 492544
rect 130160 492532 130166 492584
rect 50890 492464 50896 492516
rect 50948 492504 50954 492516
rect 84378 492504 84384 492516
rect 50948 492476 84384 492504
rect 50948 492464 50954 492476
rect 84378 492464 84384 492476
rect 84436 492464 84442 492516
rect 92474 492464 92480 492516
rect 92532 492504 92538 492516
rect 92934 492504 92940 492516
rect 92532 492476 92940 492504
rect 92532 492464 92538 492476
rect 92934 492464 92940 492476
rect 92992 492464 92998 492516
rect 102226 492464 102232 492516
rect 102284 492504 102290 492516
rect 103054 492504 103060 492516
rect 102284 492476 103060 492504
rect 102284 492464 102290 492476
rect 103054 492464 103060 492476
rect 103112 492464 103118 492516
rect 106366 492464 106372 492516
rect 106424 492504 106430 492516
rect 106918 492504 106924 492516
rect 106424 492476 106924 492504
rect 106424 492464 106430 492476
rect 106918 492464 106924 492476
rect 106976 492464 106982 492516
rect 107654 492464 107660 492516
rect 107712 492504 107718 492516
rect 107838 492504 107844 492516
rect 107712 492476 107844 492504
rect 107712 492464 107718 492476
rect 107838 492464 107844 492476
rect 107896 492464 107902 492516
rect 118694 492464 118700 492516
rect 118752 492504 118758 492516
rect 119246 492504 119252 492516
rect 118752 492476 119252 492504
rect 118752 492464 118758 492476
rect 119246 492464 119252 492476
rect 119304 492464 119310 492516
rect 120074 492464 120080 492516
rect 120132 492504 120138 492516
rect 120534 492504 120540 492516
rect 120132 492476 120540 492504
rect 120132 492464 120138 492476
rect 120534 492464 120540 492476
rect 120592 492464 120598 492516
rect 122926 492464 122932 492516
rect 122984 492504 122990 492516
rect 123294 492504 123300 492516
rect 122984 492476 123300 492504
rect 122984 492464 122990 492476
rect 123294 492464 123300 492476
rect 123352 492464 123358 492516
rect 124306 492464 124312 492516
rect 124364 492504 124370 492516
rect 124950 492504 124956 492516
rect 124364 492476 124956 492504
rect 124364 492464 124370 492476
rect 124950 492464 124956 492476
rect 125008 492464 125014 492516
rect 125686 492464 125692 492516
rect 125744 492504 125750 492516
rect 125870 492504 125876 492516
rect 125744 492476 125876 492504
rect 125744 492464 125750 492476
rect 125870 492464 125876 492476
rect 125928 492464 125934 492516
rect 126974 492464 126980 492516
rect 127032 492504 127038 492516
rect 127158 492504 127164 492516
rect 127032 492476 127164 492504
rect 127032 492464 127038 492476
rect 127158 492464 127164 492476
rect 127216 492464 127222 492516
rect 129734 492464 129740 492516
rect 129792 492504 129798 492516
rect 130654 492504 130660 492516
rect 129792 492476 130660 492504
rect 129792 492464 129798 492476
rect 130654 492464 130660 492476
rect 130712 492464 130718 492516
rect 131114 492464 131120 492516
rect 131172 492504 131178 492516
rect 131574 492504 131580 492516
rect 131172 492476 131580 492504
rect 131172 492464 131178 492476
rect 131574 492464 131580 492476
rect 131632 492464 131638 492516
rect 133966 492464 133972 492516
rect 134024 492504 134030 492516
rect 134702 492504 134708 492516
rect 134024 492476 134708 492504
rect 134024 492464 134030 492476
rect 134702 492464 134708 492476
rect 134760 492464 134766 492516
rect 135346 492464 135352 492516
rect 135404 492504 135410 492516
rect 135990 492504 135996 492516
rect 135404 492476 135996 492504
rect 135404 492464 135410 492476
rect 135990 492464 135996 492476
rect 136048 492464 136054 492516
rect 138014 492464 138020 492516
rect 138072 492504 138078 492516
rect 138658 492504 138664 492516
rect 138072 492476 138664 492504
rect 138072 492464 138078 492476
rect 138658 492464 138664 492476
rect 138716 492464 138722 492516
rect 139394 492464 139400 492516
rect 139452 492504 139458 492516
rect 140038 492504 140044 492516
rect 139452 492476 140044 492504
rect 139452 492464 139458 492476
rect 140038 492464 140044 492476
rect 140096 492464 140102 492516
rect 140958 492464 140964 492516
rect 141016 492504 141022 492516
rect 141694 492504 141700 492516
rect 141016 492476 141700 492504
rect 141016 492464 141022 492476
rect 141694 492464 141700 492476
rect 141752 492464 141758 492516
rect 143534 492464 143540 492516
rect 143592 492504 143598 492516
rect 143902 492504 143908 492516
rect 143592 492476 143908 492504
rect 143592 492464 143598 492476
rect 143902 492464 143908 492476
rect 143960 492464 143966 492516
rect 146294 492464 146300 492516
rect 146352 492504 146358 492516
rect 147030 492504 147036 492516
rect 146352 492476 147036 492504
rect 146352 492464 146358 492476
rect 147030 492464 147036 492476
rect 147088 492464 147094 492516
rect 150434 492464 150440 492516
rect 150492 492504 150498 492516
rect 151538 492504 151544 492516
rect 150492 492476 151544 492504
rect 150492 492464 150498 492476
rect 151538 492464 151544 492476
rect 151596 492464 151602 492516
rect 50522 492396 50528 492448
rect 50580 492436 50586 492448
rect 50580 492408 67588 492436
rect 50580 492396 50586 492408
rect 62022 492328 62028 492380
rect 62080 492368 62086 492380
rect 62758 492368 62764 492380
rect 62080 492340 62764 492368
rect 62080 492328 62086 492340
rect 62758 492328 62764 492340
rect 62816 492328 62822 492380
rect 64874 492328 64880 492380
rect 64932 492368 64938 492380
rect 65518 492368 65524 492380
rect 64932 492340 65524 492368
rect 64932 492328 64938 492340
rect 65518 492328 65524 492340
rect 65576 492328 65582 492380
rect 56410 492260 56416 492312
rect 56468 492300 56474 492312
rect 63034 492300 63040 492312
rect 56468 492272 63040 492300
rect 56468 492260 56474 492272
rect 63034 492260 63040 492272
rect 63092 492260 63098 492312
rect 67560 492300 67588 492408
rect 67726 492396 67732 492448
rect 67784 492436 67790 492448
rect 68186 492436 68192 492448
rect 67784 492408 68192 492436
rect 67784 492396 67790 492408
rect 68186 492396 68192 492408
rect 68244 492396 68250 492448
rect 68278 492396 68284 492448
rect 68336 492436 68342 492448
rect 68336 492408 69152 492436
rect 68336 492396 68342 492408
rect 67634 492328 67640 492380
rect 67692 492368 67698 492380
rect 67910 492368 67916 492380
rect 67692 492340 67916 492368
rect 67692 492328 67698 492340
rect 67910 492328 67916 492340
rect 67968 492328 67974 492380
rect 68370 492328 68376 492380
rect 68428 492368 68434 492380
rect 69124 492368 69152 492408
rect 71774 492396 71780 492448
rect 71832 492436 71838 492448
rect 72142 492436 72148 492448
rect 71832 492408 72148 492436
rect 71832 492396 71838 492408
rect 72142 492396 72148 492408
rect 72200 492396 72206 492448
rect 72510 492396 72516 492448
rect 72568 492436 72574 492448
rect 106274 492436 106280 492448
rect 72568 492408 106280 492436
rect 72568 492396 72574 492408
rect 106274 492396 106280 492408
rect 106332 492396 106338 492448
rect 122834 492396 122840 492448
rect 122892 492436 122898 492448
rect 123662 492436 123668 492448
rect 122892 492408 123668 492436
rect 122892 492396 122898 492408
rect 123662 492396 123668 492408
rect 123720 492396 123726 492448
rect 125594 492396 125600 492448
rect 125652 492436 125658 492448
rect 126330 492436 126336 492448
rect 125652 492408 126336 492436
rect 125652 492396 125658 492408
rect 126330 492396 126336 492408
rect 126388 492396 126394 492448
rect 131206 492396 131212 492448
rect 131264 492436 131270 492448
rect 132126 492436 132132 492448
rect 131264 492408 132132 492436
rect 131264 492396 131270 492408
rect 132126 492396 132132 492408
rect 132184 492396 132190 492448
rect 104618 492368 104624 492380
rect 68428 492340 69060 492368
rect 69124 492340 104624 492368
rect 68428 492328 68434 492340
rect 68922 492300 68928 492312
rect 67560 492272 68928 492300
rect 68922 492260 68928 492272
rect 68980 492260 68986 492312
rect 69032 492300 69060 492340
rect 104618 492328 104624 492340
rect 104676 492328 104682 492380
rect 151786 492368 151814 492612
rect 156690 492600 156696 492652
rect 156748 492640 156754 492652
rect 212810 492640 212816 492652
rect 156748 492612 212816 492640
rect 156748 492600 156754 492612
rect 212810 492600 212816 492612
rect 212868 492600 212874 492652
rect 219544 492584 219572 492736
rect 248598 492668 248604 492720
rect 248656 492708 248662 492720
rect 248656 492680 249196 492708
rect 248656 492668 248662 492680
rect 249168 492640 249196 492680
rect 255256 492680 256464 492708
rect 255256 492640 255284 492680
rect 249168 492612 255284 492640
rect 255314 492600 255320 492652
rect 255372 492640 255378 492652
rect 256326 492640 256332 492652
rect 255372 492612 256332 492640
rect 255372 492600 255378 492612
rect 256326 492600 256332 492612
rect 256384 492600 256390 492652
rect 155310 492532 155316 492584
rect 155368 492572 155374 492584
rect 211154 492572 211160 492584
rect 155368 492544 211160 492572
rect 155368 492532 155374 492544
rect 211154 492532 211160 492544
rect 211212 492532 211218 492584
rect 219526 492532 219532 492584
rect 219584 492532 219590 492584
rect 240042 492532 240048 492584
rect 240100 492572 240106 492584
rect 240100 492544 253934 492572
rect 240100 492532 240106 492544
rect 157334 492464 157340 492516
rect 157392 492504 157398 492516
rect 158070 492504 158076 492516
rect 157392 492476 158076 492504
rect 157392 492464 157398 492476
rect 158070 492464 158076 492476
rect 158128 492464 158134 492516
rect 160094 492464 160100 492516
rect 160152 492504 160158 492516
rect 160646 492504 160652 492516
rect 160152 492476 160652 492504
rect 160152 492464 160158 492476
rect 160646 492464 160652 492476
rect 160704 492464 160710 492516
rect 160756 492476 201556 492504
rect 153102 492396 153108 492448
rect 153160 492436 153166 492448
rect 160756 492436 160784 492476
rect 153160 492408 160784 492436
rect 153160 492396 153166 492408
rect 160830 492396 160836 492448
rect 160888 492436 160894 492448
rect 160888 492408 201356 492436
rect 160888 492396 160894 492408
rect 200850 492368 200856 492380
rect 151786 492340 200856 492368
rect 200850 492328 200856 492340
rect 200908 492328 200914 492380
rect 104894 492300 104900 492312
rect 69032 492272 104900 492300
rect 104894 492260 104900 492272
rect 104952 492260 104958 492312
rect 151446 492260 151452 492312
rect 151504 492300 151510 492312
rect 191098 492300 191104 492312
rect 151504 492272 191104 492300
rect 151504 492260 151510 492272
rect 191098 492260 191104 492272
rect 191156 492260 191162 492312
rect 201328 492300 201356 492408
rect 201528 492368 201556 492476
rect 201586 492464 201592 492516
rect 201644 492504 201650 492516
rect 202046 492504 202052 492516
rect 201644 492476 202052 492504
rect 201644 492464 201650 492476
rect 202046 492464 202052 492476
rect 202104 492464 202110 492516
rect 202966 492464 202972 492516
rect 203024 492504 203030 492516
rect 203886 492504 203892 492516
rect 203024 492476 203892 492504
rect 203024 492464 203030 492476
rect 203886 492464 203892 492476
rect 203944 492464 203950 492516
rect 208486 492464 208492 492516
rect 208544 492504 208550 492516
rect 208670 492504 208676 492516
rect 208544 492476 208676 492504
rect 208544 492464 208550 492476
rect 208670 492464 208676 492476
rect 208728 492464 208734 492516
rect 209866 492464 209872 492516
rect 209924 492504 209930 492516
rect 210510 492504 210516 492516
rect 209924 492476 210516 492504
rect 209924 492464 209930 492476
rect 210510 492464 210516 492476
rect 210568 492464 210574 492516
rect 212718 492464 212724 492516
rect 212776 492504 212782 492516
rect 213454 492504 213460 492516
rect 212776 492476 213460 492504
rect 212776 492464 212782 492476
rect 213454 492464 213460 492476
rect 213512 492464 213518 492516
rect 215294 492464 215300 492516
rect 215352 492504 215358 492516
rect 216214 492504 216220 492516
rect 215352 492476 216220 492504
rect 215352 492464 215358 492476
rect 216214 492464 216220 492476
rect 216272 492464 216278 492516
rect 218054 492464 218060 492516
rect 218112 492504 218118 492516
rect 218790 492504 218796 492516
rect 218112 492476 218796 492504
rect 218112 492464 218118 492476
rect 218790 492464 218796 492476
rect 218848 492464 218854 492516
rect 223574 492464 223580 492516
rect 223632 492504 223638 492516
rect 223758 492504 223764 492516
rect 223632 492476 223764 492504
rect 223632 492464 223638 492476
rect 223758 492464 223764 492476
rect 223816 492464 223822 492516
rect 253906 492504 253934 492544
rect 255406 492532 255412 492584
rect 255464 492572 255470 492584
rect 255774 492572 255780 492584
rect 255464 492544 255780 492572
rect 255464 492532 255470 492544
rect 255774 492532 255780 492544
rect 255832 492532 255838 492584
rect 256436 492572 256464 492680
rect 258166 492668 258172 492720
rect 258224 492708 258230 492720
rect 258902 492708 258908 492720
rect 258224 492680 258908 492708
rect 258224 492668 258230 492680
rect 258902 492668 258908 492680
rect 258960 492668 258966 492720
rect 262398 492668 262404 492720
rect 262456 492708 262462 492720
rect 262582 492708 262588 492720
rect 262456 492680 262588 492708
rect 262456 492668 262462 492680
rect 262582 492668 262588 492680
rect 262640 492668 262646 492720
rect 283006 492668 283012 492720
rect 283064 492708 283070 492720
rect 283558 492708 283564 492720
rect 283064 492680 283564 492708
rect 283064 492668 283070 492680
rect 283558 492668 283564 492680
rect 283616 492668 283622 492720
rect 291194 492668 291200 492720
rect 291252 492708 291258 492720
rect 291930 492708 291936 492720
rect 291252 492680 291936 492708
rect 291252 492668 291258 492680
rect 291930 492668 291936 492680
rect 291988 492668 291994 492720
rect 295334 492668 295340 492720
rect 295392 492708 295398 492720
rect 295886 492708 295892 492720
rect 295392 492680 295892 492708
rect 295392 492668 295398 492680
rect 295886 492668 295892 492680
rect 295944 492668 295950 492720
rect 256694 492600 256700 492652
rect 256752 492640 256758 492652
rect 257062 492640 257068 492652
rect 256752 492612 257068 492640
rect 256752 492600 256758 492612
rect 257062 492600 257068 492612
rect 257120 492600 257126 492652
rect 258074 492600 258080 492652
rect 258132 492640 258138 492652
rect 258534 492640 258540 492652
rect 258132 492612 258540 492640
rect 258132 492600 258138 492612
rect 258534 492600 258540 492612
rect 258592 492600 258598 492652
rect 259454 492600 259460 492652
rect 259512 492640 259518 492652
rect 260190 492640 260196 492652
rect 259512 492612 260196 492640
rect 259512 492600 259518 492612
rect 260190 492600 260196 492612
rect 260248 492600 260254 492652
rect 260834 492600 260840 492652
rect 260892 492640 260898 492652
rect 261478 492640 261484 492652
rect 260892 492612 261484 492640
rect 260892 492600 260898 492612
rect 261478 492600 261484 492612
rect 261536 492600 261542 492652
rect 262214 492600 262220 492652
rect 262272 492640 262278 492652
rect 262858 492640 262864 492652
rect 262272 492612 262864 492640
rect 262272 492600 262278 492612
rect 262858 492600 262864 492612
rect 262916 492600 262922 492652
rect 264974 492600 264980 492652
rect 265032 492640 265038 492652
rect 265894 492640 265900 492652
rect 265032 492612 265900 492640
rect 265032 492600 265038 492612
rect 265894 492600 265900 492612
rect 265952 492600 265958 492652
rect 267826 492600 267832 492652
rect 267884 492640 267890 492652
rect 268654 492640 268660 492652
rect 267884 492612 268660 492640
rect 267884 492600 267890 492612
rect 268654 492600 268660 492612
rect 268712 492600 268718 492652
rect 269114 492600 269120 492652
rect 269172 492640 269178 492652
rect 269942 492640 269948 492652
rect 269172 492612 269948 492640
rect 269172 492600 269178 492612
rect 269942 492600 269948 492612
rect 270000 492600 270006 492652
rect 270586 492600 270592 492652
rect 270644 492640 270650 492652
rect 271230 492640 271236 492652
rect 270644 492612 271236 492640
rect 270644 492600 270650 492612
rect 271230 492600 271236 492612
rect 271288 492600 271294 492652
rect 271966 492600 271972 492652
rect 272024 492640 272030 492652
rect 272518 492640 272524 492652
rect 272024 492612 272524 492640
rect 272024 492600 272030 492612
rect 272518 492600 272524 492612
rect 272576 492600 272582 492652
rect 282914 492600 282920 492652
rect 282972 492640 282978 492652
rect 283190 492640 283196 492652
rect 282972 492612 283196 492640
rect 282972 492600 282978 492612
rect 283190 492600 283196 492612
rect 283248 492600 283254 492652
rect 284294 492600 284300 492652
rect 284352 492640 284358 492652
rect 284846 492640 284852 492652
rect 284352 492612 284852 492640
rect 284352 492600 284358 492612
rect 284846 492600 284852 492612
rect 284904 492600 284910 492652
rect 285674 492600 285680 492652
rect 285732 492640 285738 492652
rect 286686 492640 286692 492652
rect 285732 492612 286692 492640
rect 285732 492600 285738 492612
rect 286686 492600 286692 492612
rect 286744 492600 286750 492652
rect 288434 492600 288440 492652
rect 288492 492640 288498 492652
rect 289262 492640 289268 492652
rect 288492 492612 289268 492640
rect 288492 492600 288498 492612
rect 289262 492600 289268 492612
rect 289320 492600 289326 492652
rect 291286 492600 291292 492652
rect 291344 492640 291350 492652
rect 291470 492640 291476 492652
rect 291344 492612 291476 492640
rect 291344 492600 291350 492612
rect 291470 492600 291476 492612
rect 291528 492600 291534 492652
rect 295518 492600 295524 492652
rect 295576 492640 295582 492652
rect 296254 492640 296260 492652
rect 295576 492612 296260 492640
rect 295576 492600 295582 492612
rect 296254 492600 296260 492612
rect 296312 492600 296318 492652
rect 296714 492600 296720 492652
rect 296772 492640 296778 492652
rect 297726 492640 297732 492652
rect 296772 492612 297732 492640
rect 296772 492600 296778 492612
rect 297726 492600 297732 492612
rect 297784 492600 297790 492652
rect 298186 492600 298192 492652
rect 298244 492640 298250 492652
rect 299014 492640 299020 492652
rect 298244 492612 299020 492640
rect 298244 492600 298250 492612
rect 299014 492600 299020 492612
rect 299072 492600 299078 492652
rect 356790 492572 356796 492584
rect 256436 492544 356796 492572
rect 356790 492532 356796 492544
rect 356848 492532 356854 492584
rect 358354 492504 358360 492516
rect 253906 492476 358360 492504
rect 358354 492464 358360 492476
rect 358412 492464 358418 492516
rect 208394 492396 208400 492448
rect 208452 492436 208458 492448
rect 209130 492436 209136 492448
rect 208452 492408 209136 492436
rect 208452 492396 208458 492408
rect 209130 492396 209136 492408
rect 209188 492396 209194 492448
rect 220906 492396 220912 492448
rect 220964 492436 220970 492448
rect 221458 492436 221464 492448
rect 220964 492408 221464 492436
rect 220964 492396 220970 492408
rect 221458 492396 221464 492408
rect 221516 492396 221522 492448
rect 239674 492396 239680 492448
rect 239732 492436 239738 492448
rect 358262 492436 358268 492448
rect 239732 492408 358268 492436
rect 239732 492396 239738 492408
rect 358262 492396 358268 492408
rect 358320 492396 358326 492448
rect 205726 492368 205732 492380
rect 201528 492340 205732 492368
rect 205726 492328 205732 492340
rect 205784 492328 205790 492380
rect 206370 492328 206376 492380
rect 206428 492368 206434 492380
rect 209222 492368 209228 492380
rect 206428 492340 209228 492368
rect 206428 492328 206434 492340
rect 209222 492328 209228 492340
rect 209280 492328 209286 492380
rect 219986 492328 219992 492380
rect 220044 492368 220050 492380
rect 222654 492368 222660 492380
rect 220044 492340 222660 492368
rect 220044 492328 220050 492340
rect 222654 492328 222660 492340
rect 222712 492328 222718 492380
rect 240778 492328 240784 492380
rect 240836 492368 240842 492380
rect 362310 492368 362316 492380
rect 240836 492340 362316 492368
rect 240836 492328 240842 492340
rect 362310 492328 362316 492340
rect 362368 492328 362374 492380
rect 201770 492300 201776 492312
rect 201328 492272 201776 492300
rect 201770 492260 201776 492272
rect 201828 492260 201834 492312
rect 240594 492260 240600 492312
rect 240652 492300 240658 492312
rect 366542 492300 366548 492312
rect 240652 492272 366548 492300
rect 240652 492260 240658 492272
rect 366542 492260 366548 492272
rect 366600 492260 366606 492312
rect 57238 492192 57244 492244
rect 57296 492232 57302 492244
rect 102410 492232 102416 492244
rect 57296 492204 102416 492232
rect 57296 492192 57302 492204
rect 102410 492192 102416 492204
rect 102468 492192 102474 492244
rect 121454 492192 121460 492244
rect 121512 492232 121518 492244
rect 121914 492232 121920 492244
rect 121512 492204 121920 492232
rect 121512 492192 121518 492204
rect 121914 492192 121920 492204
rect 121972 492192 121978 492244
rect 155218 492192 155224 492244
rect 155276 492232 155282 492244
rect 200666 492232 200672 492244
rect 155276 492204 200672 492232
rect 155276 492192 155282 492204
rect 200666 492192 200672 492204
rect 200724 492192 200730 492244
rect 226150 492232 226156 492244
rect 219406 492204 226156 492232
rect 53374 492124 53380 492176
rect 53432 492164 53438 492176
rect 100202 492164 100208 492176
rect 53432 492136 100208 492164
rect 53432 492124 53438 492136
rect 100202 492124 100208 492136
rect 100260 492124 100266 492176
rect 152274 492124 152280 492176
rect 152332 492164 152338 492176
rect 160830 492164 160836 492176
rect 152332 492136 160836 492164
rect 152332 492124 152338 492136
rect 160830 492124 160836 492136
rect 160888 492124 160894 492176
rect 160922 492124 160928 492176
rect 160980 492164 160986 492176
rect 190178 492164 190184 492176
rect 160980 492136 190184 492164
rect 160980 492124 160986 492136
rect 190178 492124 190184 492136
rect 190236 492124 190242 492176
rect 190288 492136 193214 492164
rect 49142 492056 49148 492108
rect 49200 492096 49206 492108
rect 97534 492096 97540 492108
rect 49200 492068 97540 492096
rect 49200 492056 49206 492068
rect 97534 492056 97540 492068
rect 97592 492056 97598 492108
rect 110138 492056 110144 492108
rect 110196 492096 110202 492108
rect 162118 492096 162124 492108
rect 110196 492068 162124 492096
rect 110196 492056 110202 492068
rect 162118 492056 162124 492068
rect 162176 492056 162182 492108
rect 164142 492056 164148 492108
rect 164200 492096 164206 492108
rect 190288 492096 190316 492136
rect 164200 492068 190316 492096
rect 193186 492096 193214 492136
rect 194962 492124 194968 492176
rect 195020 492164 195026 492176
rect 196986 492164 196992 492176
rect 195020 492136 196992 492164
rect 195020 492124 195026 492136
rect 196986 492124 196992 492136
rect 197044 492124 197050 492176
rect 218330 492124 218336 492176
rect 218388 492164 218394 492176
rect 219406 492164 219434 492204
rect 226150 492192 226156 492204
rect 226208 492192 226214 492244
rect 231394 492192 231400 492244
rect 231452 492232 231458 492244
rect 358170 492232 358176 492244
rect 231452 492204 358176 492232
rect 231452 492192 231458 492204
rect 358170 492192 358176 492204
rect 358228 492192 358234 492244
rect 218388 492136 219434 492164
rect 218388 492124 218394 492136
rect 226058 492124 226064 492176
rect 226116 492164 226122 492176
rect 356698 492164 356704 492176
rect 226116 492136 356704 492164
rect 226116 492124 226122 492136
rect 356698 492124 356704 492136
rect 356756 492124 356762 492176
rect 202138 492096 202144 492108
rect 193186 492068 202144 492096
rect 164200 492056 164206 492068
rect 202138 492056 202144 492068
rect 202196 492056 202202 492108
rect 202782 492056 202788 492108
rect 202840 492096 202846 492108
rect 212074 492096 212080 492108
rect 202840 492068 212080 492096
rect 202840 492056 202846 492068
rect 212074 492056 212080 492068
rect 212132 492056 212138 492108
rect 231762 492056 231768 492108
rect 231820 492096 231826 492108
rect 366358 492096 366364 492108
rect 231820 492068 366364 492096
rect 231820 492056 231826 492068
rect 366358 492056 366364 492068
rect 366416 492056 366422 492108
rect 62850 491988 62856 492040
rect 62908 492028 62914 492040
rect 129642 492028 129648 492040
rect 62908 492000 129648 492028
rect 62908 491988 62914 492000
rect 129642 491988 129648 492000
rect 129700 491988 129706 492040
rect 139854 491988 139860 492040
rect 139912 492028 139918 492040
rect 190086 492028 190092 492040
rect 139912 492000 190092 492028
rect 139912 491988 139918 492000
rect 190086 491988 190092 492000
rect 190144 491988 190150 492040
rect 190178 491988 190184 492040
rect 190236 492028 190242 492040
rect 197630 492028 197636 492040
rect 190236 492000 197636 492028
rect 190236 491988 190242 492000
rect 197630 491988 197636 492000
rect 197688 491988 197694 492040
rect 200298 491988 200304 492040
rect 200356 492028 200362 492040
rect 217410 492028 217416 492040
rect 200356 492000 217416 492028
rect 200356 491988 200362 492000
rect 217410 491988 217416 492000
rect 217468 491988 217474 492040
rect 225598 491988 225604 492040
rect 225656 492028 225662 492040
rect 362218 492028 362224 492040
rect 225656 492000 362224 492028
rect 225656 491988 225662 492000
rect 362218 491988 362224 492000
rect 362276 491988 362282 492040
rect 43898 491920 43904 491972
rect 43956 491960 43962 491972
rect 95326 491960 95332 491972
rect 43956 491932 95332 491960
rect 43956 491920 43962 491932
rect 95326 491920 95332 491932
rect 95384 491920 95390 491972
rect 110322 491920 110328 491972
rect 110380 491960 110386 491972
rect 192478 491960 192484 491972
rect 110380 491932 192484 491960
rect 110380 491920 110386 491932
rect 192478 491920 192484 491932
rect 192536 491920 192542 491972
rect 194502 491920 194508 491972
rect 194560 491960 194566 491972
rect 212442 491960 212448 491972
rect 194560 491932 212448 491960
rect 194560 491920 194566 491932
rect 212442 491920 212448 491932
rect 212500 491920 212506 491972
rect 223482 491920 223488 491972
rect 223540 491960 223546 491972
rect 363598 491960 363604 491972
rect 223540 491932 363604 491960
rect 223540 491920 223546 491932
rect 363598 491920 363604 491932
rect 363656 491920 363662 491972
rect 55030 491852 55036 491904
rect 55088 491892 55094 491904
rect 81710 491892 81716 491904
rect 55088 491864 81716 491892
rect 55088 491852 55094 491864
rect 81710 491852 81716 491864
rect 81768 491852 81774 491904
rect 157978 491852 157984 491904
rect 158036 491892 158042 491904
rect 197354 491892 197360 491904
rect 158036 491864 197360 491892
rect 158036 491852 158042 491864
rect 197354 491852 197360 491864
rect 197412 491852 197418 491904
rect 253934 491852 253940 491904
rect 253992 491892 253998 491904
rect 254210 491892 254216 491904
rect 253992 491864 254216 491892
rect 253992 491852 253998 491864
rect 254210 491852 254216 491864
rect 254268 491852 254274 491904
rect 256786 491852 256792 491904
rect 256844 491892 256850 491904
rect 257614 491892 257620 491904
rect 256844 491864 257620 491892
rect 256844 491852 256850 491864
rect 257614 491852 257620 491864
rect 257672 491852 257678 491904
rect 53742 491784 53748 491836
rect 53800 491824 53806 491836
rect 74534 491824 74540 491836
rect 53800 491796 74540 491824
rect 53800 491784 53806 491796
rect 74534 491784 74540 491796
rect 74592 491784 74598 491836
rect 153930 491784 153936 491836
rect 153988 491824 153994 491836
rect 160922 491824 160928 491836
rect 153988 491796 160928 491824
rect 153988 491784 153994 491796
rect 160922 491784 160928 491796
rect 160980 491784 160986 491836
rect 169754 491784 169760 491836
rect 169812 491824 169818 491836
rect 170030 491824 170036 491836
rect 169812 491796 170036 491824
rect 169812 491784 169818 491796
rect 170030 491784 170036 491796
rect 170088 491784 170094 491836
rect 198090 491824 198096 491836
rect 171106 491796 198096 491824
rect 52362 491716 52368 491768
rect 52420 491756 52426 491768
rect 71958 491756 71964 491768
rect 52420 491728 71964 491756
rect 52420 491716 52426 491728
rect 71958 491716 71964 491728
rect 72016 491716 72022 491768
rect 166902 491716 166908 491768
rect 166960 491756 166966 491768
rect 171106 491756 171134 491796
rect 198090 491784 198096 491796
rect 198148 491784 198154 491836
rect 292574 491784 292580 491836
rect 292632 491824 292638 491836
rect 292758 491824 292764 491836
rect 292632 491796 292764 491824
rect 292632 491784 292638 491796
rect 292758 491784 292764 491796
rect 292816 491784 292822 491836
rect 166960 491728 171134 491756
rect 166960 491716 166966 491728
rect 183462 491716 183468 491768
rect 183520 491756 183526 491768
rect 198182 491756 198188 491768
rect 183520 491728 198188 491756
rect 183520 491716 183526 491728
rect 198182 491716 198188 491728
rect 198240 491716 198246 491768
rect 253934 491716 253940 491768
rect 253992 491756 253998 491768
rect 254854 491756 254860 491768
rect 253992 491728 254860 491756
rect 253992 491716 253998 491728
rect 254854 491716 254860 491728
rect 254912 491716 254918 491768
rect 56502 491648 56508 491700
rect 56560 491688 56566 491700
rect 73798 491688 73804 491700
rect 56560 491660 73804 491688
rect 56560 491648 56566 491660
rect 73798 491648 73804 491660
rect 73856 491648 73862 491700
rect 191098 491648 191104 491700
rect 191156 491688 191162 491700
rect 197722 491688 197728 491700
rect 191156 491660 197728 491688
rect 191156 491648 191162 491660
rect 197722 491648 197728 491660
rect 197780 491648 197786 491700
rect 207198 491648 207204 491700
rect 207256 491688 207262 491700
rect 207750 491688 207756 491700
rect 207256 491660 207756 491688
rect 207256 491648 207262 491660
rect 207750 491648 207756 491660
rect 207808 491648 207814 491700
rect 190086 491580 190092 491632
rect 190144 491620 190150 491632
rect 193858 491620 193864 491632
rect 190144 491592 193864 491620
rect 190144 491580 190150 491592
rect 193858 491580 193864 491592
rect 193916 491580 193922 491632
rect 204162 491376 204168 491428
rect 204220 491416 204226 491428
rect 211614 491416 211620 491428
rect 204220 491388 211620 491416
rect 204220 491376 204226 491388
rect 211614 491376 211620 491388
rect 211672 491376 211678 491428
rect 199010 491308 199016 491360
rect 199068 491348 199074 491360
rect 202414 491348 202420 491360
rect 199068 491320 202420 491348
rect 199068 491308 199074 491320
rect 202414 491308 202420 491320
rect 202472 491308 202478 491360
rect 142154 491240 142160 491292
rect 142212 491280 142218 491292
rect 142614 491280 142620 491292
rect 142212 491252 142620 491280
rect 142212 491240 142218 491252
rect 142614 491240 142620 491252
rect 142672 491240 142678 491292
rect 267090 490764 267096 490816
rect 267148 490804 267154 490816
rect 359458 490804 359464 490816
rect 267148 490776 359464 490804
rect 267148 490764 267154 490776
rect 359458 490764 359464 490776
rect 359516 490764 359522 490816
rect 70394 490696 70400 490748
rect 70452 490736 70458 490748
rect 70854 490736 70860 490748
rect 70452 490708 70860 490736
rect 70452 490696 70458 490708
rect 70854 490696 70860 490708
rect 70912 490696 70918 490748
rect 260926 490696 260932 490748
rect 260984 490736 260990 490748
rect 368106 490736 368112 490748
rect 260984 490708 368112 490736
rect 260984 490696 260990 490708
rect 368106 490696 368112 490708
rect 368164 490696 368170 490748
rect 246482 490628 246488 490680
rect 246540 490668 246546 490680
rect 376110 490668 376116 490680
rect 246540 490640 376116 490668
rect 246540 490628 246546 490640
rect 376110 490628 376116 490640
rect 376168 490628 376174 490680
rect 58986 490560 58992 490612
rect 59044 490600 59050 490612
rect 96246 490600 96252 490612
rect 59044 490572 96252 490600
rect 59044 490560 59050 490572
rect 96246 490560 96252 490572
rect 96304 490560 96310 490612
rect 191834 490560 191840 490612
rect 191892 490600 191898 490612
rect 192386 490600 192392 490612
rect 191892 490572 192392 490600
rect 191892 490560 191898 490572
rect 192386 490560 192392 490572
rect 192444 490560 192450 490612
rect 222562 490560 222568 490612
rect 222620 490600 222626 490612
rect 376018 490600 376024 490612
rect 222620 490572 376024 490600
rect 222620 490560 222626 490572
rect 376018 490560 376024 490572
rect 376076 490560 376082 490612
rect 85758 490424 85764 490476
rect 85816 490464 85822 490476
rect 85942 490464 85948 490476
rect 85816 490436 85948 490464
rect 85816 490424 85822 490436
rect 85942 490424 85948 490436
rect 86000 490424 86006 490476
rect 87046 490424 87052 490476
rect 87104 490464 87110 490476
rect 87598 490464 87604 490476
rect 87104 490436 87604 490464
rect 87104 490424 87110 490436
rect 87598 490424 87604 490436
rect 87656 490424 87662 490476
rect 237466 490424 237472 490476
rect 237524 490464 237530 490476
rect 237742 490464 237748 490476
rect 237524 490436 237748 490464
rect 237524 490424 237530 490436
rect 237742 490424 237748 490436
rect 237800 490424 237806 490476
rect 274818 490424 274824 490476
rect 274876 490464 274882 490476
rect 275186 490464 275192 490476
rect 274876 490436 275192 490464
rect 274876 490424 274882 490436
rect 275186 490424 275192 490436
rect 275244 490424 275250 490476
rect 276014 490424 276020 490476
rect 276072 490464 276078 490476
rect 276934 490464 276940 490476
rect 276072 490436 276940 490464
rect 276072 490424 276078 490436
rect 276934 490424 276940 490436
rect 276992 490424 276998 490476
rect 80054 490356 80060 490408
rect 80112 490396 80118 490408
rect 80974 490396 80980 490408
rect 80112 490368 80980 490396
rect 80112 490356 80118 490368
rect 80974 490356 80980 490368
rect 81032 490356 81038 490408
rect 81526 490356 81532 490408
rect 81584 490396 81590 490408
rect 82262 490396 82268 490408
rect 81584 490368 82268 490396
rect 81584 490356 81590 490368
rect 82262 490356 82268 490368
rect 82320 490356 82326 490408
rect 82814 490356 82820 490408
rect 82872 490396 82878 490408
rect 83550 490396 83556 490408
rect 82872 490368 83556 490396
rect 82872 490356 82878 490368
rect 83550 490356 83556 490368
rect 83608 490356 83614 490408
rect 84286 490356 84292 490408
rect 84344 490396 84350 490408
rect 84930 490396 84936 490408
rect 84344 490368 84936 490396
rect 84344 490356 84350 490368
rect 84930 490356 84936 490368
rect 84988 490356 84994 490408
rect 85574 490356 85580 490408
rect 85632 490396 85638 490408
rect 86310 490396 86316 490408
rect 85632 490368 86316 490396
rect 85632 490356 85638 490368
rect 86310 490356 86316 490368
rect 86368 490356 86374 490408
rect 86954 490356 86960 490408
rect 87012 490396 87018 490408
rect 87230 490396 87236 490408
rect 87012 490368 87236 490396
rect 87012 490356 87018 490368
rect 87230 490356 87236 490368
rect 87288 490356 87294 490408
rect 111886 490356 111892 490408
rect 111944 490396 111950 490408
rect 112622 490396 112628 490408
rect 111944 490368 112628 490396
rect 111944 490356 111950 490368
rect 112622 490356 112628 490368
rect 112680 490356 112686 490408
rect 186314 490356 186320 490408
rect 186372 490396 186378 490408
rect 187142 490396 187148 490408
rect 186372 490368 187148 490396
rect 186372 490356 186378 490368
rect 187142 490356 187148 490368
rect 187200 490356 187206 490408
rect 192110 490356 192116 490408
rect 192168 490396 192174 490408
rect 192846 490396 192852 490408
rect 192168 490368 192852 490396
rect 192168 490356 192174 490368
rect 192846 490356 192852 490368
rect 192904 490356 192910 490408
rect 193214 490356 193220 490408
rect 193272 490396 193278 490408
rect 193766 490396 193772 490408
rect 193272 490368 193772 490396
rect 193272 490356 193278 490368
rect 193766 490356 193772 490368
rect 193824 490356 193830 490408
rect 194594 490356 194600 490408
rect 194652 490396 194658 490408
rect 195422 490396 195428 490408
rect 194652 490368 195428 490396
rect 194652 490356 194658 490368
rect 195422 490356 195428 490368
rect 195480 490356 195486 490408
rect 231854 490356 231860 490408
rect 231912 490396 231918 490408
rect 232406 490396 232412 490408
rect 231912 490368 232412 490396
rect 231912 490356 231918 490368
rect 232406 490356 232412 490368
rect 232464 490356 232470 490408
rect 233234 490356 233240 490408
rect 233292 490396 233298 490408
rect 234246 490396 234252 490408
rect 233292 490368 234252 490396
rect 233292 490356 233298 490368
rect 234246 490356 234252 490368
rect 234304 490356 234310 490408
rect 237374 490356 237380 490408
rect 237432 490396 237438 490408
rect 238202 490396 238208 490408
rect 237432 490368 238208 490396
rect 237432 490356 237438 490368
rect 238202 490356 238208 490368
rect 238260 490356 238266 490408
rect 242894 490356 242900 490408
rect 242952 490396 242958 490408
rect 243446 490396 243452 490408
rect 242952 490368 243452 490396
rect 242952 490356 242958 490368
rect 243446 490356 243452 490368
rect 243504 490356 243510 490408
rect 244366 490356 244372 490408
rect 244424 490396 244430 490408
rect 245286 490396 245292 490408
rect 244424 490368 245292 490396
rect 244424 490356 244430 490368
rect 245286 490356 245292 490368
rect 245344 490356 245350 490408
rect 245654 490356 245660 490408
rect 245712 490396 245718 490408
rect 246574 490396 246580 490408
rect 245712 490368 246580 490396
rect 245712 490356 245718 490368
rect 246574 490356 246580 490368
rect 246632 490356 246638 490408
rect 249794 490356 249800 490408
rect 249852 490396 249858 490408
rect 250530 490396 250536 490408
rect 249852 490368 250536 490396
rect 249852 490356 249858 490368
rect 250530 490356 250536 490368
rect 250588 490356 250594 490408
rect 273254 490356 273260 490408
rect 273312 490396 273318 490408
rect 273806 490396 273812 490408
rect 273312 490368 273812 490396
rect 273312 490356 273318 490368
rect 273806 490356 273812 490368
rect 273864 490356 273870 490408
rect 274634 490356 274640 490408
rect 274692 490396 274698 490408
rect 275646 490396 275652 490408
rect 274692 490368 275652 490396
rect 274692 490356 274698 490368
rect 275646 490356 275652 490368
rect 275704 490356 275710 490408
rect 276106 490356 276112 490408
rect 276164 490396 276170 490408
rect 276566 490396 276572 490408
rect 276164 490368 276572 490396
rect 276164 490356 276170 490368
rect 276566 490356 276572 490368
rect 276624 490356 276630 490408
rect 277486 490356 277492 490408
rect 277544 490396 277550 490408
rect 278222 490396 278228 490408
rect 277544 490368 278228 490396
rect 277544 490356 277550 490368
rect 278222 490356 278228 490368
rect 278280 490356 278286 490408
rect 280154 490356 280160 490408
rect 280212 490396 280218 490408
rect 280982 490396 280988 490408
rect 280212 490368 280988 490396
rect 280212 490356 280218 490368
rect 280982 490356 280988 490368
rect 281040 490356 281046 490408
rect 60734 490288 60740 490340
rect 60792 490328 60798 490340
rect 61102 490328 61108 490340
rect 60792 490300 61108 490328
rect 60792 490288 60798 490300
rect 61102 490288 61108 490300
rect 61160 490288 61166 490340
rect 187694 490152 187700 490204
rect 187752 490192 187758 490204
rect 188430 490192 188436 490204
rect 187752 490164 188436 490192
rect 187752 490152 187758 490164
rect 188430 490152 188436 490164
rect 188488 490152 188494 490204
rect 244642 490192 244648 490204
rect 244568 490164 244648 490192
rect 244568 490000 244596 490164
rect 244642 490152 244648 490164
rect 244700 490152 244706 490204
rect 244550 489948 244556 490000
rect 244608 489948 244614 490000
rect 50338 489812 50344 489864
rect 50396 489852 50402 489864
rect 98086 489852 98092 489864
rect 50396 489824 98092 489852
rect 50396 489812 50402 489824
rect 98086 489812 98092 489824
rect 98144 489812 98150 489864
rect 59814 489744 59820 489796
rect 59872 489784 59878 489796
rect 118694 489784 118700 489796
rect 59872 489756 118700 489784
rect 59872 489744 59878 489756
rect 118694 489744 118700 489756
rect 118752 489744 118758 489796
rect 48222 489676 48228 489728
rect 48280 489716 48286 489728
rect 111242 489716 111248 489728
rect 48280 489688 111248 489716
rect 48280 489676 48286 489688
rect 111242 489676 111248 489688
rect 111300 489676 111306 489728
rect 48038 489608 48044 489660
rect 48096 489648 48102 489660
rect 112070 489648 112076 489660
rect 48096 489620 112076 489648
rect 48096 489608 48102 489620
rect 112070 489608 112076 489620
rect 112128 489608 112134 489660
rect 46566 489540 46572 489592
rect 46624 489580 46630 489592
rect 111702 489580 111708 489592
rect 46624 489552 111708 489580
rect 46624 489540 46630 489552
rect 111702 489540 111708 489552
rect 111760 489540 111766 489592
rect 46290 489472 46296 489524
rect 46348 489512 46354 489524
rect 110782 489512 110788 489524
rect 46348 489484 110788 489512
rect 46348 489472 46354 489484
rect 110782 489472 110788 489484
rect 110840 489472 110846 489524
rect 138198 489472 138204 489524
rect 138256 489512 138262 489524
rect 200298 489512 200304 489524
rect 138256 489484 200304 489512
rect 138256 489472 138262 489484
rect 200298 489472 200304 489484
rect 200356 489472 200362 489524
rect 51718 489404 51724 489456
rect 51776 489444 51782 489456
rect 116026 489444 116032 489456
rect 51776 489416 116032 489444
rect 51776 489404 51782 489416
rect 116026 489404 116032 489416
rect 116084 489404 116090 489456
rect 136726 489404 136732 489456
rect 136784 489444 136790 489456
rect 198918 489444 198924 489456
rect 136784 489416 198924 489444
rect 136784 489404 136790 489416
rect 198918 489404 198924 489416
rect 198976 489404 198982 489456
rect 48958 489336 48964 489388
rect 49016 489376 49022 489388
rect 115198 489376 115204 489388
rect 49016 489348 115204 489376
rect 49016 489336 49022 489348
rect 115198 489336 115204 489348
rect 115256 489336 115262 489388
rect 138106 489336 138112 489388
rect 138164 489376 138170 489388
rect 200390 489376 200396 489388
rect 138164 489348 200396 489376
rect 138164 489336 138170 489348
rect 200390 489336 200396 489348
rect 200448 489336 200454 489388
rect 281810 489336 281816 489388
rect 281868 489376 281874 489388
rect 359550 489376 359556 489388
rect 281868 489348 359556 489376
rect 281868 489336 281874 489348
rect 359550 489336 359556 489348
rect 359608 489336 359614 489388
rect 57146 489268 57152 489320
rect 57204 489308 57210 489320
rect 132494 489308 132500 489320
rect 57204 489280 132500 489308
rect 57204 489268 57210 489280
rect 132494 489268 132500 489280
rect 132552 489268 132558 489320
rect 135438 489268 135444 489320
rect 135496 489308 135502 489320
rect 203242 489308 203248 489320
rect 135496 489280 203248 489308
rect 135496 489268 135502 489280
rect 203242 489268 203248 489280
rect 203300 489268 203306 489320
rect 247310 489268 247316 489320
rect 247368 489308 247374 489320
rect 370590 489308 370596 489320
rect 247368 489280 370596 489308
rect 247368 489268 247374 489280
rect 370590 489268 370596 489280
rect 370648 489268 370654 489320
rect 48682 489200 48688 489252
rect 48740 489240 48746 489252
rect 129734 489240 129740 489252
rect 48740 489212 129740 489240
rect 48740 489200 48746 489212
rect 129734 489200 129740 489212
rect 129792 489200 129798 489252
rect 136818 489200 136824 489252
rect 136876 489240 136882 489252
rect 205818 489240 205824 489252
rect 136876 489212 205824 489240
rect 136876 489200 136882 489212
rect 205818 489200 205824 489212
rect 205876 489200 205882 489252
rect 236730 489200 236736 489252
rect 236788 489240 236794 489252
rect 366450 489240 366456 489252
rect 236788 489212 366456 489240
rect 236788 489200 236794 489212
rect 366450 489200 366456 489212
rect 366508 489200 366514 489252
rect 61930 489132 61936 489184
rect 61988 489172 61994 489184
rect 180058 489172 180064 489184
rect 61988 489144 180064 489172
rect 61988 489132 61994 489144
rect 180058 489132 180064 489144
rect 180116 489132 180122 489184
rect 204346 489132 204352 489184
rect 204404 489172 204410 489184
rect 217318 489172 217324 489184
rect 204404 489144 217324 489172
rect 204404 489132 204410 489144
rect 217318 489132 217324 489144
rect 217376 489132 217382 489184
rect 239306 489132 239312 489184
rect 239364 489172 239370 489184
rect 376202 489172 376208 489184
rect 239364 489144 376208 489172
rect 239364 489132 239370 489144
rect 376202 489132 376208 489144
rect 376260 489132 376266 489184
rect 50430 489064 50436 489116
rect 50488 489104 50494 489116
rect 97994 489104 98000 489116
rect 50488 489076 98000 489104
rect 50488 489064 50494 489076
rect 97994 489064 98000 489076
rect 98052 489064 98058 489116
rect 54662 488996 54668 489048
rect 54720 489036 54726 489048
rect 96706 489036 96712 489048
rect 54720 489008 96712 489036
rect 54720 488996 54726 489008
rect 96706 488996 96712 489008
rect 96764 488996 96770 489048
rect 55766 488928 55772 488980
rect 55824 488968 55830 488980
rect 96798 488968 96804 488980
rect 55824 488940 96804 488968
rect 55824 488928 55830 488940
rect 96798 488928 96804 488940
rect 96856 488928 96862 488980
rect 283098 487840 283104 487892
rect 283156 487880 283162 487892
rect 359826 487880 359832 487892
rect 283156 487852 359832 487880
rect 283156 487840 283162 487852
rect 359826 487840 359832 487852
rect 359884 487840 359890 487892
rect 57698 487772 57704 487824
rect 57756 487812 57762 487824
rect 114278 487812 114284 487824
rect 57756 487784 114284 487812
rect 57756 487772 57762 487784
rect 114278 487772 114284 487784
rect 114336 487772 114342 487824
rect 158898 487772 158904 487824
rect 158956 487812 158962 487824
rect 218790 487812 218796 487824
rect 158956 487784 218796 487812
rect 158956 487772 158962 487784
rect 218790 487772 218796 487784
rect 218848 487772 218854 487824
rect 227622 487772 227628 487824
rect 227680 487812 227686 487824
rect 227806 487812 227812 487824
rect 227680 487784 227812 487812
rect 227680 487772 227686 487784
rect 227806 487772 227812 487784
rect 227864 487772 227870 487824
rect 244458 487772 244464 487824
rect 244516 487812 244522 487824
rect 244734 487812 244740 487824
rect 244516 487784 244740 487812
rect 244516 487772 244522 487784
rect 244734 487772 244740 487784
rect 244792 487772 244798 487824
rect 260926 487772 260932 487824
rect 260984 487812 260990 487824
rect 366726 487812 366732 487824
rect 260984 487784 366732 487812
rect 260984 487772 260990 487784
rect 366726 487772 366732 487784
rect 366784 487772 366790 487824
rect 226426 487296 226432 487348
rect 226484 487336 226490 487348
rect 226702 487336 226708 487348
rect 226484 487308 226708 487336
rect 226484 487296 226490 487308
rect 226702 487296 226708 487308
rect 226760 487296 226766 487348
rect 53190 487092 53196 487144
rect 53248 487132 53254 487144
rect 116946 487132 116952 487144
rect 53248 487104 116952 487132
rect 53248 487092 53254 487104
rect 116946 487092 116952 487104
rect 117004 487092 117010 487144
rect 53282 487024 53288 487076
rect 53340 487064 53346 487076
rect 116486 487064 116492 487076
rect 53340 487036 116492 487064
rect 53340 487024 53346 487036
rect 116486 487024 116492 487036
rect 116544 487024 116550 487076
rect 58618 486956 58624 487008
rect 58676 486996 58682 487008
rect 121546 486996 121552 487008
rect 58676 486968 121552 486996
rect 58676 486956 58682 486968
rect 121546 486956 121552 486968
rect 121604 486956 121610 487008
rect 59722 486888 59728 486940
rect 59780 486928 59786 486940
rect 130010 486928 130016 486940
rect 59780 486900 130016 486928
rect 59780 486888 59786 486900
rect 130010 486888 130016 486900
rect 130068 486888 130074 486940
rect 46658 486820 46664 486872
rect 46716 486860 46722 486872
rect 117406 486860 117412 486872
rect 46716 486832 117412 486860
rect 46716 486820 46722 486832
rect 117406 486820 117412 486832
rect 117464 486820 117470 486872
rect 229186 486820 229192 486872
rect 229244 486860 229250 486872
rect 229830 486860 229836 486872
rect 229244 486832 229836 486860
rect 229244 486820 229250 486832
rect 229830 486820 229836 486832
rect 229888 486820 229894 486872
rect 46382 486752 46388 486804
rect 46440 486792 46446 486804
rect 117866 486792 117872 486804
rect 46440 486764 117872 486792
rect 46440 486752 46446 486764
rect 117866 486752 117872 486764
rect 117924 486752 117930 486804
rect 189074 486752 189080 486804
rect 189132 486792 189138 486804
rect 189718 486792 189724 486804
rect 189132 486764 189724 486792
rect 189132 486752 189138 486764
rect 189718 486752 189724 486764
rect 189776 486752 189782 486804
rect 226334 486752 226340 486804
rect 226392 486792 226398 486804
rect 227254 486792 227260 486804
rect 226392 486764 227260 486792
rect 226392 486752 226398 486764
rect 227254 486752 227260 486764
rect 227312 486752 227318 486804
rect 46474 486684 46480 486736
rect 46532 486724 46538 486736
rect 118234 486724 118240 486736
rect 46532 486696 118240 486724
rect 46532 486684 46538 486696
rect 118234 486684 118240 486696
rect 118292 486684 118298 486736
rect 54386 486616 54392 486668
rect 54444 486656 54450 486668
rect 129918 486656 129924 486668
rect 54444 486628 129924 486656
rect 54444 486616 54450 486628
rect 129918 486616 129924 486628
rect 129976 486616 129982 486668
rect 50798 486548 50804 486600
rect 50856 486588 50862 486600
rect 131298 486588 131304 486600
rect 50856 486560 131304 486588
rect 50856 486548 50862 486560
rect 131298 486548 131304 486560
rect 131356 486548 131362 486600
rect 47946 486480 47952 486532
rect 48004 486520 48010 486532
rect 128538 486520 128544 486532
rect 48004 486492 128544 486520
rect 48004 486480 48010 486492
rect 128538 486480 128544 486492
rect 128596 486480 128602 486532
rect 242066 486480 242072 486532
rect 242124 486520 242130 486532
rect 370682 486520 370688 486532
rect 242124 486492 370688 486520
rect 242124 486480 242130 486492
rect 370682 486480 370688 486492
rect 370740 486480 370746 486532
rect 47854 486412 47860 486464
rect 47912 486452 47918 486464
rect 129826 486452 129832 486464
rect 47912 486424 129832 486452
rect 47912 486412 47918 486424
rect 129826 486412 129832 486424
rect 129884 486412 129890 486464
rect 223666 486412 223672 486464
rect 223724 486452 223730 486464
rect 363690 486452 363696 486464
rect 223724 486424 363696 486452
rect 223724 486412 223730 486424
rect 363690 486412 363696 486424
rect 363748 486412 363754 486464
rect 58894 486344 58900 486396
rect 58952 486384 58958 486396
rect 118786 486384 118792 486396
rect 58952 486356 118792 486384
rect 58952 486344 58958 486356
rect 118786 486344 118792 486356
rect 118844 486344 118850 486396
rect 58802 486276 58808 486328
rect 58860 486316 58866 486328
rect 118878 486316 118884 486328
rect 58860 486288 118884 486316
rect 58860 486276 58866 486288
rect 118878 486276 118884 486288
rect 118936 486276 118942 486328
rect 57882 486208 57888 486260
rect 57940 486248 57946 486260
rect 113910 486248 113916 486260
rect 57940 486220 113916 486248
rect 57940 486208 57946 486220
rect 113910 486208 113916 486220
rect 113968 486208 113974 486260
rect 256878 485188 256884 485240
rect 256936 485228 256942 485240
rect 369302 485228 369308 485240
rect 256936 485200 369308 485228
rect 256936 485188 256942 485200
rect 369302 485188 369308 485200
rect 369360 485188 369366 485240
rect 243078 485120 243084 485172
rect 243136 485160 243142 485172
rect 371970 485160 371976 485172
rect 243136 485132 371976 485160
rect 243136 485120 243142 485132
rect 371970 485120 371976 485132
rect 372028 485120 372034 485172
rect 165706 485052 165712 485104
rect 165764 485092 165770 485104
rect 209038 485092 209044 485104
rect 165764 485064 209044 485092
rect 165764 485052 165770 485064
rect 209038 485052 209044 485064
rect 209096 485052 209102 485104
rect 229278 485052 229284 485104
rect 229336 485092 229342 485104
rect 364978 485092 364984 485104
rect 229336 485064 364984 485092
rect 229336 485052 229342 485064
rect 364978 485052 364984 485064
rect 365036 485052 365042 485104
rect 57054 484304 57060 484356
rect 57112 484344 57118 484356
rect 128446 484344 128452 484356
rect 57112 484316 128452 484344
rect 57112 484304 57118 484316
rect 128446 484304 128452 484316
rect 128504 484304 128510 484356
rect 58710 484236 58716 484288
rect 58768 484276 58774 484288
rect 134058 484276 134064 484288
rect 58768 484248 134064 484276
rect 58768 484236 58774 484248
rect 134058 484236 134064 484248
rect 134116 484236 134122 484288
rect 48774 484168 48780 484220
rect 48832 484208 48838 484220
rect 124214 484208 124220 484220
rect 48832 484180 124220 484208
rect 48832 484168 48838 484180
rect 124214 484168 124220 484180
rect 124272 484168 124278 484220
rect 59630 484100 59636 484152
rect 59688 484140 59694 484152
rect 135346 484140 135352 484152
rect 59688 484112 135352 484140
rect 59688 484100 59694 484112
rect 135346 484100 135352 484112
rect 135404 484100 135410 484152
rect 45462 484032 45468 484084
rect 45520 484072 45526 484084
rect 124306 484072 124312 484084
rect 45520 484044 124312 484072
rect 45520 484032 45526 484044
rect 124306 484032 124312 484044
rect 124364 484032 124370 484084
rect 43622 483964 43628 484016
rect 43680 484004 43686 484016
rect 122926 484004 122932 484016
rect 43680 483976 122932 484004
rect 43680 483964 43686 483976
rect 122926 483964 122932 483976
rect 122984 483964 122990 484016
rect 42242 483896 42248 483948
rect 42300 483936 42306 483948
rect 124398 483936 124404 483948
rect 42300 483908 124404 483936
rect 42300 483896 42306 483908
rect 124398 483896 124404 483908
rect 124456 483896 124462 483948
rect 48866 483828 48872 483880
rect 48924 483868 48930 483880
rect 132678 483868 132684 483880
rect 48924 483840 132684 483868
rect 48924 483828 48930 483840
rect 132678 483828 132684 483840
rect 132736 483828 132742 483880
rect 46106 483760 46112 483812
rect 46164 483800 46170 483812
rect 132586 483800 132592 483812
rect 46164 483772 132592 483800
rect 46164 483760 46170 483772
rect 132586 483760 132592 483772
rect 132644 483760 132650 483812
rect 43346 483692 43352 483744
rect 43404 483732 43410 483744
rect 131206 483732 131212 483744
rect 43404 483704 131212 483732
rect 43404 483692 43410 483704
rect 131206 483692 131212 483704
rect 131264 483692 131270 483744
rect 292758 483692 292764 483744
rect 292816 483732 292822 483744
rect 379974 483732 379980 483744
rect 292816 483704 379980 483732
rect 292816 483692 292822 483704
rect 379974 483692 379980 483704
rect 380032 483692 380038 483744
rect 46014 483624 46020 483676
rect 46072 483664 46078 483676
rect 143626 483664 143632 483676
rect 46072 483636 143632 483664
rect 46072 483624 46078 483636
rect 143626 483624 143632 483636
rect 143684 483624 143690 483676
rect 167178 483624 167184 483676
rect 167236 483664 167242 483676
rect 215938 483664 215944 483676
rect 167236 483636 215944 483664
rect 167236 483624 167242 483636
rect 215938 483624 215944 483636
rect 215996 483624 216002 483676
rect 237558 483624 237564 483676
rect 237616 483664 237622 483676
rect 378870 483664 378876 483676
rect 237616 483636 378876 483664
rect 237616 483624 237622 483636
rect 378870 483624 378876 483636
rect 378928 483624 378934 483676
rect 58526 483556 58532 483608
rect 58584 483596 58590 483608
rect 128354 483596 128360 483608
rect 58584 483568 128360 483596
rect 58584 483556 58590 483568
rect 128354 483556 128360 483568
rect 128412 483556 128418 483608
rect 59354 483488 59360 483540
rect 59412 483528 59418 483540
rect 86218 483528 86224 483540
rect 59412 483500 86224 483528
rect 59412 483488 59418 483500
rect 86218 483488 86224 483500
rect 86276 483488 86282 483540
rect 262398 482400 262404 482452
rect 262456 482440 262462 482452
rect 373442 482440 373448 482452
rect 262456 482412 373448 482440
rect 262456 482400 262462 482412
rect 373442 482400 373448 482412
rect 373500 482400 373506 482452
rect 205634 482332 205640 482384
rect 205692 482372 205698 482384
rect 217594 482372 217600 482384
rect 205692 482344 217600 482372
rect 205692 482332 205698 482344
rect 217594 482332 217600 482344
rect 217652 482332 217658 482384
rect 235994 482332 236000 482384
rect 236052 482372 236058 482384
rect 367830 482372 367836 482384
rect 236052 482344 367836 482372
rect 236052 482332 236058 482344
rect 367830 482332 367836 482344
rect 367888 482332 367894 482384
rect 57606 482264 57612 482316
rect 57664 482304 57670 482316
rect 114554 482304 114560 482316
rect 57664 482276 114560 482304
rect 57664 482264 57670 482276
rect 114554 482264 114560 482276
rect 114612 482264 114618 482316
rect 168558 482264 168564 482316
rect 168616 482304 168622 482316
rect 210418 482304 210424 482316
rect 168616 482276 210424 482304
rect 168616 482264 168622 482276
rect 210418 482264 210424 482276
rect 210476 482264 210482 482316
rect 229094 482264 229100 482316
rect 229152 482304 229158 482316
rect 360930 482304 360936 482316
rect 229152 482276 360936 482304
rect 229152 482264 229158 482276
rect 360930 482264 360936 482276
rect 360988 482264 360994 482316
rect 295610 481108 295616 481160
rect 295668 481148 295674 481160
rect 376754 481148 376760 481160
rect 295668 481120 376760 481148
rect 295668 481108 295674 481120
rect 376754 481108 376760 481120
rect 376812 481108 376818 481160
rect 242986 481040 242992 481092
rect 243044 481080 243050 481092
rect 363782 481080 363788 481092
rect 243044 481052 363788 481080
rect 243044 481040 243050 481052
rect 363782 481040 363788 481052
rect 363840 481040 363846 481092
rect 149054 480972 149060 481024
rect 149112 481012 149118 481024
rect 211798 481012 211804 481024
rect 149112 480984 211804 481012
rect 149112 480972 149118 480984
rect 211798 480972 211804 480984
rect 211856 480972 211862 481024
rect 254210 480972 254216 481024
rect 254268 481012 254274 481024
rect 379054 481012 379060 481024
rect 254268 480984 379060 481012
rect 254268 480972 254274 480984
rect 379054 480972 379060 480984
rect 379112 480972 379118 481024
rect 60826 480904 60832 480956
rect 60884 480944 60890 480956
rect 199194 480944 199200 480956
rect 60884 480916 199200 480944
rect 60884 480904 60890 480916
rect 199194 480904 199200 480916
rect 199252 480904 199258 480956
rect 230474 480904 230480 480956
rect 230532 480944 230538 480956
rect 365070 480944 365076 480956
rect 230532 480916 365076 480944
rect 230532 480904 230538 480916
rect 365070 480904 365076 480916
rect 365128 480904 365134 480956
rect 296898 480156 296904 480208
rect 296956 480196 296962 480208
rect 358630 480196 358636 480208
rect 296956 480168 358636 480196
rect 296956 480156 296962 480168
rect 358630 480156 358636 480168
rect 358688 480156 358694 480208
rect 295426 480088 295432 480140
rect 295484 480128 295490 480140
rect 362678 480128 362684 480140
rect 295484 480100 362684 480128
rect 295484 480088 295490 480100
rect 362678 480088 362684 480100
rect 362736 480088 362742 480140
rect 295334 480020 295340 480072
rect 295392 480060 295398 480072
rect 364150 480060 364156 480072
rect 295392 480032 364156 480060
rect 295392 480020 295398 480032
rect 364150 480020 364156 480032
rect 364208 480020 364214 480072
rect 295518 479952 295524 480004
rect 295576 479992 295582 480004
rect 366910 479992 366916 480004
rect 295576 479964 366916 479992
rect 295576 479952 295582 479964
rect 366910 479952 366916 479964
rect 366968 479952 366974 480004
rect 294138 479884 294144 479936
rect 294196 479924 294202 479936
rect 365622 479924 365628 479936
rect 294196 479896 365628 479924
rect 294196 479884 294202 479896
rect 365622 479884 365628 479896
rect 365680 479884 365686 479936
rect 296806 479816 296812 479868
rect 296864 479856 296870 479868
rect 369578 479856 369584 479868
rect 296864 479828 369584 479856
rect 296864 479816 296870 479828
rect 369578 479816 369584 479828
rect 369636 479816 369642 479868
rect 298278 479748 298284 479800
rect 298336 479788 298342 479800
rect 379514 479788 379520 479800
rect 298336 479760 379520 479788
rect 298336 479748 298342 479760
rect 379514 479748 379520 479760
rect 379572 479748 379578 479800
rect 287238 479680 287244 479732
rect 287296 479720 287302 479732
rect 373718 479720 373724 479732
rect 287296 479692 373724 479720
rect 287296 479680 287302 479692
rect 373718 479680 373724 479692
rect 373776 479680 373782 479732
rect 284478 479612 284484 479664
rect 284536 479652 284542 479664
rect 377398 479652 377404 479664
rect 284536 479624 377404 479652
rect 284536 479612 284542 479624
rect 377398 479612 377404 479624
rect 377456 479612 377462 479664
rect 178218 479544 178224 479596
rect 178276 479584 178282 479596
rect 210602 479584 210608 479596
rect 178276 479556 210608 479584
rect 178276 479544 178282 479556
rect 210602 479544 210608 479556
rect 210660 479544 210666 479596
rect 252738 479544 252744 479596
rect 252796 479584 252802 479596
rect 374822 479584 374828 479596
rect 252796 479556 374828 479584
rect 252796 479544 252802 479556
rect 374822 479544 374828 479556
rect 374880 479544 374886 479596
rect 161750 479476 161756 479528
rect 161808 479516 161814 479528
rect 216030 479516 216036 479528
rect 161808 479488 216036 479516
rect 161808 479476 161814 479488
rect 216030 479476 216036 479488
rect 216088 479476 216094 479528
rect 244550 479476 244556 479528
rect 244608 479516 244614 479528
rect 369118 479516 369124 479528
rect 244608 479488 369124 479516
rect 244608 479476 244614 479488
rect 369118 479476 369124 479488
rect 369176 479476 369182 479528
rect 256786 478252 256792 478304
rect 256844 478292 256850 478304
rect 361298 478292 361304 478304
rect 256844 478264 361304 478292
rect 256844 478252 256850 478264
rect 361298 478252 361304 478264
rect 361356 478252 361362 478304
rect 252646 478184 252652 478236
rect 252704 478224 252710 478236
rect 369394 478224 369400 478236
rect 252704 478196 369400 478224
rect 252704 478184 252710 478196
rect 369394 478184 369400 478196
rect 369452 478184 369458 478236
rect 146386 478116 146392 478168
rect 146444 478156 146450 478168
rect 211890 478156 211896 478168
rect 146444 478128 211896 478156
rect 146444 478116 146450 478128
rect 211890 478116 211896 478128
rect 211948 478116 211954 478168
rect 244458 478116 244464 478168
rect 244516 478156 244522 478168
rect 374638 478156 374644 478168
rect 244516 478128 374644 478156
rect 244516 478116 244522 478128
rect 374638 478116 374644 478128
rect 374696 478116 374702 478168
rect 292666 477436 292672 477488
rect 292724 477476 292730 477488
rect 357158 477476 357164 477488
rect 292724 477448 357164 477476
rect 292724 477436 292730 477448
rect 357158 477436 357164 477448
rect 357216 477436 357222 477488
rect 294046 477368 294052 477420
rect 294104 477408 294110 477420
rect 368382 477408 368388 477420
rect 294104 477380 368388 477408
rect 294104 477368 294110 477380
rect 368382 477368 368388 477380
rect 368440 477368 368446 477420
rect 293954 477300 293960 477352
rect 294012 477340 294018 477352
rect 371142 477340 371148 477352
rect 294012 477312 371148 477340
rect 294012 477300 294018 477312
rect 371142 477300 371148 477312
rect 371200 477300 371206 477352
rect 291378 477232 291384 477284
rect 291436 477272 291442 477284
rect 374454 477272 374460 477284
rect 291436 477244 374460 477272
rect 291436 477232 291442 477244
rect 374454 477232 374460 477244
rect 374512 477232 374518 477284
rect 291286 477164 291292 477216
rect 291344 477204 291350 477216
rect 376478 477204 376484 477216
rect 291344 477176 376484 477204
rect 291344 477164 291350 477176
rect 376478 477164 376484 477176
rect 376536 477164 376542 477216
rect 285950 477096 285956 477148
rect 286008 477136 286014 477148
rect 371786 477136 371792 477148
rect 286008 477108 371792 477136
rect 286008 477096 286014 477108
rect 371786 477096 371792 477108
rect 371844 477096 371850 477148
rect 281626 477028 281632 477080
rect 281684 477068 281690 477080
rect 368290 477068 368296 477080
rect 281684 477040 368296 477068
rect 281684 477028 281690 477040
rect 368290 477028 368296 477040
rect 368348 477028 368354 477080
rect 289998 476960 290004 477012
rect 290056 477000 290062 477012
rect 377214 477000 377220 477012
rect 290056 476972 377220 477000
rect 290056 476960 290062 476972
rect 377214 476960 377220 476972
rect 377272 476960 377278 477012
rect 256694 476892 256700 476944
rect 256752 476932 256758 476944
rect 365346 476932 365352 476944
rect 256752 476904 365352 476932
rect 256752 476892 256758 476904
rect 365346 476892 365352 476904
rect 365404 476892 365410 476944
rect 244366 476824 244372 476876
rect 244424 476864 244430 476876
rect 373258 476864 373264 476876
rect 244424 476836 373264 476864
rect 244424 476824 244430 476836
rect 373258 476824 373264 476836
rect 373316 476824 373322 476876
rect 158806 476756 158812 476808
rect 158864 476796 158870 476808
rect 203610 476796 203616 476808
rect 158864 476768 203616 476796
rect 158864 476756 158870 476768
rect 203610 476756 203616 476768
rect 203668 476756 203674 476808
rect 226518 476756 226524 476808
rect 226576 476796 226582 476808
rect 378778 476796 378784 476808
rect 226576 476768 378784 476796
rect 226576 476756 226582 476768
rect 378778 476756 378784 476768
rect 378836 476756 378842 476808
rect 262306 475464 262312 475516
rect 262364 475504 262370 475516
rect 379238 475504 379244 475516
rect 262364 475476 379244 475504
rect 262364 475464 262370 475476
rect 379238 475464 379244 475476
rect 379296 475464 379302 475516
rect 252554 475396 252560 475448
rect 252612 475436 252618 475448
rect 374914 475436 374920 475448
rect 252612 475408 374920 475436
rect 252612 475396 252618 475408
rect 374914 475396 374920 475408
rect 374972 475396 374978 475448
rect 62758 475328 62764 475380
rect 62816 475368 62822 475380
rect 199378 475368 199384 475380
rect 62816 475340 199384 475368
rect 62816 475328 62822 475340
rect 199378 475328 199384 475340
rect 199436 475328 199442 475380
rect 227898 475328 227904 475380
rect 227956 475368 227962 475380
rect 367738 475368 367744 475380
rect 227956 475340 367744 475368
rect 227956 475328 227962 475340
rect 367738 475328 367744 475340
rect 367796 475328 367802 475380
rect 289906 474580 289912 474632
rect 289964 474620 289970 474632
rect 373166 474620 373172 474632
rect 289964 474592 373172 474620
rect 289964 474580 289970 474592
rect 373166 474580 373172 474592
rect 373224 474580 373230 474632
rect 267826 474512 267832 474564
rect 267884 474552 267890 474564
rect 359642 474552 359648 474564
rect 267884 474524 359648 474552
rect 267884 474512 267890 474524
rect 359642 474512 359648 474524
rect 359700 474512 359706 474564
rect 270678 474444 270684 474496
rect 270736 474484 270742 474496
rect 362770 474484 362776 474496
rect 270736 474456 362776 474484
rect 270736 474444 270742 474456
rect 362770 474444 362776 474456
rect 362828 474444 362834 474496
rect 267918 474376 267924 474428
rect 267976 474416 267982 474428
rect 361390 474416 361396 474428
rect 267976 474388 361396 474416
rect 267976 474376 267982 474388
rect 361390 474376 361396 474388
rect 361448 474376 361454 474428
rect 270586 474308 270592 474360
rect 270644 474348 270650 474360
rect 364886 474348 364892 474360
rect 270644 474320 364892 474348
rect 270644 474308 270650 474320
rect 364886 474308 364892 474320
rect 364944 474308 364950 474360
rect 269298 474240 269304 474292
rect 269356 474280 269362 474292
rect 369670 474280 369676 474292
rect 269356 474252 369676 474280
rect 269356 474240 269362 474252
rect 369670 474240 369676 474252
rect 369728 474240 369734 474292
rect 269206 474172 269212 474224
rect 269264 474212 269270 474224
rect 372430 474212 372436 474224
rect 269264 474184 372436 474212
rect 269264 474172 269270 474184
rect 372430 474172 372436 474184
rect 372488 474172 372494 474224
rect 259638 474104 259644 474156
rect 259696 474144 259702 474156
rect 372246 474144 372252 474156
rect 259696 474116 372252 474144
rect 259696 474104 259702 474116
rect 372246 474104 372252 474116
rect 372304 474104 372310 474156
rect 244274 474036 244280 474088
rect 244332 474076 244338 474088
rect 358446 474076 358452 474088
rect 244332 474048 358452 474076
rect 244332 474036 244338 474048
rect 358446 474036 358452 474048
rect 358504 474036 358510 474088
rect 161658 473968 161664 474020
rect 161716 474008 161722 474020
rect 213178 474008 213184 474020
rect 161716 473980 213184 474008
rect 161716 473968 161722 473980
rect 213178 473968 213184 473980
rect 213236 473968 213242 474020
rect 237466 473968 237472 474020
rect 237524 474008 237530 474020
rect 372062 474008 372068 474020
rect 237524 473980 372068 474008
rect 237524 473968 237530 473980
rect 372062 473968 372068 473980
rect 372120 473968 372126 474020
rect 185026 472744 185032 472796
rect 185084 472784 185090 472796
rect 210694 472784 210700 472796
rect 185084 472756 210700 472784
rect 185084 472744 185090 472756
rect 210694 472744 210700 472756
rect 210752 472744 210758 472796
rect 258258 472744 258264 472796
rect 258316 472784 258322 472796
rect 373534 472784 373540 472796
rect 258316 472756 373540 472784
rect 258316 472744 258322 472756
rect 373534 472744 373540 472756
rect 373592 472744 373598 472796
rect 178126 472676 178132 472728
rect 178184 472716 178190 472728
rect 205082 472716 205088 472728
rect 178184 472688 205088 472716
rect 178184 472676 178190 472688
rect 205082 472676 205088 472688
rect 205140 472676 205146 472728
rect 245746 472676 245752 472728
rect 245804 472716 245810 472728
rect 361114 472716 361120 472728
rect 245804 472688 361120 472716
rect 245804 472676 245810 472688
rect 361114 472676 361120 472688
rect 361172 472676 361178 472728
rect 3602 472608 3608 472660
rect 3660 472648 3666 472660
rect 307018 472648 307024 472660
rect 3660 472620 307024 472648
rect 3660 472608 3666 472620
rect 307018 472608 307024 472620
rect 307076 472608 307082 472660
rect 3510 471928 3516 471980
rect 3568 471968 3574 471980
rect 429194 471968 429200 471980
rect 3568 471940 429200 471968
rect 3568 471928 3574 471940
rect 429194 471928 429200 471940
rect 429252 471928 429258 471980
rect 273438 471860 273444 471912
rect 273496 471900 273502 471912
rect 359734 471900 359740 471912
rect 273496 471872 359740 471900
rect 273496 471860 273502 471872
rect 359734 471860 359740 471872
rect 359792 471860 359798 471912
rect 276198 471792 276204 471844
rect 276256 471832 276262 471844
rect 364242 471832 364248 471844
rect 276256 471804 364248 471832
rect 276256 471792 276262 471804
rect 364242 471792 364248 471804
rect 364300 471792 364306 471844
rect 277578 471724 277584 471776
rect 277636 471764 277642 471776
rect 369026 471764 369032 471776
rect 277636 471736 369032 471764
rect 277636 471724 277642 471736
rect 369026 471724 369032 471736
rect 369084 471724 369090 471776
rect 274910 471656 274916 471708
rect 274968 471696 274974 471708
rect 367646 471696 367652 471708
rect 274968 471668 367652 471696
rect 274968 471656 274974 471668
rect 367646 471656 367652 471668
rect 367704 471656 367710 471708
rect 284386 471588 284392 471640
rect 284444 471628 284450 471640
rect 377674 471628 377680 471640
rect 284444 471600 377680 471628
rect 284444 471588 284450 471600
rect 377674 471588 377680 471600
rect 377732 471588 377738 471640
rect 267734 471520 267740 471572
rect 267792 471560 267798 471572
rect 361482 471560 361488 471572
rect 267792 471532 361488 471560
rect 267792 471520 267798 471532
rect 361482 471520 361488 471532
rect 361540 471520 361546 471572
rect 272058 471452 272064 471504
rect 272116 471492 272122 471504
rect 367002 471492 367008 471504
rect 272116 471464 367008 471492
rect 272116 471452 272122 471464
rect 367002 471452 367008 471464
rect 367060 471452 367066 471504
rect 273346 471384 273352 471436
rect 273404 471424 273410 471436
rect 377490 471424 377496 471436
rect 273404 471396 377496 471424
rect 273404 471384 273410 471396
rect 377490 471384 377496 471396
rect 377548 471384 377554 471436
rect 176838 471316 176844 471368
rect 176896 471356 176902 471368
rect 206554 471356 206560 471368
rect 176896 471328 206560 471356
rect 176896 471316 176902 471328
rect 206554 471316 206560 471328
rect 206612 471316 206618 471368
rect 259546 471316 259552 471368
rect 259604 471356 259610 471368
rect 370866 471356 370872 471368
rect 259604 471328 370872 471356
rect 259604 471316 259610 471328
rect 370866 471316 370872 471328
rect 370924 471316 370930 471368
rect 164418 471248 164424 471300
rect 164476 471288 164482 471300
rect 211982 471288 211988 471300
rect 164476 471260 211988 471288
rect 164476 471248 164482 471260
rect 211982 471248 211988 471260
rect 212040 471248 212046 471300
rect 251358 471248 251364 471300
rect 251416 471288 251422 471300
rect 363966 471288 363972 471300
rect 251416 471260 363972 471288
rect 251416 471248 251422 471260
rect 363966 471248 363972 471260
rect 364024 471248 364030 471300
rect 284294 470024 284300 470076
rect 284352 470064 284358 470076
rect 377766 470064 377772 470076
rect 284352 470036 377772 470064
rect 284352 470024 284358 470036
rect 377766 470024 377772 470036
rect 377824 470024 377830 470076
rect 251266 469956 251272 470008
rect 251324 469996 251330 470008
rect 362402 469996 362408 470008
rect 251324 469968 362408 469996
rect 251324 469956 251330 469968
rect 362402 469956 362408 469968
rect 362460 469956 362466 470008
rect 176746 469888 176752 469940
rect 176804 469928 176810 469940
rect 212166 469928 212172 469940
rect 176804 469900 212172 469928
rect 176804 469888 176810 469900
rect 212166 469888 212172 469900
rect 212224 469888 212230 469940
rect 241606 469888 241612 469940
rect 241664 469928 241670 469940
rect 365162 469928 365168 469940
rect 241664 469900 365168 469928
rect 241664 469888 241670 469900
rect 365162 469888 365168 469900
rect 365220 469888 365226 469940
rect 4798 469820 4804 469872
rect 4856 469860 4862 469872
rect 391934 469860 391940 469872
rect 4856 469832 391940 469860
rect 4856 469820 4862 469832
rect 391934 469820 391940 469832
rect 391992 469820 391998 469872
rect 48130 469140 48136 469192
rect 48188 469180 48194 469192
rect 72418 469180 72424 469192
rect 48188 469152 72424 469180
rect 48188 469140 48194 469152
rect 72418 469140 72424 469152
rect 72476 469140 72482 469192
rect 285858 469140 285864 469192
rect 285916 469180 285922 469192
rect 370406 469180 370412 469192
rect 285916 469152 370412 469180
rect 285916 469140 285922 469152
rect 370406 469140 370412 469152
rect 370464 469140 370470 469192
rect 42610 469072 42616 469124
rect 42668 469112 42674 469124
rect 67818 469112 67824 469124
rect 42668 469084 67824 469112
rect 42668 469072 42674 469084
rect 67818 469072 67824 469084
rect 67876 469072 67882 469124
rect 266446 469072 266452 469124
rect 266504 469112 266510 469124
rect 360746 469112 360752 469124
rect 266504 469084 360752 469112
rect 266504 469072 266510 469084
rect 360746 469072 360752 469084
rect 360804 469072 360810 469124
rect 42518 469004 42524 469056
rect 42576 469044 42582 469056
rect 70578 469044 70584 469056
rect 42576 469016 70584 469044
rect 42576 469004 42582 469016
rect 70578 469004 70584 469016
rect 70636 469004 70642 469056
rect 276106 469004 276112 469056
rect 276164 469044 276170 469056
rect 375098 469044 375104 469056
rect 276164 469016 375104 469044
rect 276164 469004 276170 469016
rect 375098 469004 375104 469016
rect 375156 469004 375162 469056
rect 42426 468936 42432 468988
rect 42484 468976 42490 468988
rect 94038 468976 94044 468988
rect 42484 468948 94044 468976
rect 42484 468936 42490 468948
rect 94038 468936 94044 468948
rect 94096 468936 94102 468988
rect 259454 468936 259460 468988
rect 259512 468976 259518 468988
rect 362494 468976 362500 468988
rect 259512 468948 362500 468976
rect 259512 468936 259518 468948
rect 362494 468936 362500 468948
rect 362552 468936 362558 468988
rect 46198 468868 46204 468920
rect 46256 468908 46262 468920
rect 104986 468908 104992 468920
rect 46256 468880 104992 468908
rect 46256 468868 46262 468880
rect 104986 468868 104992 468880
rect 105044 468868 105050 468920
rect 254026 468868 254032 468920
rect 254084 468908 254090 468920
rect 362586 468908 362592 468920
rect 254084 468880 362592 468908
rect 254084 468868 254090 468880
rect 362586 468868 362592 468880
rect 362644 468868 362650 468920
rect 43530 468800 43536 468852
rect 43588 468840 43594 468852
rect 103606 468840 103612 468852
rect 43588 468812 103612 468840
rect 43588 468800 43594 468812
rect 103606 468800 103612 468812
rect 103664 468800 103670 468852
rect 255314 468800 255320 468852
rect 255372 468840 255378 468852
rect 365438 468840 365444 468852
rect 255372 468812 365444 468840
rect 255372 468800 255378 468812
rect 365438 468800 365444 468812
rect 365496 468800 365502 468852
rect 42150 468732 42156 468784
rect 42208 468772 42214 468784
rect 102226 468772 102232 468784
rect 42208 468744 102232 468772
rect 42208 468732 42214 468744
rect 102226 468732 102232 468744
rect 102284 468732 102290 468784
rect 254118 468732 254124 468784
rect 254176 468772 254182 468784
rect 368198 468772 368204 468784
rect 254176 468744 368204 468772
rect 254176 468732 254182 468744
rect 368198 468732 368204 468744
rect 368256 468732 368262 468784
rect 45370 468664 45376 468716
rect 45428 468704 45434 468716
rect 106366 468704 106372 468716
rect 45428 468676 106372 468704
rect 45428 468664 45434 468676
rect 106366 468664 106372 468676
rect 106424 468664 106430 468716
rect 255498 468664 255504 468716
rect 255556 468704 255562 468716
rect 373626 468704 373632 468716
rect 255556 468676 373632 468704
rect 255556 468664 255562 468676
rect 373626 468664 373632 468676
rect 373684 468664 373690 468716
rect 45278 468596 45284 468648
rect 45336 468636 45342 468648
rect 106458 468636 106464 468648
rect 45336 468608 106464 468636
rect 45336 468596 45342 468608
rect 106458 468596 106464 468608
rect 106516 468596 106522 468648
rect 255406 468596 255412 468648
rect 255464 468636 255470 468648
rect 376294 468636 376300 468648
rect 255464 468608 376300 468636
rect 255464 468596 255470 468608
rect 376294 468596 376300 468608
rect 376352 468596 376358 468648
rect 43438 468528 43444 468580
rect 43496 468568 43502 468580
rect 105078 468568 105084 468580
rect 43496 468540 105084 468568
rect 43496 468528 43502 468540
rect 105078 468528 105084 468540
rect 105136 468528 105142 468580
rect 174078 468528 174084 468580
rect 174136 468568 174142 468580
rect 214650 468568 214656 468580
rect 174136 468540 214656 468568
rect 174136 468528 174142 468540
rect 214650 468528 214656 468540
rect 214708 468528 214714 468580
rect 247126 468528 247132 468580
rect 247184 468568 247190 468580
rect 378962 468568 378968 468580
rect 247184 468540 378968 468568
rect 247184 468528 247190 468540
rect 378962 468528 378968 468540
rect 379020 468528 379026 468580
rect 18598 468460 18604 468512
rect 18656 468500 18662 468512
rect 378134 468500 378140 468512
rect 18656 468472 378140 468500
rect 18656 468460 18662 468472
rect 378134 468460 378140 468472
rect 378192 468460 378198 468512
rect 44082 468392 44088 468444
rect 44140 468432 44146 468444
rect 66346 468432 66352 468444
rect 44140 468404 66352 468432
rect 44140 468392 44146 468404
rect 66346 468392 66352 468404
rect 66404 468392 66410 468444
rect 288618 468392 288624 468444
rect 288676 468432 288682 468444
rect 367554 468432 367560 468444
rect 288676 468404 367560 468432
rect 288676 468392 288682 468404
rect 367554 468392 367560 468404
rect 367612 468392 367618 468444
rect 175458 467236 175464 467288
rect 175516 467276 175522 467288
rect 200850 467276 200856 467288
rect 175516 467248 200856 467276
rect 175516 467236 175522 467248
rect 200850 467236 200856 467248
rect 200908 467236 200914 467288
rect 175366 467168 175372 467220
rect 175424 467208 175430 467220
rect 202230 467208 202236 467220
rect 175424 467180 202236 467208
rect 175424 467168 175430 467180
rect 202230 467168 202236 467180
rect 202288 467168 202294 467220
rect 57514 467100 57520 467152
rect 57572 467140 57578 467152
rect 111886 467140 111892 467152
rect 57572 467112 111892 467140
rect 57572 467100 57578 467112
rect 111886 467100 111892 467112
rect 111944 467100 111950 467152
rect 162946 467100 162952 467152
rect 163004 467140 163010 467152
rect 209130 467140 209136 467152
rect 163004 467112 209136 467140
rect 163004 467100 163010 467112
rect 209130 467100 209136 467112
rect 209188 467100 209194 467152
rect 209222 467100 209228 467152
rect 209280 467140 209286 467152
rect 217778 467140 217784 467152
rect 209280 467112 217784 467140
rect 209280 467100 209286 467112
rect 217778 467100 217784 467112
rect 217836 467100 217842 467152
rect 227806 467100 227812 467152
rect 227864 467140 227870 467152
rect 371878 467140 371884 467152
rect 227864 467112 371884 467140
rect 227864 467100 227870 467112
rect 371878 467100 371884 467112
rect 371936 467100 371942 467152
rect 45186 466352 45192 466404
rect 45244 466392 45250 466404
rect 68278 466392 68284 466404
rect 45244 466364 68284 466392
rect 45244 466352 45250 466364
rect 68278 466352 68284 466364
rect 68336 466352 68342 466404
rect 190638 466352 190644 466404
rect 190696 466392 190702 466404
rect 212902 466392 212908 466404
rect 190696 466364 212908 466392
rect 190696 466352 190702 466364
rect 212902 466352 212908 466364
rect 212960 466352 212966 466404
rect 280338 466352 280344 466404
rect 280396 466392 280402 466404
rect 357250 466392 357256 466404
rect 280396 466364 357256 466392
rect 280396 466352 280402 466364
rect 357250 466352 357256 466364
rect 357308 466352 357314 466404
rect 45094 466284 45100 466336
rect 45152 466324 45158 466336
rect 68370 466324 68376 466336
rect 45152 466296 68376 466324
rect 45152 466284 45158 466296
rect 68370 466284 68376 466296
rect 68428 466284 68434 466336
rect 176654 466284 176660 466336
rect 176712 466324 176718 466336
rect 209314 466324 209320 466336
rect 176712 466296 209320 466324
rect 176712 466284 176718 466296
rect 209314 466284 209320 466296
rect 209372 466284 209378 466336
rect 298186 466284 298192 466336
rect 298244 466324 298250 466336
rect 376570 466324 376576 466336
rect 298244 466296 376576 466324
rect 298244 466284 298250 466296
rect 376570 466284 376576 466296
rect 376628 466284 376634 466336
rect 52086 466216 52092 466268
rect 52144 466256 52150 466268
rect 82814 466256 82820 466268
rect 52144 466228 82820 466256
rect 52144 466216 52150 466228
rect 82814 466216 82820 466228
rect 82872 466216 82878 466268
rect 173986 466216 173992 466268
rect 174044 466256 174050 466268
rect 207842 466256 207848 466268
rect 174044 466228 207848 466256
rect 174044 466216 174050 466228
rect 207842 466216 207848 466228
rect 207900 466216 207906 466268
rect 289814 466216 289820 466268
rect 289872 466256 289878 466268
rect 373074 466256 373080 466268
rect 289872 466228 373080 466256
rect 289872 466216 289878 466228
rect 373074 466216 373080 466228
rect 373132 466216 373138 466268
rect 50706 466148 50712 466200
rect 50764 466188 50770 466200
rect 82998 466188 83004 466200
rect 50764 466160 83004 466188
rect 50764 466148 50770 466160
rect 82998 466148 83004 466160
rect 83056 466148 83062 466200
rect 140774 466148 140780 466200
rect 140832 466188 140838 466200
rect 197814 466188 197820 466200
rect 140832 466160 197820 466188
rect 140832 466148 140838 466160
rect 197814 466148 197820 466160
rect 197872 466148 197878 466200
rect 271966 466148 271972 466200
rect 272024 466188 272030 466200
rect 358722 466188 358728 466200
rect 272024 466160 358728 466188
rect 272024 466148 272030 466160
rect 358722 466148 358728 466160
rect 358780 466148 358786 466200
rect 49510 466080 49516 466132
rect 49568 466120 49574 466132
rect 82906 466120 82912 466132
rect 49568 466092 82912 466120
rect 49568 466080 49574 466092
rect 82906 466080 82912 466092
rect 82964 466080 82970 466132
rect 139394 466080 139400 466132
rect 139452 466120 139458 466132
rect 197078 466120 197084 466132
rect 139452 466092 197084 466120
rect 139452 466080 139458 466092
rect 197078 466080 197084 466092
rect 197136 466080 197142 466132
rect 263778 466080 263784 466132
rect 263836 466120 263842 466132
rect 356882 466120 356888 466132
rect 263836 466092 356888 466120
rect 263836 466080 263842 466092
rect 356882 466080 356888 466092
rect 356940 466080 356946 466132
rect 57790 466012 57796 466064
rect 57848 466052 57854 466064
rect 102318 466052 102324 466064
rect 57848 466024 102324 466052
rect 57848 466012 57854 466024
rect 102318 466012 102324 466024
rect 102376 466012 102382 466064
rect 140866 466012 140872 466064
rect 140924 466052 140930 466064
rect 200482 466052 200488 466064
rect 140924 466024 200488 466052
rect 140924 466012 140930 466024
rect 200482 466012 200488 466024
rect 200540 466012 200546 466064
rect 263686 466012 263692 466064
rect 263744 466052 263750 466064
rect 366818 466052 366824 466064
rect 263744 466024 366824 466052
rect 263744 466012 263750 466024
rect 366818 466012 366824 466024
rect 366876 466012 366882 466064
rect 54570 465944 54576 465996
rect 54628 465984 54634 465996
rect 100938 465984 100944 465996
rect 54628 465956 100944 465984
rect 54628 465944 54634 465956
rect 100938 465944 100944 465956
rect 100996 465944 101002 465996
rect 140958 465944 140964 465996
rect 141016 465984 141022 465996
rect 201770 465984 201776 465996
rect 141016 465956 201776 465984
rect 141016 465944 141022 465956
rect 201770 465944 201776 465956
rect 201828 465944 201834 465996
rect 265250 465944 265256 465996
rect 265308 465984 265314 465996
rect 372338 465984 372344 465996
rect 265308 465956 372344 465984
rect 265308 465944 265314 465956
rect 372338 465944 372344 465956
rect 372396 465944 372402 465996
rect 53098 465876 53104 465928
rect 53156 465916 53162 465928
rect 100846 465916 100852 465928
rect 53156 465888 100852 465916
rect 53156 465876 53162 465888
rect 100846 465876 100852 465888
rect 100904 465876 100910 465928
rect 141050 465876 141056 465928
rect 141108 465916 141114 465928
rect 203334 465916 203340 465928
rect 141108 465888 203340 465916
rect 141108 465876 141114 465888
rect 203334 465876 203340 465888
rect 203392 465876 203398 465928
rect 265158 465876 265164 465928
rect 265216 465916 265222 465928
rect 375006 465916 375012 465928
rect 265216 465888 375012 465916
rect 265216 465876 265222 465888
rect 375006 465876 375012 465888
rect 375064 465876 375070 465928
rect 57422 465808 57428 465860
rect 57480 465848 57486 465860
rect 113358 465848 113364 465860
rect 57480 465820 113364 465848
rect 57480 465808 57486 465820
rect 113358 465808 113364 465820
rect 113416 465808 113422 465860
rect 139486 465808 139492 465860
rect 139544 465848 139550 465860
rect 204530 465848 204536 465860
rect 139544 465820 204536 465848
rect 139544 465808 139550 465820
rect 204530 465808 204536 465820
rect 204588 465808 204594 465860
rect 260834 465808 260840 465860
rect 260892 465848 260898 465860
rect 376386 465848 376392 465860
rect 260892 465820 376392 465848
rect 260892 465808 260898 465820
rect 376386 465808 376392 465820
rect 376444 465808 376450 465860
rect 50246 465740 50252 465792
rect 50304 465780 50310 465792
rect 98178 465780 98184 465792
rect 50304 465752 98184 465780
rect 50304 465740 50310 465752
rect 98178 465740 98184 465752
rect 98236 465740 98242 465792
rect 107838 465740 107844 465792
rect 107896 465780 107902 465792
rect 204346 465780 204352 465792
rect 107896 465752 204352 465780
rect 107896 465740 107902 465752
rect 204346 465740 204352 465752
rect 204404 465740 204410 465792
rect 226334 465740 226340 465792
rect 226392 465780 226398 465792
rect 361022 465780 361028 465792
rect 226392 465752 361028 465780
rect 226392 465740 226398 465752
rect 361022 465740 361028 465752
rect 361080 465740 361086 465792
rect 51626 465672 51632 465724
rect 51684 465712 51690 465724
rect 99466 465712 99472 465724
rect 51684 465684 99472 465712
rect 51684 465672 51690 465684
rect 99466 465672 99472 465684
rect 99524 465672 99530 465724
rect 109034 465672 109040 465724
rect 109092 465712 109098 465724
rect 205634 465712 205640 465724
rect 109092 465684 205640 465712
rect 109092 465672 109098 465684
rect 205634 465672 205640 465684
rect 205692 465672 205698 465724
rect 227714 465672 227720 465724
rect 227772 465712 227778 465724
rect 370498 465712 370504 465724
rect 227772 465684 370504 465712
rect 227772 465672 227778 465684
rect 370498 465672 370504 465684
rect 370556 465672 370562 465724
rect 44726 465604 44732 465656
rect 44784 465644 44790 465656
rect 65058 465644 65064 465656
rect 44784 465616 65064 465644
rect 44784 465604 44790 465616
rect 65058 465604 65064 465616
rect 65116 465604 65122 465656
rect 187878 465604 187884 465656
rect 187936 465644 187942 465656
rect 206646 465644 206652 465656
rect 187936 465616 206652 465644
rect 187936 465604 187942 465616
rect 206646 465604 206652 465616
rect 206704 465604 206710 465656
rect 44818 465536 44824 465588
rect 44876 465576 44882 465588
rect 64966 465576 64972 465588
rect 44876 465548 64972 465576
rect 44876 465536 44882 465548
rect 64966 465536 64972 465548
rect 65024 465536 65030 465588
rect 182358 465536 182364 465588
rect 182416 465576 182422 465588
rect 200942 465576 200948 465588
rect 182416 465548 200948 465576
rect 182416 465536 182422 465548
rect 200942 465536 200948 465548
rect 201000 465536 201006 465588
rect 44910 465468 44916 465520
rect 44968 465508 44974 465520
rect 64874 465508 64880 465520
rect 44968 465480 64880 465508
rect 44968 465468 44974 465480
rect 64874 465468 64880 465480
rect 64932 465468 64938 465520
rect 192110 465468 192116 465520
rect 192168 465508 192174 465520
rect 205358 465508 205364 465520
rect 192168 465480 205364 465508
rect 192168 465468 192174 465480
rect 205358 465468 205364 465480
rect 205416 465468 205422 465520
rect 287146 464448 287152 464500
rect 287204 464488 287210 464500
rect 370314 464488 370320 464500
rect 287204 464460 370320 464488
rect 287204 464448 287210 464460
rect 370314 464448 370320 464460
rect 370372 464448 370378 464500
rect 164234 464380 164240 464432
rect 164292 464420 164298 464432
rect 216122 464420 216128 464432
rect 164292 464392 216128 464420
rect 164292 464380 164298 464392
rect 216122 464380 216128 464392
rect 216180 464380 216186 464432
rect 274818 464380 274824 464432
rect 274876 464420 274882 464432
rect 364794 464420 364800 464432
rect 274876 464392 364800 464420
rect 274876 464380 274882 464392
rect 364794 464380 364800 464392
rect 364852 464380 364858 464432
rect 160186 464312 160192 464364
rect 160244 464352 160250 464364
rect 214558 464352 214564 464364
rect 160244 464324 214564 464352
rect 160244 464312 160250 464324
rect 214558 464312 214564 464324
rect 214616 464312 214622 464364
rect 285766 464312 285772 464364
rect 285824 464352 285830 464364
rect 377582 464352 377588 464364
rect 285824 464324 377588 464352
rect 285824 464312 285830 464324
rect 377582 464312 377588 464324
rect 377640 464312 377646 464364
rect 59906 463632 59912 463684
rect 59964 463672 59970 463684
rect 91186 463672 91192 463684
rect 59964 463644 91192 463672
rect 59964 463632 59970 463644
rect 91186 463632 91192 463644
rect 91244 463632 91250 463684
rect 190546 463632 190552 463684
rect 190604 463672 190610 463684
rect 214374 463672 214380 463684
rect 190604 463644 214380 463672
rect 190604 463632 190610 463644
rect 214374 463632 214380 463644
rect 214432 463632 214438 463684
rect 54938 463564 54944 463616
rect 54996 463604 55002 463616
rect 86954 463604 86960 463616
rect 54996 463576 86960 463604
rect 54996 463564 55002 463576
rect 86954 463564 86960 463576
rect 87012 463564 87018 463616
rect 190454 463564 190460 463616
rect 190512 463604 190518 463616
rect 217502 463604 217508 463616
rect 190512 463576 217508 463604
rect 190512 463564 190518 463576
rect 217502 463564 217508 463576
rect 217560 463564 217566 463616
rect 277486 463564 277492 463616
rect 277544 463604 277550 463616
rect 357342 463604 357348 463616
rect 277544 463576 357348 463604
rect 277544 463564 277550 463576
rect 357342 463564 357348 463576
rect 357400 463564 357406 463616
rect 49602 463496 49608 463548
rect 49660 463536 49666 463548
rect 81618 463536 81624 463548
rect 49660 463508 81624 463536
rect 49660 463496 49666 463508
rect 81618 463496 81624 463508
rect 81676 463496 81682 463548
rect 184934 463496 184940 463548
rect 184992 463536 184998 463548
rect 213270 463536 213276 463548
rect 184992 463508 213276 463536
rect 184992 463496 184998 463508
rect 213270 463496 213276 463508
rect 213328 463496 213334 463548
rect 288526 463496 288532 463548
rect 288584 463536 288590 463548
rect 368934 463536 368940 463548
rect 288584 463508 368940 463536
rect 288584 463496 288590 463508
rect 368934 463496 368940 463508
rect 368992 463496 368998 463548
rect 55950 463428 55956 463480
rect 56008 463468 56014 463480
rect 88610 463468 88616 463480
rect 56008 463440 88616 463468
rect 56008 463428 56014 463440
rect 88610 463428 88616 463440
rect 88668 463428 88674 463480
rect 183738 463428 183744 463480
rect 183796 463468 183802 463480
rect 212258 463468 212264 463480
rect 183796 463440 212264 463468
rect 183796 463428 183802 463440
rect 212258 463428 212264 463440
rect 212316 463428 212322 463480
rect 277394 463428 277400 463480
rect 277452 463468 277458 463480
rect 366266 463468 366272 463480
rect 277452 463440 366272 463468
rect 277452 463428 277458 463440
rect 366266 463428 366272 463440
rect 366324 463428 366330 463480
rect 51994 463360 52000 463412
rect 52052 463400 52058 463412
rect 85666 463400 85672 463412
rect 52052 463372 85672 463400
rect 52052 463360 52058 463372
rect 85666 463360 85672 463372
rect 85724 463360 85730 463412
rect 175274 463360 175280 463412
rect 175332 463400 175338 463412
rect 207934 463400 207940 463412
rect 175332 463372 207940 463400
rect 175332 463360 175338 463372
rect 207934 463360 207940 463372
rect 207992 463360 207998 463412
rect 276014 463360 276020 463412
rect 276072 463400 276078 463412
rect 371694 463400 371700 463412
rect 276072 463372 371700 463400
rect 276072 463360 276078 463372
rect 371694 463360 371700 463372
rect 371752 463360 371758 463412
rect 56226 463292 56232 463344
rect 56284 463332 56290 463344
rect 89806 463332 89812 463344
rect 56284 463304 89812 463332
rect 56284 463292 56290 463304
rect 89806 463292 89812 463304
rect 89864 463292 89870 463344
rect 180978 463292 180984 463344
rect 181036 463332 181042 463344
rect 216214 463332 216220 463344
rect 181036 463304 216220 463332
rect 181036 463292 181042 463304
rect 216214 463292 216220 463304
rect 216272 463292 216278 463344
rect 269114 463292 269120 463344
rect 269172 463332 269178 463344
rect 366174 463332 366180 463344
rect 269172 463304 366180 463332
rect 269172 463292 269178 463304
rect 366174 463292 366180 463304
rect 366232 463292 366238 463344
rect 54846 463224 54852 463276
rect 54904 463264 54910 463276
rect 88518 463264 88524 463276
rect 54904 463236 88524 463264
rect 54904 463224 54910 463236
rect 88518 463224 88524 463236
rect 88576 463224 88582 463276
rect 160094 463224 160100 463276
rect 160152 463264 160158 463276
rect 200758 463264 200764 463276
rect 160152 463236 200764 463264
rect 160152 463224 160158 463236
rect 200758 463224 200764 463236
rect 200816 463224 200822 463276
rect 263594 463224 263600 463276
rect 263652 463264 263658 463276
rect 363874 463264 363880 463276
rect 263652 463236 363880 463264
rect 263652 463224 263658 463236
rect 363874 463224 363880 463236
rect 363932 463224 363938 463276
rect 54754 463156 54760 463208
rect 54812 463196 54818 463208
rect 88426 463196 88432 463208
rect 54812 463168 88432 463196
rect 54812 463156 54818 463168
rect 88426 463156 88432 463168
rect 88484 463156 88490 463208
rect 168466 463156 168472 463208
rect 168524 463196 168530 463208
rect 210510 463196 210516 463208
rect 168524 463168 210516 463196
rect 168524 463156 168530 463168
rect 210510 463156 210516 463168
rect 210568 463156 210574 463208
rect 262214 463156 262220 463208
rect 262272 463196 262278 463208
rect 365530 463196 365536 463208
rect 262272 463168 365536 463196
rect 262272 463156 262278 463168
rect 365530 463156 365536 463168
rect 365588 463156 365594 463208
rect 53006 463088 53012 463140
rect 53064 463128 53070 463140
rect 87138 463128 87144 463140
rect 53064 463100 87144 463128
rect 53064 463088 53070 463100
rect 87138 463088 87144 463100
rect 87196 463088 87202 463140
rect 142338 463088 142344 463140
rect 142396 463128 142402 463140
rect 199102 463128 199108 463140
rect 142396 463100 199108 463128
rect 142396 463088 142402 463100
rect 199102 463088 199108 463100
rect 199160 463088 199166 463140
rect 241514 463088 241520 463140
rect 241572 463128 241578 463140
rect 358538 463128 358544 463140
rect 241572 463100 358544 463128
rect 241572 463088 241578 463100
rect 358538 463088 358544 463100
rect 358596 463088 358602 463140
rect 59078 463020 59084 463072
rect 59136 463060 59142 463072
rect 95418 463060 95424 463072
rect 59136 463032 95424 463060
rect 59136 463020 59142 463032
rect 95418 463020 95424 463032
rect 95476 463020 95482 463072
rect 142246 463020 142252 463072
rect 142304 463060 142310 463072
rect 207474 463060 207480 463072
rect 142304 463032 207480 463060
rect 142304 463020 142310 463032
rect 207474 463020 207480 463032
rect 207532 463020 207538 463072
rect 251174 463020 251180 463072
rect 251232 463060 251238 463072
rect 370774 463060 370780 463072
rect 251232 463032 370780 463060
rect 251232 463020 251238 463032
rect 370774 463020 370780 463032
rect 370832 463020 370838 463072
rect 52822 462952 52828 463004
rect 52880 462992 52886 463004
rect 100754 462992 100760 463004
rect 52880 462964 100760 462992
rect 52880 462952 52886 462964
rect 100754 462952 100760 462964
rect 100812 462952 100818 463004
rect 107746 462952 107752 463004
rect 107804 462992 107810 463004
rect 197630 462992 197636 463004
rect 107804 462964 197636 462992
rect 107804 462952 107810 462964
rect 197630 462952 197636 462964
rect 197688 462952 197694 463004
rect 240134 462952 240140 463004
rect 240192 462992 240198 463004
rect 361206 462992 361212 463004
rect 240192 462964 361212 462992
rect 240192 462952 240198 462964
rect 361206 462952 361212 462964
rect 361264 462952 361270 463004
rect 56042 462884 56048 462936
rect 56100 462924 56106 462936
rect 87046 462924 87052 462936
rect 56100 462896 87052 462924
rect 56100 462884 56106 462896
rect 87046 462884 87052 462896
rect 87104 462884 87110 462936
rect 180886 462884 180892 462936
rect 180944 462924 180950 462936
rect 203702 462924 203708 462936
rect 180944 462896 203708 462924
rect 180944 462884 180950 462896
rect 203702 462884 203708 462896
rect 203760 462884 203766 462936
rect 55858 462816 55864 462868
rect 55916 462856 55922 462868
rect 85574 462856 85580 462868
rect 55916 462828 85580 462856
rect 55916 462816 55922 462828
rect 85574 462816 85580 462828
rect 85632 462816 85638 462868
rect 187786 462816 187792 462868
rect 187844 462856 187850 462868
rect 205174 462856 205180 462868
rect 187844 462828 205180 462856
rect 187844 462816 187850 462828
rect 205174 462816 205180 462828
rect 205232 462816 205238 462868
rect 44634 462748 44640 462800
rect 44692 462788 44698 462800
rect 63678 462788 63684 462800
rect 44692 462760 63684 462788
rect 44692 462748 44698 462760
rect 63678 462748 63684 462760
rect 63736 462748 63742 462800
rect 193306 462748 193312 462800
rect 193364 462788 193370 462800
rect 206830 462788 206836 462800
rect 193364 462760 206836 462788
rect 193364 462748 193370 462760
rect 206830 462748 206836 462760
rect 206888 462748 206894 462800
rect 207014 462340 207020 462392
rect 207072 462380 207078 462392
rect 207290 462380 207296 462392
rect 207072 462352 207296 462380
rect 207072 462340 207078 462352
rect 207290 462340 207296 462352
rect 207348 462380 207354 462392
rect 217686 462380 217692 462392
rect 207348 462352 217692 462380
rect 207348 462340 207354 462352
rect 217686 462340 217692 462352
rect 217744 462340 217750 462392
rect 86218 462272 86224 462324
rect 86276 462312 86282 462324
rect 178310 462312 178316 462324
rect 86276 462284 178316 462312
rect 86276 462272 86282 462284
rect 178310 462272 178316 462284
rect 178368 462272 178374 462324
rect 180058 462272 180064 462324
rect 180116 462312 180122 462324
rect 199562 462312 199568 462324
rect 180116 462284 199568 462312
rect 180116 462272 180122 462284
rect 199562 462272 199568 462284
rect 199620 462272 199626 462324
rect 203150 462272 203156 462324
rect 203208 462312 203214 462324
rect 206278 462312 206284 462324
rect 203208 462284 206284 462312
rect 203208 462272 203214 462284
rect 206278 462272 206284 462284
rect 206336 462272 206342 462324
rect 192478 462204 192484 462256
rect 192536 462244 192542 462256
rect 210050 462244 210056 462256
rect 192536 462216 210056 462244
rect 192536 462204 192542 462216
rect 210050 462204 210056 462216
rect 210108 462204 210114 462256
rect 186406 462136 186412 462188
rect 186464 462176 186470 462188
rect 205266 462176 205272 462188
rect 186464 462148 205272 462176
rect 186464 462136 186470 462148
rect 205266 462136 205272 462148
rect 205324 462136 205330 462188
rect 191926 462068 191932 462120
rect 191984 462108 191990 462120
rect 215846 462108 215852 462120
rect 191984 462080 215852 462108
rect 191984 462068 191990 462080
rect 215846 462068 215852 462080
rect 215904 462068 215910 462120
rect 283006 462068 283012 462120
rect 283064 462108 283070 462120
rect 360838 462108 360844 462120
rect 283064 462080 360844 462108
rect 283064 462068 283070 462080
rect 360838 462068 360844 462080
rect 360896 462068 360902 462120
rect 192018 462000 192024 462052
rect 192076 462040 192082 462052
rect 218422 462040 218428 462052
rect 192076 462012 218428 462040
rect 192076 462000 192082 462012
rect 218422 462000 218428 462012
rect 218480 462000 218486 462052
rect 278774 462000 278780 462052
rect 278832 462040 278838 462052
rect 357894 462040 357900 462052
rect 278832 462012 357900 462040
rect 278832 462000 278838 462012
rect 357894 462000 357900 462012
rect 357952 462000 357958 462052
rect 182266 461932 182272 461984
rect 182324 461972 182330 461984
rect 209406 461972 209412 461984
rect 182324 461944 209412 461972
rect 182324 461932 182330 461944
rect 209406 461932 209412 461944
rect 209464 461932 209470 461984
rect 287054 461932 287060 461984
rect 287112 461972 287118 461984
rect 372522 461972 372528 461984
rect 287112 461944 372528 461972
rect 287112 461932 287118 461944
rect 372522 461932 372528 461944
rect 372580 461932 372586 461984
rect 182174 461864 182180 461916
rect 182232 461904 182238 461916
rect 211430 461904 211436 461916
rect 182232 461876 211436 461904
rect 182232 461864 182238 461876
rect 211430 461864 211436 461876
rect 211488 461864 211494 461916
rect 285674 461864 285680 461916
rect 285732 461904 285738 461916
rect 373994 461904 374000 461916
rect 285732 461876 374000 461904
rect 285732 461864 285738 461876
rect 373994 461864 374000 461876
rect 374052 461864 374058 461916
rect 511258 461864 511264 461916
rect 511316 461904 511322 461916
rect 517514 461904 517520 461916
rect 511316 461876 517520 461904
rect 511316 461864 511322 461876
rect 517514 461864 517520 461876
rect 517572 461864 517578 461916
rect 171226 461796 171232 461848
rect 171284 461836 171290 461848
rect 212074 461836 212080 461848
rect 171284 461808 212080 461836
rect 171284 461796 171290 461808
rect 212074 461796 212080 461808
rect 212132 461796 212138 461848
rect 271874 461796 271880 461848
rect 271932 461836 271938 461848
rect 363506 461836 363512 461848
rect 271932 461808 363512 461836
rect 271932 461796 271938 461808
rect 363506 461796 363512 461808
rect 363564 461796 363570 461848
rect 57330 461728 57336 461780
rect 57388 461768 57394 461780
rect 111978 461768 111984 461780
rect 57388 461740 111984 461768
rect 57388 461728 57394 461740
rect 111978 461728 111984 461740
rect 112036 461728 112042 461780
rect 165614 461728 165620 461780
rect 165672 461768 165678 461780
rect 218882 461768 218888 461780
rect 165672 461740 218888 461768
rect 165672 461728 165678 461740
rect 218882 461728 218888 461740
rect 218940 461728 218946 461780
rect 280246 461728 280252 461780
rect 280304 461768 280310 461780
rect 375742 461768 375748 461780
rect 280304 461740 375748 461768
rect 280304 461728 280310 461740
rect 375742 461728 375748 461740
rect 375800 461728 375806 461780
rect 62206 461660 62212 461712
rect 62264 461700 62270 461712
rect 199470 461700 199476 461712
rect 62264 461672 199476 461700
rect 62264 461660 62270 461672
rect 199470 461660 199476 461672
rect 199528 461660 199534 461712
rect 199562 461660 199568 461712
rect 199620 461700 199626 461712
rect 339678 461700 339684 461712
rect 199620 461672 339684 461700
rect 199620 461660 199626 461672
rect 339678 461660 339684 461672
rect 339736 461660 339742 461712
rect 47578 461592 47584 461644
rect 47636 461632 47642 461644
rect 207014 461632 207020 461644
rect 47636 461604 207020 461632
rect 47636 461592 47642 461604
rect 207014 461592 207020 461604
rect 207072 461592 207078 461644
rect 274726 461592 274732 461644
rect 274784 461632 274790 461644
rect 371050 461632 371056 461644
rect 274784 461604 371056 461632
rect 274784 461592 274790 461604
rect 371050 461592 371056 461604
rect 371108 461592 371114 461644
rect 339678 461048 339684 461100
rect 339736 461088 339742 461100
rect 360102 461088 360108 461100
rect 339736 461060 360108 461088
rect 339736 461048 339742 461060
rect 360102 461048 360108 461060
rect 360160 461088 360166 461100
rect 499850 461088 499856 461100
rect 360160 461060 499856 461088
rect 360160 461048 360166 461060
rect 499850 461048 499856 461060
rect 499908 461088 499914 461100
rect 500862 461088 500868 461100
rect 499908 461060 500868 461088
rect 499908 461048 499914 461060
rect 500862 461048 500868 461060
rect 500920 461048 500926 461100
rect 178310 460980 178316 461032
rect 178368 461020 178374 461032
rect 200574 461020 200580 461032
rect 178368 460992 200580 461020
rect 178368 460980 178374 460992
rect 200574 460980 200580 460992
rect 200632 461020 200638 461032
rect 338298 461020 338304 461032
rect 200632 460992 338304 461020
rect 200632 460980 200638 460992
rect 338298 460980 338304 460992
rect 338356 461020 338362 461032
rect 357066 461020 357072 461032
rect 338356 460992 357072 461020
rect 338356 460980 338362 460992
rect 357066 460980 357072 460992
rect 357124 461020 357130 461032
rect 498470 461020 498476 461032
rect 357124 460992 498476 461020
rect 357124 460980 357130 460992
rect 498470 460980 498476 460992
rect 498528 461020 498534 461032
rect 517790 461020 517796 461032
rect 498528 460992 517796 461020
rect 498528 460980 498534 460992
rect 517790 460980 517796 460992
rect 517848 460980 517854 461032
rect 190914 460912 190920 460964
rect 190972 460952 190978 460964
rect 207014 460952 207020 460964
rect 190972 460924 207020 460952
rect 190972 460912 190978 460924
rect 207014 460912 207020 460924
rect 207072 460912 207078 460964
rect 350994 460912 351000 460964
rect 351052 460952 351058 460964
rect 361574 460952 361580 460964
rect 351052 460924 361580 460952
rect 351052 460912 351058 460924
rect 361574 460912 361580 460924
rect 361632 460912 361638 460964
rect 500862 460912 500868 460964
rect 500920 460952 500926 460964
rect 517606 460952 517612 460964
rect 500920 460924 517612 460952
rect 500920 460912 500926 460924
rect 517606 460912 517612 460924
rect 517664 460912 517670 460964
rect 49234 460844 49240 460896
rect 49292 460884 49298 460896
rect 78858 460884 78864 460896
rect 49292 460856 78864 460884
rect 49292 460844 49298 460856
rect 78858 460844 78864 460856
rect 78916 460844 78922 460896
rect 183554 460844 183560 460896
rect 183612 460884 183618 460896
rect 202322 460884 202328 460896
rect 183612 460856 202328 460884
rect 183612 460844 183618 460856
rect 202322 460844 202328 460856
rect 202380 460844 202386 460896
rect 299474 460844 299480 460896
rect 299532 460884 299538 460896
rect 379422 460884 379428 460896
rect 299532 460856 379428 460884
rect 299532 460844 299538 460856
rect 379422 460844 379428 460856
rect 379480 460844 379486 460896
rect 50982 460776 50988 460828
rect 51040 460816 51046 460828
rect 78674 460816 78680 460828
rect 51040 460788 78680 460816
rect 51040 460776 51046 460788
rect 78674 460776 78680 460788
rect 78732 460776 78738 460828
rect 193858 460776 193864 460828
rect 193916 460816 193922 460828
rect 212994 460816 213000 460828
rect 193916 460788 213000 460816
rect 193916 460776 193922 460788
rect 212994 460776 213000 460788
rect 213052 460776 213058 460828
rect 266354 460776 266360 460828
rect 266412 460816 266418 460828
rect 358078 460816 358084 460828
rect 266412 460788 358084 460816
rect 266412 460776 266418 460788
rect 358078 460776 358084 460788
rect 358136 460776 358142 460828
rect 53466 460708 53472 460760
rect 53524 460748 53530 460760
rect 77294 460748 77300 460760
rect 53524 460720 77300 460748
rect 53524 460708 53530 460720
rect 77294 460708 77300 460720
rect 77352 460708 77358 460760
rect 189258 460708 189264 460760
rect 189316 460748 189322 460760
rect 210234 460748 210240 460760
rect 189316 460720 210240 460748
rect 189316 460708 189322 460720
rect 210234 460708 210240 460720
rect 210292 460708 210298 460760
rect 281534 460708 281540 460760
rect 281592 460748 281598 460760
rect 379330 460748 379336 460760
rect 281592 460720 379336 460748
rect 281592 460708 281598 460720
rect 379330 460708 379336 460720
rect 379388 460708 379394 460760
rect 52270 460640 52276 460692
rect 52328 460680 52334 460692
rect 75914 460680 75920 460692
rect 52328 460652 75920 460680
rect 52328 460640 52334 460652
rect 75914 460640 75920 460652
rect 75972 460640 75978 460692
rect 172606 460640 172612 460692
rect 172664 460680 172670 460692
rect 207750 460680 207756 460692
rect 172664 460652 207756 460680
rect 172664 460640 172670 460652
rect 207750 460640 207756 460652
rect 207808 460640 207814 460692
rect 258074 460640 258080 460692
rect 258132 460680 258138 460692
rect 364058 460680 364064 460692
rect 258132 460652 364064 460680
rect 258132 460640 258138 460652
rect 364058 460640 364064 460652
rect 364116 460640 364122 460692
rect 55490 460572 55496 460624
rect 55548 460612 55554 460624
rect 78766 460612 78772 460624
rect 55548 460584 78772 460612
rect 55548 460572 55554 460584
rect 78766 460572 78772 460584
rect 78824 460572 78830 460624
rect 179506 460572 179512 460624
rect 179564 460612 179570 460624
rect 214742 460612 214748 460624
rect 179564 460584 214748 460612
rect 179564 460572 179570 460584
rect 214742 460572 214748 460584
rect 214800 460572 214806 460624
rect 248414 460572 248420 460624
rect 248472 460612 248478 460624
rect 366634 460612 366640 460624
rect 248472 460584 366640 460612
rect 248472 460572 248478 460584
rect 366634 460572 366640 460584
rect 366692 460572 366698 460624
rect 55122 460504 55128 460556
rect 55180 460544 55186 460556
rect 71866 460544 71872 460556
rect 55180 460516 71872 460544
rect 55180 460504 55186 460516
rect 71866 460504 71872 460516
rect 71924 460504 71930 460556
rect 179414 460504 179420 460556
rect 179472 460544 179478 460556
rect 214834 460544 214840 460556
rect 179472 460516 214840 460544
rect 179472 460504 179478 460516
rect 214834 460504 214840 460516
rect 214892 460504 214898 460556
rect 249794 460504 249800 460556
rect 249852 460544 249858 460556
rect 368014 460544 368020 460556
rect 249852 460516 368020 460544
rect 249852 460504 249858 460516
rect 368014 460504 368020 460516
rect 368072 460504 368078 460556
rect 52362 460436 52368 460488
rect 52420 460476 52426 460488
rect 70394 460476 70400 460488
rect 52420 460448 70400 460476
rect 52420 460436 52426 460448
rect 70394 460436 70400 460448
rect 70452 460436 70458 460488
rect 162118 460436 162124 460488
rect 162176 460476 162182 460488
rect 197722 460476 197728 460488
rect 162176 460448 197728 460476
rect 162176 460436 162182 460448
rect 197722 460436 197728 460448
rect 197780 460436 197786 460488
rect 249978 460436 249984 460488
rect 250036 460476 250042 460488
rect 369210 460476 369216 460488
rect 250036 460448 369216 460476
rect 250036 460436 250042 460448
rect 369210 460436 369216 460448
rect 369268 460436 369274 460488
rect 43990 460368 43996 460420
rect 44048 460408 44054 460420
rect 67634 460408 67640 460420
rect 44048 460380 67640 460408
rect 44048 460368 44054 460380
rect 67634 460368 67640 460380
rect 67692 460368 67698 460420
rect 167086 460368 167092 460420
rect 167144 460408 167150 460420
rect 204990 460408 204996 460420
rect 167144 460380 204996 460408
rect 167144 460368 167150 460380
rect 204990 460368 204996 460380
rect 205048 460368 205054 460420
rect 242894 460368 242900 460420
rect 242952 460408 242958 460420
rect 365254 460408 365260 460420
rect 242952 460380 365260 460408
rect 242952 460368 242958 460380
rect 365254 460368 365260 460380
rect 365312 460368 365318 460420
rect 51902 460300 51908 460352
rect 51960 460340 51966 460352
rect 92566 460340 92572 460352
rect 51960 460312 92572 460340
rect 51960 460300 51966 460312
rect 92566 460300 92572 460312
rect 92624 460300 92630 460352
rect 168374 460300 168380 460352
rect 168432 460340 168438 460352
rect 206370 460340 206376 460352
rect 168432 460312 206376 460340
rect 168432 460300 168438 460312
rect 206370 460300 206376 460312
rect 206428 460300 206434 460352
rect 249886 460300 249892 460352
rect 249944 460340 249950 460352
rect 373350 460340 373356 460352
rect 249944 460312 373356 460340
rect 249944 460300 249950 460312
rect 373350 460300 373356 460312
rect 373408 460300 373414 460352
rect 45002 460232 45008 460284
rect 45060 460272 45066 460284
rect 103698 460272 103704 460284
rect 45060 460244 103704 460272
rect 45060 460232 45066 460244
rect 103698 460232 103704 460244
rect 103756 460232 103762 460284
rect 125594 460232 125600 460284
rect 125652 460272 125658 460284
rect 196894 460272 196900 460284
rect 125652 460244 196900 460272
rect 125652 460232 125658 460244
rect 196894 460232 196900 460244
rect 196952 460232 196958 460284
rect 248506 460232 248512 460284
rect 248564 460272 248570 460284
rect 372154 460272 372160 460284
rect 248564 460244 372160 460272
rect 248564 460232 248570 460244
rect 372154 460232 372160 460244
rect 372212 460232 372218 460284
rect 47670 460164 47676 460216
rect 47728 460204 47734 460216
rect 63494 460204 63500 460216
rect 47728 460176 63500 460204
rect 47728 460164 47734 460176
rect 63494 460164 63500 460176
rect 63552 460164 63558 460216
rect 63586 460164 63592 460216
rect 63644 460204 63650 460216
rect 199010 460204 199016 460216
rect 63644 460176 199016 460204
rect 63644 460164 63650 460176
rect 199010 460164 199016 460176
rect 199068 460164 199074 460216
rect 237374 460164 237380 460216
rect 237432 460204 237438 460216
rect 374730 460204 374736 460216
rect 237432 460176 374736 460204
rect 237432 460164 237438 460176
rect 374730 460164 374736 460176
rect 374788 460164 374794 460216
rect 50154 460096 50160 460148
rect 50212 460136 50218 460148
rect 66254 460136 66260 460148
rect 50212 460108 66260 460136
rect 50212 460096 50218 460108
rect 66254 460096 66260 460108
rect 66312 460096 66318 460148
rect 187694 460096 187700 460148
rect 187752 460136 187758 460148
rect 203794 460136 203800 460148
rect 187752 460108 203800 460136
rect 187752 460096 187758 460108
rect 203794 460096 203800 460108
rect 203852 460096 203858 460148
rect 280154 460096 280160 460148
rect 280212 460136 280218 460148
rect 357986 460136 357992 460148
rect 280212 460108 357992 460136
rect 280212 460096 280218 460108
rect 357986 460096 357992 460108
rect 358044 460096 358050 460148
rect 47762 460028 47768 460080
rect 47820 460068 47826 460080
rect 62114 460068 62120 460080
rect 47820 460040 62120 460068
rect 47820 460028 47826 460040
rect 62114 460028 62120 460040
rect 62172 460028 62178 460080
rect 193214 460028 193220 460080
rect 193272 460068 193278 460080
rect 208854 460068 208860 460080
rect 193272 460040 208860 460068
rect 193272 460028 193278 460040
rect 208854 460028 208860 460040
rect 208912 460028 208918 460080
rect 194686 459960 194692 460012
rect 194744 460000 194750 460012
rect 203518 460000 203524 460012
rect 194744 459972 203524 460000
rect 194744 459960 194750 459972
rect 203518 459960 203524 459972
rect 203576 459960 203582 460012
rect 214282 459620 214288 459672
rect 214340 459660 214346 459672
rect 220906 459660 220912 459672
rect 214340 459632 220912 459660
rect 214340 459620 214346 459632
rect 220906 459620 220912 459632
rect 220964 459620 220970 459672
rect 216306 459552 216312 459604
rect 216364 459592 216370 459604
rect 220814 459592 220820 459604
rect 216364 459564 220820 459592
rect 216364 459552 216370 459564
rect 220814 459552 220820 459564
rect 220872 459552 220878 459604
rect 191834 459484 191840 459536
rect 191892 459524 191898 459536
rect 208026 459524 208032 459536
rect 191892 459496 208032 459524
rect 191892 459484 191898 459496
rect 208026 459484 208032 459496
rect 208084 459484 208090 459536
rect 194594 459416 194600 459468
rect 194652 459456 194658 459468
rect 211522 459456 211528 459468
rect 194652 459428 211528 459456
rect 194652 459416 194658 459428
rect 211522 459416 211528 459428
rect 211580 459416 211586 459468
rect 291194 459416 291200 459468
rect 291252 459456 291258 459468
rect 360654 459456 360660 459468
rect 291252 459428 360660 459456
rect 291252 459416 291258 459428
rect 360654 459416 360660 459428
rect 360712 459416 360718 459468
rect 189166 459348 189172 459400
rect 189224 459388 189230 459400
rect 209498 459388 209504 459400
rect 189224 459360 209504 459388
rect 189224 459348 189230 459360
rect 209498 459348 209504 459360
rect 209556 459348 209562 459400
rect 282914 459348 282920 459400
rect 282972 459388 282978 459400
rect 359918 459388 359924 459400
rect 282972 459360 359924 459388
rect 282972 459348 282978 459360
rect 359918 459348 359924 459360
rect 359976 459348 359982 459400
rect 180794 459280 180800 459332
rect 180852 459320 180858 459332
rect 210786 459320 210792 459332
rect 180852 459292 210792 459320
rect 180852 459280 180858 459292
rect 210786 459280 210792 459292
rect 210844 459280 210850 459332
rect 288434 459280 288440 459332
rect 288492 459320 288498 459332
rect 374546 459320 374552 459332
rect 288492 459292 374552 459320
rect 288492 459280 288498 459292
rect 374546 459280 374552 459292
rect 374604 459280 374610 459332
rect 59170 459212 59176 459264
rect 59228 459252 59234 459264
rect 92474 459252 92480 459264
rect 59228 459224 92480 459252
rect 59228 459212 59234 459224
rect 92474 459212 92480 459224
rect 92532 459212 92538 459264
rect 173894 459212 173900 459264
rect 173952 459252 173958 459264
rect 206738 459252 206744 459264
rect 173952 459224 206744 459252
rect 173952 459212 173958 459224
rect 206738 459212 206744 459224
rect 206796 459212 206802 459264
rect 274634 459212 274640 459264
rect 274692 459252 274698 459264
rect 362862 459252 362868 459264
rect 274692 459224 362868 459252
rect 274692 459212 274698 459224
rect 362862 459212 362868 459224
rect 362920 459212 362926 459264
rect 51534 459144 51540 459196
rect 51592 459184 51598 459196
rect 99558 459184 99564 459196
rect 51592 459156 99564 459184
rect 51592 459144 51598 459156
rect 99558 459144 99564 459156
rect 99616 459144 99622 459196
rect 178034 459144 178040 459196
rect 178092 459184 178098 459196
rect 218974 459184 218980 459196
rect 178092 459156 218980 459184
rect 178092 459144 178098 459156
rect 218974 459144 218980 459156
rect 219032 459144 219038 459196
rect 270494 459144 270500 459196
rect 270552 459184 270558 459196
rect 363414 459184 363420 459196
rect 270552 459156 363420 459184
rect 270552 459144 270558 459156
rect 363414 459144 363420 459156
rect 363472 459144 363478 459196
rect 52730 459076 52736 459128
rect 52788 459116 52794 459128
rect 120074 459116 120080 459128
rect 52788 459088 120080 459116
rect 52788 459076 52794 459088
rect 120074 459076 120080 459088
rect 120132 459076 120138 459128
rect 142154 459076 142160 459128
rect 142212 459116 142218 459128
rect 197998 459116 198004 459128
rect 142212 459088 198004 459116
rect 142212 459076 142218 459088
rect 197998 459076 198004 459088
rect 198056 459076 198062 459128
rect 273254 459076 273260 459128
rect 273312 459116 273318 459128
rect 372982 459116 372988 459128
rect 273312 459088 372988 459116
rect 273312 459076 273318 459088
rect 372982 459076 372988 459088
rect 373040 459076 373046 459128
rect 54294 459008 54300 459060
rect 54352 459048 54358 459060
rect 131114 459048 131120 459060
rect 54352 459020 131120 459048
rect 54352 459008 54358 459020
rect 131114 459008 131120 459020
rect 131172 459008 131178 459060
rect 136634 459008 136640 459060
rect 136692 459048 136698 459060
rect 199286 459048 199292 459060
rect 136692 459020 199292 459048
rect 136692 459008 136698 459020
rect 199286 459008 199292 459020
rect 199344 459008 199350 459060
rect 264974 459008 264980 459060
rect 265032 459048 265038 459060
rect 369486 459048 369492 459060
rect 265032 459020 369492 459048
rect 265032 459008 265038 459020
rect 369486 459008 369492 459020
rect 369544 459008 369550 459060
rect 56226 458940 56232 458992
rect 56284 458980 56290 458992
rect 133966 458980 133972 458992
rect 56284 458952 133972 458980
rect 56284 458940 56290 458952
rect 133966 458940 133972 458952
rect 134024 458940 134030 458992
rect 135254 458940 135260 458992
rect 135312 458980 135318 458992
rect 197906 458980 197912 458992
rect 135312 458952 197912 458980
rect 135312 458940 135318 458952
rect 197906 458940 197912 458952
rect 197964 458940 197970 458992
rect 253934 458940 253940 458992
rect 253992 458980 253998 458992
rect 370958 458980 370964 458992
rect 253992 458952 370964 458980
rect 253992 458940 253998 458952
rect 370958 458940 370964 458952
rect 371016 458940 371022 458992
rect 52270 458872 52276 458924
rect 52328 458912 52334 458924
rect 133874 458912 133880 458924
rect 52328 458884 133880 458912
rect 52328 458872 52334 458884
rect 133874 458872 133880 458884
rect 133932 458872 133938 458924
rect 138014 458872 138020 458924
rect 138072 458912 138078 458924
rect 201862 458912 201868 458924
rect 138072 458884 201868 458912
rect 138072 458872 138078 458884
rect 201862 458872 201868 458884
rect 201920 458872 201926 458924
rect 247034 458872 247040 458924
rect 247092 458912 247098 458924
rect 367922 458912 367928 458924
rect 247092 458884 367928 458912
rect 247092 458872 247098 458884
rect 367922 458872 367928 458884
rect 367980 458872 367986 458924
rect 60734 458804 60740 458856
rect 60792 458844 60798 458856
rect 199562 458844 199568 458856
rect 60792 458816 199568 458844
rect 60792 458804 60798 458816
rect 199562 458804 199568 458816
rect 199620 458804 199626 458856
rect 245654 458804 245660 458856
rect 245712 458844 245718 458856
rect 379146 458844 379152 458856
rect 245712 458816 379152 458844
rect 245712 458804 245718 458816
rect 379146 458804 379152 458816
rect 379204 458804 379210 458856
rect 189074 458736 189080 458788
rect 189132 458776 189138 458788
rect 201034 458776 201040 458788
rect 189132 458748 201040 458776
rect 189132 458736 189138 458748
rect 201034 458736 201040 458748
rect 201092 458736 201098 458788
rect 199010 458328 199016 458380
rect 199068 458368 199074 458380
rect 199068 458340 354674 458368
rect 199068 458328 199074 458340
rect 47486 458260 47492 458312
rect 47544 458300 47550 458312
rect 354646 458300 354674 458340
rect 358814 458300 358820 458312
rect 47544 458272 200114 458300
rect 354646 458272 358820 458300
rect 47544 458260 47550 458272
rect 200086 458232 200114 458272
rect 358814 458260 358820 458272
rect 358872 458300 358878 458312
rect 516594 458300 516600 458312
rect 358872 458272 516600 458300
rect 358872 458260 358878 458272
rect 516594 458260 516600 458272
rect 516652 458260 516658 458312
rect 207382 458232 207388 458244
rect 200086 458204 207388 458232
rect 207382 458192 207388 458204
rect 207440 458232 207446 458244
rect 208118 458232 208124 458244
rect 207440 458204 208124 458232
rect 207440 458192 207446 458204
rect 208118 458192 208124 458204
rect 208176 458192 208182 458244
rect 53006 457784 53012 457836
rect 53064 457824 53070 457836
rect 53466 457824 53472 457836
rect 53064 457796 53472 457824
rect 53064 457784 53070 457796
rect 53466 457784 53472 457796
rect 53524 457784 53530 457836
rect 49234 456084 49240 456136
rect 49292 456124 49298 456136
rect 49602 456124 49608 456136
rect 49292 456096 49608 456124
rect 49292 456084 49298 456096
rect 49602 456084 49608 456096
rect 49660 456084 49666 456136
rect 518158 441532 518164 441584
rect 518216 441572 518222 441584
rect 579890 441572 579896 441584
rect 518216 441544 579896 441572
rect 518216 441532 518222 441544
rect 579890 441532 579896 441544
rect 579948 441532 579954 441584
rect 3142 422220 3148 422272
rect 3200 422260 3206 422272
rect 18598 422260 18604 422272
rect 3200 422232 18604 422260
rect 3200 422220 3206 422232
rect 18598 422220 18604 422232
rect 18656 422220 18662 422272
rect 54478 416644 54484 416696
rect 54536 416684 54542 416696
rect 57238 416684 57244 416696
rect 54536 416656 57244 416684
rect 54536 416644 54542 416656
rect 57238 416644 57244 416656
rect 57296 416644 57302 416696
rect 56226 415352 56232 415404
rect 56284 415392 56290 415404
rect 56594 415392 56600 415404
rect 56284 415364 56600 415392
rect 56284 415352 56290 415364
rect 56594 415352 56600 415364
rect 56652 415352 56658 415404
rect 47578 412564 47584 412616
rect 47636 412604 47642 412616
rect 57238 412604 57244 412616
rect 47636 412576 57244 412604
rect 47636 412564 47642 412576
rect 57238 412564 57244 412576
rect 57296 412564 57302 412616
rect 47486 411204 47492 411256
rect 47544 411244 47550 411256
rect 57238 411244 57244 411256
rect 47544 411216 57244 411244
rect 47544 411204 47550 411216
rect 57238 411204 57244 411216
rect 57296 411204 57302 411256
rect 50798 411068 50804 411120
rect 50856 411108 50862 411120
rect 55674 411108 55680 411120
rect 50856 411080 55680 411108
rect 50856 411068 50862 411080
rect 55674 411068 55680 411080
rect 55732 411068 55738 411120
rect 208118 410524 208124 410576
rect 208176 410564 208182 410576
rect 216766 410564 216772 410576
rect 208176 410536 216772 410564
rect 208176 410524 208182 410536
rect 216766 410524 216772 410536
rect 216824 410524 216830 410576
rect 205726 409096 205732 409148
rect 205784 409136 205790 409148
rect 216766 409136 216772 409148
rect 205784 409108 216772 409136
rect 205784 409096 205790 409108
rect 216766 409096 216772 409108
rect 216824 409096 216830 409148
rect 56226 408552 56232 408604
rect 56284 408592 56290 408604
rect 56594 408592 56600 408604
rect 56284 408564 56600 408592
rect 56284 408552 56290 408564
rect 56594 408552 56600 408564
rect 56652 408552 56658 408604
rect 57054 408552 57060 408604
rect 57112 408592 57118 408604
rect 57974 408592 57980 408604
rect 57112 408564 57980 408592
rect 57112 408552 57118 408564
rect 57974 408552 57980 408564
rect 58032 408552 58038 408604
rect 47578 408484 47584 408536
rect 47636 408524 47642 408536
rect 57238 408524 57244 408536
rect 47636 408496 57244 408524
rect 47636 408484 47642 408496
rect 57238 408484 57244 408496
rect 57296 408484 57302 408536
rect 58526 407736 58532 407788
rect 58584 407776 58590 407788
rect 59354 407776 59360 407788
rect 58584 407748 59360 407776
rect 58584 407736 58590 407748
rect 59354 407736 59360 407748
rect 59412 407736 59418 407788
rect 57054 407464 57060 407516
rect 57112 407504 57118 407516
rect 59630 407504 59636 407516
rect 57112 407476 59636 407504
rect 57112 407464 57118 407476
rect 59630 407464 59636 407476
rect 59688 407464 59694 407516
rect 47486 407124 47492 407176
rect 47544 407164 47550 407176
rect 57238 407164 57244 407176
rect 47544 407136 57244 407164
rect 47544 407124 47550 407136
rect 57238 407124 57244 407136
rect 57296 407124 57302 407176
rect 360838 406376 360844 406428
rect 360896 406416 360902 406428
rect 377398 406416 377404 406428
rect 360896 406388 377404 406416
rect 360896 406376 360902 406388
rect 377398 406376 377404 406388
rect 377456 406376 377462 406428
rect 47394 405696 47400 405748
rect 47452 405736 47458 405748
rect 57238 405736 57244 405748
rect 47452 405708 57244 405736
rect 47452 405696 47458 405708
rect 57238 405696 57244 405708
rect 57296 405696 57302 405748
rect 204438 404948 204444 405000
rect 204496 404988 204502 405000
rect 216858 404988 216864 405000
rect 204496 404960 216864 404988
rect 204496 404948 204502 404960
rect 216858 404948 216864 404960
rect 216916 404948 216922 405000
rect 359918 404948 359924 405000
rect 359976 404988 359982 405000
rect 377674 404988 377680 405000
rect 359976 404960 377680 404988
rect 359976 404948 359982 404960
rect 377674 404948 377680 404960
rect 377732 404948 377738 405000
rect 50798 404336 50804 404388
rect 50856 404376 50862 404388
rect 57238 404376 57244 404388
rect 50856 404348 57244 404376
rect 50856 404336 50862 404348
rect 57238 404336 57244 404348
rect 57296 404336 57302 404388
rect 359826 403588 359832 403640
rect 359884 403628 359890 403640
rect 377766 403628 377772 403640
rect 359884 403600 377772 403628
rect 359884 403588 359890 403600
rect 377766 403588 377772 403600
rect 377824 403588 377830 403640
rect 50982 402976 50988 403028
rect 51040 403016 51046 403028
rect 57238 403016 57244 403028
rect 51040 402988 57244 403016
rect 51040 402976 51046 402988
rect 57238 402976 57244 402988
rect 57296 402976 57302 403028
rect 360102 389308 360108 389360
rect 360160 389348 360166 389360
rect 361666 389348 361672 389360
rect 360160 389320 361672 389348
rect 360160 389308 360166 389320
rect 361666 389308 361672 389320
rect 361724 389308 361730 389360
rect 46014 384956 46020 385008
rect 46072 384996 46078 385008
rect 57238 384996 57244 385008
rect 46072 384968 57244 384996
rect 46072 384956 46078 384968
rect 57238 384956 57244 384968
rect 57296 384956 57302 385008
rect 206278 384956 206284 385008
rect 206336 384996 206342 385008
rect 216674 384996 216680 385008
rect 206336 384968 216680 384996
rect 206336 384956 206342 384968
rect 216674 384956 216680 384968
rect 216732 384956 216738 385008
rect 359550 384956 359556 385008
rect 359608 384996 359614 385008
rect 376938 384996 376944 385008
rect 359608 384968 376944 384996
rect 359608 384956 359614 384968
rect 376938 384956 376944 384968
rect 376996 384956 377002 385008
rect 47946 383596 47952 383648
rect 48004 383636 48010 383648
rect 56870 383636 56876 383648
rect 48004 383608 56876 383636
rect 48004 383596 48010 383608
rect 56870 383596 56876 383608
rect 56928 383596 56934 383648
rect 207014 383596 207020 383648
rect 207072 383636 207078 383648
rect 216674 383636 216680 383648
rect 207072 383608 216680 383636
rect 207072 383596 207078 383608
rect 216674 383596 216680 383608
rect 216732 383596 216738 383648
rect 361574 383596 361580 383648
rect 361632 383636 361638 383648
rect 376938 383636 376944 383648
rect 361632 383608 376944 383636
rect 361632 383596 361638 383608
rect 376938 383596 376944 383608
rect 376996 383596 377002 383648
rect 57146 383528 57152 383580
rect 57204 383568 57210 383580
rect 57606 383568 57612 383580
rect 57204 383540 57612 383568
rect 57204 383528 57210 383540
rect 57606 383528 57612 383540
rect 57664 383528 57670 383580
rect 209498 383528 209504 383580
rect 209556 383568 209562 383580
rect 217042 383568 217048 383580
rect 209556 383540 217048 383568
rect 209556 383528 209562 383540
rect 217042 383528 217048 383540
rect 217100 383528 217106 383580
rect 359458 383528 359464 383580
rect 359516 383568 359522 383580
rect 376846 383568 376852 383580
rect 359516 383540 376852 383568
rect 359516 383528 359522 383540
rect 376846 383528 376852 383540
rect 376904 383528 376910 383580
rect 56962 382304 56968 382356
rect 57020 382344 57026 382356
rect 57238 382344 57244 382356
rect 57020 382316 57244 382344
rect 57020 382304 57026 382316
rect 57238 382304 57244 382316
rect 57296 382304 57302 382356
rect 206278 382236 206284 382288
rect 206336 382276 206342 382288
rect 207014 382276 207020 382288
rect 206336 382248 207020 382276
rect 206336 382236 206342 382248
rect 207014 382236 207020 382248
rect 207072 382236 207078 382288
rect 360838 382236 360844 382288
rect 360896 382276 360902 382288
rect 361574 382276 361580 382288
rect 360896 382248 361580 382276
rect 360896 382236 360902 382248
rect 361574 382236 361580 382248
rect 361632 382236 361638 382288
rect 42702 382168 42708 382220
rect 42760 382208 42766 382220
rect 57238 382208 57244 382220
rect 42760 382180 57244 382208
rect 42760 382168 42766 382180
rect 57238 382168 57244 382180
rect 57296 382208 57302 382220
rect 57514 382208 57520 382220
rect 57296 382180 57520 382208
rect 57296 382168 57302 382180
rect 57514 382168 57520 382180
rect 57572 382168 57578 382220
rect 47946 380876 47952 380928
rect 48004 380916 48010 380928
rect 48774 380916 48780 380928
rect 48004 380888 48780 380916
rect 48004 380876 48010 380888
rect 48774 380876 48780 380888
rect 48832 380876 48838 380928
rect 212902 380672 212908 380724
rect 212960 380672 212966 380724
rect 212920 380520 212948 380672
rect 212902 380468 212908 380520
rect 212960 380468 212966 380520
rect 57146 377748 57152 377800
rect 57204 377788 57210 377800
rect 57606 377788 57612 377800
rect 57204 377760 57612 377788
rect 57204 377748 57210 377760
rect 57606 377748 57612 377760
rect 57664 377748 57670 377800
rect 216766 375300 216772 375352
rect 216824 375340 216830 375352
rect 217778 375340 217784 375352
rect 216824 375312 217784 375340
rect 216824 375300 216830 375312
rect 217778 375300 217784 375312
rect 217836 375300 217842 375352
rect 47578 375028 47584 375080
rect 47636 375068 47642 375080
rect 216766 375068 216772 375080
rect 47636 375040 216772 375068
rect 47636 375028 47642 375040
rect 216766 375028 216772 375040
rect 216824 375028 216830 375080
rect 47486 374960 47492 375012
rect 47544 375000 47550 375012
rect 217226 375000 217232 375012
rect 47544 374972 217232 375000
rect 47544 374960 47550 374972
rect 217226 374960 217232 374972
rect 217284 374960 217290 375012
rect 58802 374892 58808 374944
rect 58860 374932 58866 374944
rect 60734 374932 60740 374944
rect 58860 374904 60740 374932
rect 58860 374892 58866 374904
rect 60734 374892 60740 374904
rect 60792 374892 60798 374944
rect 58894 374824 58900 374876
rect 58952 374864 58958 374876
rect 62114 374864 62120 374876
rect 58952 374836 62120 374864
rect 58952 374824 58958 374836
rect 62114 374824 62120 374836
rect 62172 374824 62178 374876
rect 208946 374824 208952 374876
rect 209004 374864 209010 374876
rect 218238 374864 218244 374876
rect 209004 374836 218244 374864
rect 209004 374824 209010 374836
rect 218238 374824 218244 374836
rect 218296 374824 218302 374876
rect 140958 374756 140964 374808
rect 141016 374796 141022 374808
rect 201862 374796 201868 374808
rect 141016 374768 201868 374796
rect 141016 374756 141022 374768
rect 201862 374756 201868 374768
rect 201920 374756 201926 374808
rect 203058 374756 203064 374808
rect 203116 374796 203122 374808
rect 281442 374796 281448 374808
rect 203116 374768 281448 374796
rect 203116 374756 203122 374768
rect 281442 374756 281448 374768
rect 281500 374756 281506 374808
rect 359734 374756 359740 374808
rect 359792 374796 359798 374808
rect 440326 374796 440332 374808
rect 359792 374768 440332 374796
rect 359792 374756 359798 374768
rect 440326 374756 440332 374768
rect 440384 374756 440390 374808
rect 201494 374688 201500 374740
rect 201552 374728 201558 374740
rect 311802 374728 311808 374740
rect 201552 374700 311808 374728
rect 201552 374688 201558 374700
rect 311802 374688 311808 374700
rect 311860 374688 311866 374740
rect 358630 374688 358636 374740
rect 358688 374728 358694 374740
rect 372890 374728 372896 374740
rect 358688 374700 372896 374728
rect 358688 374688 358694 374700
rect 372890 374688 372896 374700
rect 372948 374688 372954 374740
rect 201678 374620 201684 374672
rect 201736 374660 201742 374672
rect 314562 374660 314568 374672
rect 201736 374632 314568 374660
rect 201736 374620 201742 374632
rect 314562 374620 314568 374632
rect 314620 374620 314626 374672
rect 372430 374620 372436 374672
rect 372488 374660 372494 374672
rect 418246 374660 418252 374672
rect 372488 374632 418252 374660
rect 372488 374620 372494 374632
rect 418246 374620 418252 374632
rect 418304 374620 418310 374672
rect 165982 374552 165988 374604
rect 166040 374592 166046 374604
rect 199102 374592 199108 374604
rect 166040 374564 199108 374592
rect 166040 374552 166046 374564
rect 199102 374552 199108 374564
rect 199160 374552 199166 374604
rect 360746 374552 360752 374604
rect 360804 374592 360810 374604
rect 407758 374592 407764 374604
rect 360804 374564 407764 374592
rect 360804 374552 360810 374564
rect 407758 374552 407764 374564
rect 407816 374552 407822 374604
rect 163406 374484 163412 374536
rect 163464 374524 163470 374536
rect 197998 374524 198004 374536
rect 163464 374496 198004 374524
rect 163464 374484 163470 374496
rect 197998 374484 198004 374496
rect 198056 374484 198062 374536
rect 361482 374484 361488 374536
rect 361540 374524 361546 374536
rect 410702 374524 410708 374536
rect 361540 374496 410708 374524
rect 361540 374484 361546 374496
rect 410702 374484 410708 374496
rect 410760 374484 410766 374536
rect 158530 374416 158536 374468
rect 158588 374456 158594 374468
rect 201770 374456 201776 374468
rect 158588 374428 201776 374456
rect 158588 374416 158594 374428
rect 201770 374416 201776 374428
rect 201828 374416 201834 374468
rect 213546 374416 213552 374468
rect 213604 374456 213610 374468
rect 244274 374456 244280 374468
rect 213604 374428 244280 374456
rect 213604 374416 213610 374428
rect 244274 374416 244280 374428
rect 244332 374416 244338 374468
rect 372890 374416 372896 374468
rect 372948 374456 372954 374468
rect 373810 374456 373816 374468
rect 372948 374428 373816 374456
rect 372948 374416 372954 374428
rect 373810 374416 373816 374428
rect 373868 374456 373874 374468
rect 433334 374456 433340 374468
rect 373868 374428 433340 374456
rect 373868 374416 373874 374428
rect 433334 374416 433340 374428
rect 433392 374416 433398 374468
rect 160922 374348 160928 374400
rect 160980 374388 160986 374400
rect 207474 374388 207480 374400
rect 160980 374360 207480 374388
rect 160980 374348 160986 374360
rect 207474 374348 207480 374360
rect 207532 374348 207538 374400
rect 241238 374348 241244 374400
rect 241296 374388 241302 374400
rect 248690 374388 248696 374400
rect 241296 374360 248696 374388
rect 241296 374348 241302 374360
rect 248690 374348 248696 374360
rect 248748 374348 248754 374400
rect 377490 374348 377496 374400
rect 377548 374388 377554 374400
rect 443086 374388 443092 374400
rect 377548 374360 443092 374388
rect 377548 374348 377554 374360
rect 443086 374348 443092 374360
rect 443144 374348 443150 374400
rect 153470 374280 153476 374332
rect 153528 374320 153534 374332
rect 200482 374320 200488 374332
rect 153528 374292 200488 374320
rect 153528 374280 153534 374292
rect 200482 374280 200488 374292
rect 200540 374280 200546 374332
rect 241146 374280 241152 374332
rect 241204 374320 241210 374332
rect 250070 374320 250076 374332
rect 241204 374292 250076 374320
rect 241204 374280 241210 374292
rect 250070 374280 250076 374292
rect 250128 374280 250134 374332
rect 367002 374280 367008 374332
rect 367060 374320 367066 374332
rect 434806 374320 434812 374332
rect 367060 374292 434812 374320
rect 367060 374280 367066 374292
rect 434806 374280 434812 374292
rect 434864 374280 434870 374332
rect 148962 374212 148968 374264
rect 149020 374252 149026 374264
rect 197078 374252 197084 374264
rect 149020 374224 197084 374252
rect 149020 374212 149026 374224
rect 197078 374212 197084 374224
rect 197136 374212 197142 374264
rect 215478 374212 215484 374264
rect 215536 374252 215542 374264
rect 263686 374252 263692 374264
rect 215536 374224 263692 374252
rect 215536 374212 215542 374224
rect 263686 374212 263692 374224
rect 263744 374212 263750 374264
rect 363506 374212 363512 374264
rect 363564 374252 363570 374264
rect 433610 374252 433616 374264
rect 363564 374224 433616 374252
rect 363564 374212 363570 374224
rect 433610 374212 433616 374224
rect 433668 374212 433674 374264
rect 146202 374144 146208 374196
rect 146260 374184 146266 374196
rect 204530 374184 204536 374196
rect 146260 374156 204536 374184
rect 146260 374144 146266 374156
rect 204530 374144 204536 374156
rect 204588 374144 204594 374196
rect 218238 374144 218244 374196
rect 218296 374184 218302 374196
rect 271138 374184 271144 374196
rect 218296 374156 271144 374184
rect 218296 374144 218302 374156
rect 271138 374144 271144 374156
rect 271196 374144 271202 374196
rect 372982 374144 372988 374196
rect 373040 374184 373046 374196
rect 445938 374184 445944 374196
rect 373040 374156 445944 374184
rect 373040 374144 373046 374156
rect 445938 374144 445944 374156
rect 445996 374144 446002 374196
rect 143534 374076 143540 374128
rect 143592 374116 143598 374128
rect 213086 374116 213092 374128
rect 143592 374088 213092 374116
rect 143592 374076 143598 374088
rect 213086 374076 213092 374088
rect 213144 374076 213150 374128
rect 219618 374076 219624 374128
rect 219676 374116 219682 374128
rect 222010 374116 222016 374128
rect 219676 374088 222016 374116
rect 219676 374076 219682 374088
rect 222010 374076 222016 374088
rect 222068 374076 222074 374128
rect 270310 374076 270316 374128
rect 270368 374116 270374 374128
rect 275830 374116 275836 374128
rect 270368 374088 275836 374116
rect 270368 374076 270374 374088
rect 275830 374076 275836 374088
rect 275888 374076 275894 374128
rect 371050 374076 371056 374128
rect 371108 374116 371114 374128
rect 448238 374116 448244 374128
rect 371108 374088 448244 374116
rect 371108 374076 371114 374088
rect 448238 374076 448244 374088
rect 448296 374076 448302 374128
rect 56962 374008 56968 374060
rect 57020 374048 57026 374060
rect 105446 374048 105452 374060
rect 57020 374020 105452 374048
rect 57020 374008 57026 374020
rect 105446 374008 105452 374020
rect 105504 374008 105510 374060
rect 201586 374008 201592 374060
rect 201644 374048 201650 374060
rect 320910 374048 320916 374060
rect 201644 374020 320916 374048
rect 201644 374008 201650 374020
rect 320910 374008 320916 374020
rect 320968 374008 320974 374060
rect 373902 374008 373908 374060
rect 373960 374048 373966 374060
rect 373960 374020 375328 374048
rect 373960 374008 373966 374020
rect 47394 373940 47400 373992
rect 47452 373980 47458 373992
rect 217594 373980 217600 373992
rect 47452 373952 217600 373980
rect 47452 373940 47458 373952
rect 217594 373940 217600 373952
rect 217652 373940 217658 373992
rect 375300 373980 375328 374020
rect 404814 373980 404820 373992
rect 375300 373952 404820 373980
rect 404814 373940 404820 373952
rect 404872 373940 404878 373992
rect 58710 373872 58716 373924
rect 58768 373912 58774 373924
rect 116118 373912 116124 373924
rect 58768 373884 116124 373912
rect 58768 373872 58774 373884
rect 116118 373872 116124 373884
rect 116176 373872 116182 373924
rect 139210 373872 139216 373924
rect 139268 373912 139274 373924
rect 200298 373912 200304 373924
rect 139268 373884 200304 373912
rect 139268 373872 139274 373884
rect 200298 373872 200304 373884
rect 200356 373872 200362 373924
rect 369670 373872 369676 373924
rect 369728 373912 369734 373924
rect 421006 373912 421012 373924
rect 369728 373884 421012 373912
rect 369728 373872 369734 373884
rect 421006 373872 421012 373884
rect 421064 373872 421070 373924
rect 43346 373804 43352 373856
rect 43404 373844 43410 373856
rect 103514 373844 103520 373856
rect 43404 373816 103520 373844
rect 43404 373804 43410 373816
rect 103514 373804 103520 373816
rect 103572 373804 103578 373856
rect 136450 373804 136456 373856
rect 136508 373844 136514 373856
rect 200390 373844 200396 373856
rect 136508 373816 200396 373844
rect 136508 373804 136514 373816
rect 200390 373804 200396 373816
rect 200448 373804 200454 373856
rect 366174 373804 366180 373856
rect 366232 373844 366238 373856
rect 423030 373844 423036 373856
rect 366232 373816 423036 373844
rect 366232 373804 366238 373816
rect 423030 373804 423036 373816
rect 423088 373804 423094 373856
rect 52270 373736 52276 373788
rect 52328 373776 52334 373788
rect 113542 373776 113548 373788
rect 52328 373748 113548 373776
rect 52328 373736 52334 373748
rect 113542 373736 113548 373748
rect 113600 373736 113606 373788
rect 131022 373736 131028 373788
rect 131080 373776 131086 373788
rect 199286 373776 199292 373788
rect 131080 373748 199292 373776
rect 131080 373736 131086 373748
rect 199286 373736 199292 373748
rect 199344 373736 199350 373788
rect 219434 373736 219440 373788
rect 219492 373776 219498 373788
rect 219618 373776 219624 373788
rect 219492 373748 219624 373776
rect 219492 373736 219498 373748
rect 219618 373736 219624 373748
rect 219676 373736 219682 373788
rect 368382 373736 368388 373788
rect 368440 373776 368446 373788
rect 376846 373776 376852 373788
rect 368440 373748 376852 373776
rect 368440 373736 368446 373748
rect 376846 373736 376852 373748
rect 376904 373736 376910 373788
rect 379422 373736 379428 373788
rect 379480 373776 379486 373788
rect 439406 373776 439412 373788
rect 379480 373748 439412 373776
rect 379480 373736 379486 373748
rect 439406 373736 439412 373748
rect 439464 373736 439470 373788
rect 56226 373668 56232 373720
rect 56284 373708 56290 373720
rect 118326 373708 118332 373720
rect 56284 373680 118332 373708
rect 56284 373668 56290 373680
rect 118326 373668 118332 373680
rect 118384 373668 118390 373720
rect 128906 373668 128912 373720
rect 128964 373708 128970 373720
rect 198918 373708 198924 373720
rect 128964 373680 198924 373708
rect 128964 373668 128970 373680
rect 198918 373668 198924 373680
rect 198976 373668 198982 373720
rect 215294 373668 215300 373720
rect 215352 373708 215358 373720
rect 215570 373708 215576 373720
rect 215352 373680 215576 373708
rect 215352 373668 215358 373680
rect 215570 373668 215576 373680
rect 215628 373708 215634 373720
rect 219250 373708 219256 373720
rect 215628 373680 219256 373708
rect 215628 373668 215634 373680
rect 219250 373668 219256 373680
rect 219308 373668 219314 373720
rect 363414 373668 363420 373720
rect 363472 373708 363478 373720
rect 425422 373708 425428 373720
rect 363472 373680 425428 373708
rect 363472 373668 363478 373680
rect 425422 373668 425428 373680
rect 425480 373668 425486 373720
rect 57054 373600 57060 373652
rect 57112 373640 57118 373652
rect 125686 373640 125692 373652
rect 57112 373612 125692 373640
rect 57112 373600 57118 373612
rect 125686 373600 125692 373612
rect 125744 373600 125750 373652
rect 133690 373600 133696 373652
rect 133748 373640 133754 373652
rect 205818 373640 205824 373652
rect 133748 373612 205824 373640
rect 133748 373600 133754 373612
rect 205818 373600 205824 373612
rect 205876 373600 205882 373652
rect 367646 373600 367652 373652
rect 367704 373640 367710 373652
rect 450262 373640 450268 373652
rect 367704 373612 450268 373640
rect 367704 373600 367710 373612
rect 450262 373600 450268 373612
rect 450320 373600 450326 373652
rect 48866 373532 48872 373584
rect 48924 373572 48930 373584
rect 110414 373572 110420 373584
rect 48924 373544 110420 373572
rect 48924 373532 48930 373544
rect 110414 373532 110420 373544
rect 110472 373532 110478 373584
rect 121362 373532 121368 373584
rect 121420 373572 121426 373584
rect 197906 373572 197912 373584
rect 121420 373544 197912 373572
rect 121420 373532 121426 373544
rect 197906 373532 197912 373544
rect 197964 373532 197970 373584
rect 215294 373532 215300 373584
rect 215352 373572 215358 373584
rect 216490 373572 216496 373584
rect 215352 373544 216496 373572
rect 215352 373532 215358 373544
rect 216490 373532 216496 373544
rect 216548 373572 216554 373584
rect 236454 373572 236460 373584
rect 216548 373544 236460 373572
rect 216548 373532 216554 373544
rect 236454 373532 236460 373544
rect 236512 373532 236518 373584
rect 375098 373532 375104 373584
rect 375156 373572 375162 373584
rect 460934 373572 460940 373584
rect 375156 373544 460940 373572
rect 375156 373532 375162 373544
rect 460934 373532 460940 373544
rect 460992 373532 460998 373584
rect 46106 373464 46112 373516
rect 46164 373504 46170 373516
rect 107838 373504 107844 373516
rect 46164 373476 107844 373504
rect 46164 373464 46170 373476
rect 107838 373464 107844 373476
rect 107896 373464 107902 373516
rect 124122 373464 124128 373516
rect 124180 373504 124186 373516
rect 203242 373504 203248 373516
rect 124180 373476 203248 373504
rect 124180 373464 124186 373476
rect 203242 373464 203248 373476
rect 203300 373464 203306 373516
rect 209774 373464 209780 373516
rect 209832 373504 209838 373516
rect 211062 373504 211068 373516
rect 209832 373476 211068 373504
rect 209832 373464 209838 373476
rect 211062 373464 211068 373476
rect 211120 373504 211126 373516
rect 214926 373504 214932 373516
rect 211120 373476 214932 373504
rect 211120 373464 211126 373476
rect 214926 373464 214932 373476
rect 214984 373504 214990 373516
rect 224218 373504 224224 373516
rect 214984 373476 224224 373504
rect 214984 373464 214990 373476
rect 224218 373464 224224 373476
rect 224276 373464 224282 373516
rect 364794 373464 364800 373516
rect 364852 373504 364858 373516
rect 452838 373504 452844 373516
rect 364852 373476 452844 373504
rect 364852 373464 364858 373476
rect 452838 373464 452844 373476
rect 452896 373464 452902 373516
rect 55674 373396 55680 373448
rect 55732 373436 55738 373448
rect 98270 373436 98276 373448
rect 55732 373408 98276 373436
rect 55732 373396 55738 373408
rect 98270 373396 98276 373408
rect 98328 373396 98334 373448
rect 98362 373396 98368 373448
rect 98420 373436 98426 373448
rect 212718 373436 212724 373448
rect 98420 373408 212724 373436
rect 98420 373396 98426 373408
rect 212718 373396 212724 373408
rect 212776 373396 212782 373448
rect 215018 373396 215024 373448
rect 215076 373436 215082 373448
rect 242894 373436 242900 373448
rect 215076 373408 242900 373436
rect 215076 373396 215082 373408
rect 242894 373396 242900 373408
rect 242952 373396 242958 373448
rect 371694 373396 371700 373448
rect 371752 373436 371758 373448
rect 462774 373436 462780 373448
rect 371752 373408 462780 373436
rect 371752 373396 371758 373408
rect 462774 373396 462780 373408
rect 462832 373396 462838 373448
rect 48682 373328 48688 373380
rect 48740 373368 48746 373380
rect 96062 373368 96068 373380
rect 48740 373340 96068 373368
rect 48740 373328 48746 373340
rect 96062 373328 96068 373340
rect 96120 373328 96126 373380
rect 96154 373328 96160 373380
rect 96212 373368 96218 373380
rect 212626 373368 212632 373380
rect 96212 373340 212632 373368
rect 96212 373328 96218 373340
rect 212626 373328 212632 373340
rect 212684 373328 212690 373380
rect 215266 373340 219204 373368
rect 47854 373260 47860 373312
rect 47912 373300 47918 373312
rect 90174 373300 90180 373312
rect 47912 373272 90180 373300
rect 47912 373260 47918 373272
rect 90174 373260 90180 373272
rect 90232 373260 90238 373312
rect 95050 373260 95056 373312
rect 95108 373300 95114 373312
rect 212534 373300 212540 373312
rect 95108 373272 212540 373300
rect 95108 373260 95114 373272
rect 212534 373260 212540 373272
rect 212592 373300 212598 373312
rect 215266 373300 215294 373340
rect 212592 373272 215294 373300
rect 212592 373260 212598 373272
rect 219176 373244 219204 373340
rect 362862 373328 362868 373380
rect 362920 373368 362926 373380
rect 455414 373368 455420 373380
rect 362920 373340 455420 373368
rect 362920 373328 362926 373340
rect 455414 373328 455420 373340
rect 455472 373328 455478 373380
rect 219342 373260 219348 373312
rect 219400 373300 219406 373312
rect 269206 373300 269212 373312
rect 219400 373272 269212 373300
rect 219400 373260 219406 373272
rect 269206 373260 269212 373272
rect 269264 373260 269270 373312
rect 364242 373260 364248 373312
rect 364300 373300 364306 373312
rect 458174 373300 458180 373312
rect 364300 373272 458180 373300
rect 364300 373260 364306 373272
rect 458174 373260 458180 373272
rect 458232 373260 458238 373312
rect 54294 373192 54300 373244
rect 54352 373232 54358 373244
rect 100846 373232 100852 373244
rect 54352 373204 100852 373232
rect 54352 373192 54358 373204
rect 100846 373192 100852 373204
rect 100904 373192 100910 373244
rect 151722 373192 151728 373244
rect 151780 373232 151786 373244
rect 197814 373232 197820 373244
rect 151780 373204 197820 373232
rect 151780 373192 151786 373204
rect 197814 373192 197820 373204
rect 197872 373192 197878 373244
rect 219158 373192 219164 373244
rect 219216 373232 219222 373244
rect 253934 373232 253940 373244
rect 219216 373204 253940 373232
rect 219216 373192 219222 373204
rect 253934 373192 253940 373204
rect 253992 373192 253998 373244
rect 365622 373192 365628 373244
rect 365680 373232 365686 373244
rect 380894 373232 380900 373244
rect 365680 373204 380900 373232
rect 365680 373192 365686 373204
rect 380894 373192 380900 373204
rect 380952 373192 380958 373244
rect 54386 373124 54392 373176
rect 54444 373164 54450 373176
rect 88334 373164 88340 373176
rect 54444 373136 88340 373164
rect 54444 373124 54450 373136
rect 88334 373124 88340 373136
rect 88392 373124 88398 373176
rect 156506 373124 156512 373176
rect 156564 373164 156570 373176
rect 203334 373164 203340 373176
rect 156564 373136 203340 373164
rect 156564 373124 156570 373136
rect 203334 373124 203340 373136
rect 203392 373124 203398 373176
rect 212626 373124 212632 373176
rect 212684 373164 212690 373176
rect 217962 373164 217968 373176
rect 212684 373136 217968 373164
rect 212684 373124 212690 373136
rect 217962 373124 217968 373136
rect 218020 373164 218026 373176
rect 255406 373164 255412 373176
rect 218020 373136 255412 373164
rect 218020 373124 218026 373136
rect 255406 373124 255412 373136
rect 255464 373124 255470 373176
rect 59722 373056 59728 373108
rect 59780 373096 59786 373108
rect 93670 373096 93676 373108
rect 59780 373068 93676 373096
rect 59780 373056 59786 373068
rect 93670 373056 93676 373068
rect 93728 373056 93734 373108
rect 212718 373056 212724 373108
rect 212776 373096 212782 373108
rect 219066 373096 219072 373108
rect 212776 373068 219072 373096
rect 212776 373056 212782 373068
rect 219066 373056 219072 373068
rect 219124 373096 219130 373108
rect 258074 373096 258080 373108
rect 219124 373068 258080 373096
rect 219124 373056 219130 373068
rect 258074 373056 258080 373068
rect 258132 373056 258138 373108
rect 212810 372988 212816 373040
rect 212868 373028 212874 373040
rect 213638 373028 213644 373040
rect 212868 373000 213644 373028
rect 212868 372988 212874 373000
rect 213638 372988 213644 373000
rect 213696 373028 213702 373040
rect 256694 373028 256700 373040
rect 213696 373000 256700 373028
rect 213696 372988 213702 373000
rect 256694 372988 256700 373000
rect 256752 372988 256758 373040
rect 214006 372920 214012 372972
rect 214064 372960 214070 372972
rect 259638 372960 259644 372972
rect 214064 372932 259644 372960
rect 214064 372920 214070 372932
rect 259638 372920 259644 372932
rect 259696 372920 259702 372972
rect 216950 372852 216956 372904
rect 217008 372892 217014 372904
rect 217594 372892 217600 372904
rect 217008 372864 217600 372892
rect 217008 372852 217014 372864
rect 217594 372852 217600 372864
rect 217652 372852 217658 372904
rect 259454 372892 259460 372904
rect 217704 372864 259460 372892
rect 100018 372784 100024 372836
rect 100076 372824 100082 372836
rect 213914 372824 213920 372836
rect 100076 372796 213920 372824
rect 100076 372784 100082 372796
rect 213914 372784 213920 372796
rect 213972 372824 213978 372836
rect 215202 372824 215208 372836
rect 213972 372796 215208 372824
rect 213972 372784 213978 372796
rect 215202 372784 215208 372796
rect 215260 372824 215266 372836
rect 217704 372824 217732 372864
rect 259454 372852 259460 372864
rect 259512 372852 259518 372904
rect 220722 372824 220728 372836
rect 215260 372796 217732 372824
rect 218072 372796 220728 372824
rect 215260 372784 215266 372796
rect 204254 372716 204260 372768
rect 204312 372756 204318 372768
rect 215294 372756 215300 372768
rect 204312 372728 215300 372756
rect 204312 372716 204318 372728
rect 215294 372716 215300 372728
rect 215352 372716 215358 372768
rect 207198 372648 207204 372700
rect 207256 372688 207262 372700
rect 215018 372688 215024 372700
rect 207256 372660 215024 372688
rect 207256 372648 207262 372660
rect 215018 372648 215024 372660
rect 215076 372648 215082 372700
rect 215386 372648 215392 372700
rect 215444 372688 215450 372700
rect 216398 372688 216404 372700
rect 215444 372660 216404 372688
rect 215444 372648 215450 372660
rect 216398 372648 216404 372660
rect 216456 372688 216462 372700
rect 218072 372688 218100 372796
rect 220722 372784 220728 372796
rect 220780 372784 220786 372836
rect 264974 372824 264980 372836
rect 220832 372796 264980 372824
rect 219250 372716 219256 372768
rect 219308 372756 219314 372768
rect 220832 372756 220860 372796
rect 264974 372784 264980 372796
rect 265032 372784 265038 372836
rect 219308 372728 220860 372756
rect 219308 372716 219314 372728
rect 220906 372716 220912 372768
rect 220964 372756 220970 372768
rect 266354 372756 266360 372768
rect 220964 372728 266360 372756
rect 220964 372716 220970 372728
rect 266354 372716 266360 372728
rect 266412 372716 266418 372768
rect 261294 372688 261300 372700
rect 216456 372660 218100 372688
rect 219406 372660 261300 372688
rect 216456 372648 216462 372660
rect 214098 372580 214104 372632
rect 214156 372620 214162 372632
rect 219406 372620 219434 372660
rect 261294 372648 261300 372660
rect 261352 372648 261358 372700
rect 380894 372648 380900 372700
rect 380952 372688 380958 372700
rect 426434 372688 426440 372700
rect 380952 372660 426440 372688
rect 380952 372648 380958 372660
rect 426434 372648 426440 372660
rect 426492 372648 426498 372700
rect 516686 372688 516692 372700
rect 509206 372660 516692 372688
rect 214156 372592 219434 372620
rect 214156 372580 214162 372592
rect 220722 372580 220728 372632
rect 220780 372620 220786 372632
rect 262214 372620 262220 372632
rect 220780 372592 262220 372620
rect 220780 372580 220786 372592
rect 262214 372580 262220 372592
rect 262272 372580 262278 372632
rect 275830 372580 275836 372632
rect 275888 372620 275894 372632
rect 356606 372620 356612 372632
rect 275888 372592 356612 372620
rect 275888 372580 275894 372592
rect 356606 372580 356612 372592
rect 356664 372580 356670 372632
rect 369762 372580 369768 372632
rect 369820 372620 369826 372632
rect 369820 372592 376524 372620
rect 369820 372580 369826 372592
rect 84746 372512 84752 372564
rect 84804 372552 84810 372564
rect 208486 372552 208492 372564
rect 84804 372524 208492 372552
rect 84804 372512 84810 372524
rect 208486 372512 208492 372524
rect 208544 372552 208550 372564
rect 210970 372552 210976 372564
rect 208544 372524 210976 372552
rect 208544 372512 208550 372524
rect 210970 372512 210976 372524
rect 211028 372512 211034 372564
rect 212718 372512 212724 372564
rect 212776 372552 212782 372564
rect 219434 372552 219440 372564
rect 212776 372524 219440 372552
rect 212776 372512 212782 372524
rect 219434 372512 219440 372524
rect 219492 372552 219498 372564
rect 273254 372552 273260 372564
rect 219492 372524 273260 372552
rect 219492 372512 219498 372524
rect 273254 372512 273260 372524
rect 273312 372512 273318 372564
rect 281442 372512 281448 372564
rect 281500 372552 281506 372564
rect 326062 372552 326068 372564
rect 281500 372524 326068 372552
rect 281500 372512 281506 372524
rect 326062 372512 326068 372524
rect 326120 372512 326126 372564
rect 370314 372512 370320 372564
rect 370372 372552 370378 372564
rect 375098 372552 375104 372564
rect 370372 372524 375104 372552
rect 370372 372512 370378 372524
rect 375098 372512 375104 372524
rect 375156 372512 375162 372564
rect 86770 372444 86776 372496
rect 86828 372484 86834 372496
rect 208394 372484 208400 372496
rect 86828 372456 208400 372484
rect 86828 372444 86834 372456
rect 208394 372444 208400 372456
rect 208452 372444 208458 372496
rect 210326 372444 210332 372496
rect 210384 372484 210390 372496
rect 218054 372484 218060 372496
rect 210384 372456 218060 372484
rect 210384 372444 210390 372456
rect 218054 372444 218060 372456
rect 218112 372484 218118 372496
rect 271874 372484 271880 372496
rect 218112 372456 271880 372484
rect 218112 372444 218118 372456
rect 271874 372444 271880 372456
rect 271932 372444 271938 372496
rect 376496 372484 376524 372592
rect 376846 372580 376852 372632
rect 376904 372620 376910 372632
rect 378042 372620 378048 372632
rect 376904 372592 378048 372620
rect 376904 372580 376910 372592
rect 378042 372580 378048 372592
rect 378100 372620 378106 372632
rect 425054 372620 425060 372632
rect 378100 372592 425060 372620
rect 378100 372580 378106 372592
rect 425054 372580 425060 372592
rect 425112 372580 425118 372632
rect 439406 372580 439412 372632
rect 439464 372620 439470 372632
rect 509206 372620 509234 372660
rect 516686 372648 516692 372660
rect 516744 372648 516750 372700
rect 439464 372592 509234 372620
rect 439464 372580 439470 372592
rect 511902 372580 511908 372632
rect 511960 372620 511966 372632
rect 517514 372620 517520 372632
rect 511960 372592 517520 372620
rect 511960 372580 511966 372592
rect 517514 372580 517520 372592
rect 517572 372580 517578 372632
rect 376570 372512 376576 372564
rect 376628 372552 376634 372564
rect 438210 372552 438216 372564
rect 376628 372524 438216 372552
rect 376628 372512 376634 372524
rect 438210 372512 438216 372524
rect 438268 372512 438274 372564
rect 376754 372484 376760 372496
rect 376496 372456 376760 372484
rect 376754 372444 376760 372456
rect 376812 372484 376818 372496
rect 427814 372484 427820 372496
rect 376812 372456 427820 372484
rect 376812 372444 376818 372456
rect 427814 372444 427820 372456
rect 427872 372444 427878 372496
rect 91554 372376 91560 372428
rect 91612 372416 91618 372428
rect 208412 372416 208440 372444
rect 213362 372416 213368 372428
rect 91612 372388 205634 372416
rect 208412 372388 213368 372416
rect 91612 372376 91618 372388
rect 92382 372308 92388 372360
rect 92440 372348 92446 372360
rect 204162 372348 204168 372360
rect 92440 372320 204168 372348
rect 92440 372308 92446 372320
rect 204162 372308 204168 372320
rect 204220 372308 204226 372360
rect 93394 372240 93400 372292
rect 93452 372280 93458 372292
rect 202782 372280 202788 372292
rect 93452 372252 202788 372280
rect 93452 372240 93458 372252
rect 202782 372240 202788 372252
rect 202840 372240 202846 372292
rect 52914 372172 52920 372224
rect 52972 372212 52978 372224
rect 54386 372212 54392 372224
rect 52972 372184 54392 372212
rect 52972 372172 52978 372184
rect 54386 372172 54392 372184
rect 54444 372172 54450 372224
rect 79502 372172 79508 372224
rect 79560 372212 79566 372224
rect 205606 372212 205634 372388
rect 213362 372376 213368 372388
rect 213420 372376 213426 372428
rect 368934 372308 368940 372360
rect 368992 372348 368998 372360
rect 379606 372348 379612 372360
rect 368992 372320 379612 372348
rect 368992 372308 368998 372320
rect 379606 372308 379612 372320
rect 379664 372308 379670 372360
rect 210970 372240 210976 372292
rect 211028 372280 211034 372292
rect 244274 372280 244280 372292
rect 211028 372252 244280 372280
rect 211028 372240 211034 372252
rect 244274 372240 244280 372252
rect 244332 372240 244338 372292
rect 211338 372212 211344 372224
rect 79560 372184 200114 372212
rect 205606 372184 211344 372212
rect 79560 372172 79566 372184
rect 200086 372144 200114 372184
rect 211338 372172 211344 372184
rect 211396 372212 211402 372224
rect 219894 372212 219900 372224
rect 211396 372184 219900 372212
rect 211396 372172 211402 372184
rect 219894 372172 219900 372184
rect 219952 372212 219958 372224
rect 220538 372212 220544 372224
rect 219952 372184 220544 372212
rect 219952 372172 219958 372184
rect 220538 372172 220544 372184
rect 220596 372172 220602 372224
rect 251174 372212 251180 372224
rect 229066 372184 251180 372212
rect 215294 372144 215300 372156
rect 200086 372116 215300 372144
rect 215294 372104 215300 372116
rect 215352 372104 215358 372156
rect 220446 372104 220452 372156
rect 220504 372144 220510 372156
rect 229066 372144 229094 372184
rect 251174 372172 251180 372184
rect 251232 372172 251238 372224
rect 220504 372116 229094 372144
rect 220504 372104 220510 372116
rect 373074 372104 373080 372156
rect 373132 372144 373138 372156
rect 379514 372144 379520 372156
rect 373132 372116 379520 372144
rect 373132 372104 373138 372116
rect 379514 372104 379520 372116
rect 379572 372104 379578 372156
rect 202782 372036 202788 372088
rect 202840 372076 202846 372088
rect 220814 372076 220820 372088
rect 202840 372048 220820 372076
rect 202840 372036 202846 372048
rect 220814 372036 220820 372048
rect 220872 372076 220878 372088
rect 221918 372076 221924 372088
rect 220872 372048 221924 372076
rect 220872 372036 220878 372048
rect 221918 372036 221924 372048
rect 221976 372036 221982 372088
rect 367554 372036 367560 372088
rect 367612 372076 367618 372088
rect 376754 372076 376760 372088
rect 367612 372048 376760 372076
rect 367612 372036 367618 372048
rect 376754 372036 376760 372048
rect 376812 372036 376818 372088
rect 112990 371968 112996 372020
rect 113048 372008 113054 372020
rect 210326 372008 210332 372020
rect 113048 371980 210332 372008
rect 113048 371968 113054 371980
rect 210326 371968 210332 371980
rect 210384 371968 210390 372020
rect 220630 371968 220636 372020
rect 220688 372008 220694 372020
rect 241238 372008 241244 372020
rect 220688 371980 241244 372008
rect 220688 371968 220694 371980
rect 241238 371968 241244 371980
rect 241296 371968 241302 372020
rect 379330 371968 379336 372020
rect 379388 372008 379394 372020
rect 396074 372008 396080 372020
rect 379388 371980 396080 372008
rect 379388 371968 379394 371980
rect 396074 371968 396080 371980
rect 396132 371968 396138 372020
rect 204162 371900 204168 371952
rect 204220 371940 204226 371952
rect 219526 371940 219532 371952
rect 204220 371912 219532 371940
rect 204220 371900 204226 371912
rect 219526 371900 219532 371912
rect 219584 371940 219590 371952
rect 220446 371940 220452 371952
rect 219584 371912 220452 371940
rect 219584 371900 219590 371912
rect 220446 371900 220452 371912
rect 220504 371900 220510 371952
rect 241146 371940 241152 371952
rect 222764 371912 241152 371940
rect 219802 371872 219808 371884
rect 212828 371844 219808 371872
rect 182726 371764 182732 371816
rect 182784 371804 182790 371816
rect 202966 371804 202972 371816
rect 182784 371776 202972 371804
rect 182784 371764 182790 371776
rect 202966 371764 202972 371776
rect 203024 371804 203030 371816
rect 204162 371804 204168 371816
rect 203024 371776 204168 371804
rect 203024 371764 203030 371776
rect 204162 371764 204168 371776
rect 204220 371764 204226 371816
rect 114462 371696 114468 371748
rect 114520 371736 114526 371748
rect 212718 371736 212724 371748
rect 114520 371708 212724 371736
rect 114520 371696 114526 371708
rect 212718 371696 212724 371708
rect 212776 371696 212782 371748
rect 88058 371628 88064 371680
rect 88116 371668 88122 371680
rect 211062 371668 211068 371680
rect 88116 371640 211068 371668
rect 88116 371628 88122 371640
rect 211062 371628 211068 371640
rect 211120 371628 211126 371680
rect 90910 371560 90916 371612
rect 90968 371600 90974 371612
rect 209866 371600 209872 371612
rect 90968 371572 209872 371600
rect 90968 371560 90974 371572
rect 209866 371560 209872 371572
rect 209924 371600 209930 371612
rect 212828 371600 212856 371844
rect 219802 371832 219808 371844
rect 219860 371872 219866 371884
rect 222764 371872 222792 371912
rect 241146 371900 241152 371912
rect 241204 371900 241210 371952
rect 371050 371900 371056 371952
rect 371108 371940 371114 371952
rect 398834 371940 398840 371952
rect 371108 371912 398840 371940
rect 371108 371900 371114 371912
rect 398834 371900 398840 371912
rect 398892 371900 398898 371952
rect 219860 371844 222792 371872
rect 219860 371832 219866 371844
rect 224218 371832 224224 371884
rect 224276 371872 224282 371884
rect 247126 371872 247132 371884
rect 224276 371844 247132 371872
rect 224276 371832 224282 371844
rect 247126 371832 247132 371844
rect 247184 371832 247190 371884
rect 372522 371832 372528 371884
rect 372580 371872 372586 371884
rect 405734 371872 405740 371884
rect 372580 371844 405740 371872
rect 372580 371832 372586 371844
rect 405734 371832 405740 371844
rect 405792 371832 405798 371884
rect 215294 371764 215300 371816
rect 215352 371804 215358 371816
rect 216306 371804 216312 371816
rect 215352 371776 216312 371804
rect 215352 371764 215358 371776
rect 216306 371764 216312 371776
rect 216364 371804 216370 371816
rect 239122 371804 239128 371816
rect 216364 371776 239128 371804
rect 216364 371764 216370 371776
rect 239122 371764 239128 371776
rect 239180 371804 239186 371816
rect 240042 371804 240048 371816
rect 239180 371776 240048 371804
rect 239180 371764 239186 371776
rect 240042 371764 240048 371776
rect 240100 371764 240106 371816
rect 369670 371804 369676 371816
rect 364306 371776 369676 371804
rect 213362 371696 213368 371748
rect 213420 371736 213426 371748
rect 245654 371736 245660 371748
rect 213420 371708 245660 371736
rect 213420 371696 213426 371708
rect 245654 371696 245660 371708
rect 245712 371696 245718 371748
rect 220538 371628 220544 371680
rect 220596 371668 220602 371680
rect 251174 371668 251180 371680
rect 220596 371640 251180 371668
rect 220596 371628 220602 371640
rect 251174 371628 251180 371640
rect 251232 371628 251238 371680
rect 274634 371628 274640 371680
rect 274692 371668 274698 371680
rect 302234 371668 302240 371680
rect 274692 371640 302240 371668
rect 274692 371628 274698 371640
rect 302234 371628 302240 371640
rect 302292 371628 302298 371680
rect 209924 371572 212856 371600
rect 209924 371560 209930 371572
rect 280062 371560 280068 371612
rect 280120 371600 280126 371612
rect 359274 371600 359280 371612
rect 280120 371572 359280 371600
rect 280120 371560 280126 371572
rect 359274 371560 359280 371572
rect 359332 371560 359338 371612
rect 89346 371492 89352 371544
rect 89404 371532 89410 371544
rect 209958 371532 209964 371544
rect 89404 371504 209964 371532
rect 89404 371492 89410 371504
rect 209958 371492 209964 371504
rect 210016 371532 210022 371544
rect 219710 371532 219716 371544
rect 210016 371504 219716 371532
rect 210016 371492 210022 371504
rect 219710 371492 219716 371504
rect 219768 371532 219774 371544
rect 220630 371532 220636 371544
rect 219768 371504 220636 371532
rect 219768 371492 219774 371504
rect 220630 371492 220636 371504
rect 220688 371492 220694 371544
rect 221918 371492 221924 371544
rect 221976 371532 221982 371544
rect 252554 371532 252560 371544
rect 221976 371504 252560 371532
rect 221976 371492 221982 371504
rect 252554 371492 252560 371504
rect 252612 371492 252618 371544
rect 276014 371492 276020 371544
rect 276072 371532 276078 371544
rect 356974 371532 356980 371544
rect 276072 371504 356980 371532
rect 276072 371492 276078 371504
rect 356974 371492 356980 371504
rect 357032 371492 357038 371544
rect 44634 371424 44640 371476
rect 44692 371464 44698 371476
rect 47486 371464 47492 371476
rect 44692 371436 47492 371464
rect 44692 371424 44698 371436
rect 47486 371424 47492 371436
rect 47544 371464 47550 371476
rect 78306 371464 78312 371476
rect 47544 371436 78312 371464
rect 47544 371424 47550 371436
rect 78306 371424 78312 371436
rect 78364 371464 78370 371476
rect 364306 371464 364334 371776
rect 369670 371764 369676 371776
rect 369728 371804 369734 371816
rect 397454 371804 397460 371816
rect 369728 371776 397460 371804
rect 369728 371764 369734 371776
rect 397454 371764 397460 371776
rect 397512 371764 397518 371816
rect 379606 371696 379612 371748
rect 379664 371736 379670 371748
rect 379790 371736 379796 371748
rect 379664 371708 379796 371736
rect 379664 371696 379670 371708
rect 379790 371696 379796 371708
rect 379848 371736 379854 371748
rect 409874 371736 409880 371748
rect 379848 371708 409880 371736
rect 379848 371696 379854 371708
rect 409874 371696 409880 371708
rect 409932 371696 409938 371748
rect 374546 371628 374552 371680
rect 374604 371668 374610 371680
rect 380066 371668 380072 371680
rect 374604 371640 380072 371668
rect 374604 371628 374610 371640
rect 380066 371628 380072 371640
rect 380124 371668 380130 371680
rect 411254 371668 411260 371680
rect 380124 371640 411260 371668
rect 380124 371628 380130 371640
rect 411254 371628 411260 371640
rect 411312 371628 411318 371680
rect 375098 371560 375104 371612
rect 375156 371600 375162 371612
rect 407114 371600 407120 371612
rect 375156 371572 407120 371600
rect 375156 371560 375162 371572
rect 407114 371560 407120 371572
rect 407172 371560 407178 371612
rect 379514 371492 379520 371544
rect 379572 371532 379578 371544
rect 379882 371532 379888 371544
rect 379572 371504 379888 371532
rect 379572 371492 379578 371504
rect 379882 371492 379888 371504
rect 379940 371532 379946 371544
rect 412634 371532 412640 371544
rect 379940 371504 412640 371532
rect 379940 371492 379946 371504
rect 412634 371492 412640 371504
rect 412692 371492 412698 371544
rect 78364 371436 200114 371464
rect 78364 371424 78370 371436
rect 44726 371356 44732 371408
rect 44784 371396 44790 371408
rect 47578 371396 47584 371408
rect 44784 371368 47584 371396
rect 44784 371356 44790 371368
rect 47578 371356 47584 371368
rect 47636 371396 47642 371408
rect 80054 371396 80060 371408
rect 47636 371368 80060 371396
rect 47636 371356 47642 371368
rect 80054 371356 80060 371368
rect 80112 371356 80118 371408
rect 200086 371396 200114 371436
rect 238726 371436 364334 371464
rect 210878 371396 210884 371408
rect 200086 371368 210884 371396
rect 210878 371356 210884 371368
rect 210936 371396 210942 371408
rect 238110 371396 238116 371408
rect 210936 371368 238116 371396
rect 210936 371356 210942 371368
rect 238110 371356 238116 371368
rect 238168 371396 238174 371408
rect 238726 371396 238754 371436
rect 373166 371424 373172 371476
rect 373224 371464 373230 371476
rect 373718 371464 373724 371476
rect 373224 371436 373724 371464
rect 373224 371424 373230 371436
rect 373718 371424 373724 371436
rect 373776 371424 373782 371476
rect 376754 371424 376760 371476
rect 376812 371464 376818 371476
rect 378042 371464 378048 371476
rect 376812 371436 378048 371464
rect 376812 371424 376818 371436
rect 378042 371424 378048 371436
rect 378100 371464 378106 371476
rect 411254 371464 411260 371476
rect 378100 371436 411260 371464
rect 378100 371424 378106 371436
rect 411254 371424 411260 371436
rect 411312 371424 411318 371476
rect 238168 371368 238754 371396
rect 238168 371356 238174 371368
rect 240042 371356 240048 371408
rect 240100 371396 240106 371408
rect 371050 371396 371056 371408
rect 240100 371368 371056 371396
rect 240100 371356 240106 371368
rect 371050 371356 371056 371368
rect 371108 371356 371114 371408
rect 379974 371356 379980 371408
rect 380032 371396 380038 371408
rect 380986 371396 380992 371408
rect 380032 371368 380992 371396
rect 380032 371356 380038 371368
rect 380986 371356 380992 371368
rect 381044 371396 381050 371408
rect 422294 371396 422300 371408
rect 381044 371368 422300 371396
rect 381044 371356 381050 371368
rect 422294 371356 422300 371368
rect 422352 371356 422358 371408
rect 438210 371356 438216 371408
rect 438268 371396 438274 371408
rect 516594 371396 516600 371408
rect 438268 371368 516600 371396
rect 438268 371356 438274 371368
rect 516594 371356 516600 371368
rect 516652 371356 516658 371408
rect 44818 371288 44824 371340
rect 44876 371328 44882 371340
rect 46106 371328 46112 371340
rect 44876 371300 46112 371328
rect 44876 371288 44882 371300
rect 46106 371288 46112 371300
rect 46164 371328 46170 371340
rect 79502 371328 79508 371340
rect 46164 371300 79508 371328
rect 46164 371288 46170 371300
rect 79502 371288 79508 371300
rect 79560 371288 79566 371340
rect 204162 371288 204168 371340
rect 204220 371328 204226 371340
rect 343174 371328 343180 371340
rect 204220 371300 343180 371328
rect 204220 371288 204226 371300
rect 343174 371288 343180 371300
rect 343232 371328 343238 371340
rect 360286 371328 360292 371340
rect 343232 371300 360292 371328
rect 343232 371288 343238 371300
rect 360286 371288 360292 371300
rect 360344 371328 360350 371340
rect 503162 371328 503168 371340
rect 360344 371300 503168 371328
rect 360344 371288 360350 371300
rect 503162 371288 503168 371300
rect 503220 371328 503226 371340
rect 517882 371328 517888 371340
rect 503220 371300 517888 371328
rect 503220 371288 503226 371300
rect 517882 371288 517888 371300
rect 517940 371288 517946 371340
rect 44910 371220 44916 371272
rect 44968 371260 44974 371272
rect 47854 371260 47860 371272
rect 44968 371232 47860 371260
rect 44968 371220 44974 371232
rect 47854 371220 47860 371232
rect 47912 371260 47918 371272
rect 81434 371260 81440 371272
rect 47912 371232 81440 371260
rect 47912 371220 47918 371232
rect 81434 371220 81440 371232
rect 81492 371220 81498 371272
rect 84562 371220 84568 371272
rect 84620 371260 84626 371272
rect 106182 371260 106188 371272
rect 84620 371232 106188 371260
rect 84620 371220 84626 371232
rect 106182 371220 106188 371232
rect 106240 371220 106246 371272
rect 201586 371260 201592 371272
rect 183480 371232 201592 371260
rect 3510 371152 3516 371204
rect 3568 371192 3574 371204
rect 40678 371192 40684 371204
rect 3568 371164 40684 371192
rect 3568 371152 3574 371164
rect 40678 371152 40684 371164
rect 40736 371152 40742 371204
rect 47670 371152 47676 371204
rect 47728 371192 47734 371204
rect 183278 371192 183284 371204
rect 47728 371164 183284 371192
rect 47728 371152 47734 371164
rect 183278 371152 183284 371164
rect 183336 371192 183342 371204
rect 183480 371192 183508 371232
rect 201586 371220 201592 371232
rect 201644 371260 201650 371272
rect 343450 371260 343456 371272
rect 201644 371232 343456 371260
rect 201644 371220 201650 371232
rect 343450 371220 343456 371232
rect 343508 371260 343514 371272
rect 357434 371260 357440 371272
rect 343508 371232 357440 371260
rect 343508 371220 343514 371232
rect 357434 371220 357440 371232
rect 357492 371260 357498 371272
rect 502334 371260 502340 371272
rect 357492 371232 502340 371260
rect 357492 371220 357498 371232
rect 502334 371220 502340 371232
rect 502392 371220 502398 371272
rect 183336 371164 183508 371192
rect 183336 371152 183342 371164
rect 198826 371152 198832 371204
rect 198884 371192 198890 371204
rect 304994 371192 305000 371204
rect 198884 371164 305000 371192
rect 198884 371152 198890 371164
rect 304994 371152 305000 371164
rect 305052 371152 305058 371204
rect 357894 371152 357900 371204
rect 357952 371192 357958 371204
rect 473354 371192 473360 371204
rect 357952 371164 473360 371192
rect 357952 371152 357958 371164
rect 473354 371152 473360 371164
rect 473412 371152 473418 371204
rect 47762 371084 47768 371136
rect 47820 371124 47826 371136
rect 182726 371124 182732 371136
rect 47820 371096 182732 371124
rect 47820 371084 47826 371096
rect 182726 371084 182732 371096
rect 182784 371084 182790 371136
rect 197538 371084 197544 371136
rect 197596 371124 197602 371136
rect 298094 371124 298100 371136
rect 197596 371096 298100 371124
rect 197596 371084 197602 371096
rect 298094 371084 298100 371096
rect 298152 371084 298158 371136
rect 357342 371084 357348 371136
rect 357400 371124 357406 371136
rect 470594 371124 470600 371136
rect 357400 371096 470600 371124
rect 357400 371084 357406 371096
rect 470594 371084 470600 371096
rect 470652 371084 470658 371136
rect 104618 371016 104624 371068
rect 104676 371056 104682 371068
rect 215478 371056 215484 371068
rect 104676 371028 215484 371056
rect 104676 371016 104682 371028
rect 215478 371016 215484 371028
rect 215536 371016 215542 371068
rect 217410 371016 217416 371068
rect 217468 371056 217474 371068
rect 307754 371056 307760 371068
rect 217468 371028 307760 371056
rect 217468 371016 217474 371028
rect 307754 371016 307760 371028
rect 307812 371016 307818 371068
rect 366266 371016 366272 371068
rect 366324 371056 366330 371068
rect 465074 371056 465080 371068
rect 366324 371028 465080 371056
rect 366324 371016 366330 371028
rect 465074 371016 465080 371028
rect 465132 371016 465138 371068
rect 196710 370948 196716 371000
rect 196768 370988 196774 371000
rect 287238 370988 287244 371000
rect 196768 370960 287244 370988
rect 196768 370948 196774 370960
rect 287238 370948 287244 370960
rect 287296 370948 287302 371000
rect 369026 370948 369032 371000
rect 369084 370988 369090 371000
rect 467834 370988 467840 371000
rect 369084 370960 467840 370988
rect 369084 370948 369090 370960
rect 467834 370948 467840 370960
rect 467892 370948 467898 371000
rect 202414 370880 202420 370932
rect 202472 370920 202478 370932
rect 300854 370920 300860 370932
rect 202472 370892 300860 370920
rect 202472 370880 202478 370892
rect 300854 370880 300860 370892
rect 300912 370880 300918 370932
rect 358722 370880 358728 370932
rect 358780 370920 358786 370932
rect 437474 370920 437480 370932
rect 358780 370892 437480 370920
rect 358780 370880 358786 370892
rect 437474 370880 437480 370892
rect 437532 370880 437538 370932
rect 197446 370812 197452 370864
rect 197504 370852 197510 370864
rect 295334 370852 295340 370864
rect 197504 370824 295340 370852
rect 197504 370812 197510 370824
rect 295334 370812 295340 370824
rect 295392 370812 295398 370864
rect 359642 370812 359648 370864
rect 359700 370852 359706 370864
rect 415394 370852 415400 370864
rect 359700 370824 415400 370852
rect 359700 370812 359706 370824
rect 415394 370812 415400 370824
rect 415452 370812 415458 370864
rect 198274 370744 198280 370796
rect 198332 370784 198338 370796
rect 292574 370784 292580 370796
rect 198332 370756 292580 370784
rect 198332 370744 198338 370756
rect 292574 370744 292580 370756
rect 292632 370744 292638 370796
rect 361390 370744 361396 370796
rect 361448 370784 361454 370796
rect 412818 370784 412824 370796
rect 361448 370756 412824 370784
rect 361448 370744 361454 370756
rect 412818 370744 412824 370756
rect 412876 370744 412882 370796
rect 196802 370676 196808 370728
rect 196860 370716 196866 370728
rect 289814 370716 289820 370728
rect 196860 370688 289820 370716
rect 196860 370676 196866 370688
rect 289814 370676 289820 370688
rect 289872 370676 289878 370728
rect 368290 370676 368296 370728
rect 368348 370716 368354 370728
rect 374546 370716 374552 370728
rect 368348 370688 374552 370716
rect 368348 370676 368354 370688
rect 374546 370676 374552 370688
rect 374604 370676 374610 370728
rect 377122 370676 377128 370728
rect 377180 370716 377186 370728
rect 416774 370716 416780 370728
rect 377180 370688 416780 370716
rect 377180 370676 377186 370688
rect 416774 370676 416780 370688
rect 416832 370676 416838 370728
rect 196618 370608 196624 370660
rect 196676 370648 196682 370660
rect 285674 370648 285680 370660
rect 196676 370620 285680 370648
rect 196676 370608 196682 370620
rect 285674 370608 285680 370620
rect 285732 370608 285738 370660
rect 373074 370608 373080 370660
rect 373132 370648 373138 370660
rect 379606 370648 379612 370660
rect 373132 370620 379612 370648
rect 373132 370608 373138 370620
rect 379606 370608 379612 370620
rect 379664 370648 379670 370660
rect 414014 370648 414020 370660
rect 379664 370620 414020 370648
rect 379664 370608 379670 370620
rect 414014 370608 414020 370620
rect 414072 370608 414078 370660
rect 196986 370540 196992 370592
rect 197044 370580 197050 370592
rect 277394 370580 277400 370592
rect 197044 370552 277400 370580
rect 197044 370540 197050 370552
rect 277394 370540 277400 370552
rect 277452 370540 277458 370592
rect 374546 370540 374552 370592
rect 374604 370580 374610 370592
rect 396074 370580 396080 370592
rect 374604 370552 396080 370580
rect 374604 370540 374610 370552
rect 396074 370540 396080 370552
rect 396132 370540 396138 370592
rect 52914 370472 52920 370524
rect 52972 370512 52978 370524
rect 58618 370512 58624 370524
rect 52972 370484 58624 370512
rect 52972 370472 52978 370484
rect 58618 370472 58624 370484
rect 58676 370472 58682 370524
rect 198734 370472 198740 370524
rect 198792 370512 198798 370524
rect 274634 370512 274640 370524
rect 198792 370484 274640 370512
rect 198792 370472 198798 370484
rect 274634 370472 274640 370484
rect 274692 370472 274698 370524
rect 374454 370472 374460 370524
rect 374512 370512 374518 370524
rect 377122 370512 377128 370524
rect 374512 370484 377128 370512
rect 374512 370472 374518 370484
rect 377122 370472 377128 370484
rect 377180 370472 377186 370524
rect 402974 370512 402980 370524
rect 377232 370484 402980 370512
rect 206830 370404 206836 370456
rect 206888 370444 206894 370456
rect 270494 370444 270500 370456
rect 206888 370416 270500 370444
rect 206888 370404 206894 370416
rect 270494 370404 270500 370416
rect 270552 370404 270558 370456
rect 106182 370336 106188 370388
rect 106240 370376 106246 370388
rect 106240 370348 205634 370376
rect 106240 370336 106246 370348
rect 205606 370240 205634 370348
rect 212442 370336 212448 370388
rect 212500 370376 212506 370388
rect 276014 370376 276020 370388
rect 212500 370348 276020 370376
rect 212500 370336 212506 370348
rect 276014 370336 276020 370348
rect 276072 370336 276078 370388
rect 370406 370336 370412 370388
rect 370464 370376 370470 370388
rect 376662 370376 376668 370388
rect 370464 370348 376668 370376
rect 370464 370336 370470 370348
rect 376662 370336 376668 370348
rect 376720 370376 376726 370388
rect 377232 370376 377260 370484
rect 402974 370472 402980 370484
rect 403032 370472 403038 370524
rect 403250 370376 403256 370388
rect 376720 370348 377260 370376
rect 379486 370348 403256 370376
rect 376720 370336 376726 370348
rect 208026 370268 208032 370320
rect 208084 370308 208090 370320
rect 264974 370308 264980 370320
rect 208084 370280 264980 370308
rect 208084 370268 208090 370280
rect 264974 370268 264980 370280
rect 265032 370268 265038 370320
rect 371786 370268 371792 370320
rect 371844 370308 371850 370320
rect 377490 370308 377496 370320
rect 371844 370280 377496 370308
rect 371844 370268 371850 370280
rect 377490 370268 377496 370280
rect 377548 370308 377554 370320
rect 379486 370308 379514 370348
rect 403250 370336 403256 370348
rect 403308 370336 403314 370388
rect 377548 370280 379514 370308
rect 377548 370268 377554 370280
rect 208578 370240 208584 370252
rect 205606 370212 208584 370240
rect 208578 370200 208584 370212
rect 208636 370240 208642 370252
rect 213546 370240 213552 370252
rect 208636 370212 213552 370240
rect 208636 370200 208642 370212
rect 213546 370200 213552 370212
rect 213604 370200 213610 370252
rect 215478 369860 215484 369912
rect 215536 369900 215542 369912
rect 217226 369900 217232 369912
rect 215536 369872 217232 369900
rect 215536 369860 215542 369872
rect 217226 369860 217232 369872
rect 217284 369860 217290 369912
rect 202874 369792 202880 369844
rect 202932 369832 202938 369844
rect 322934 369832 322940 369844
rect 202932 369804 322940 369832
rect 202932 369792 202938 369804
rect 322934 369792 322940 369804
rect 322992 369792 322998 369844
rect 357986 369792 357992 369844
rect 358044 369832 358050 369844
rect 485774 369832 485780 369844
rect 358044 369804 485780 369832
rect 358044 369792 358050 369804
rect 485774 369792 485780 369804
rect 485832 369792 485838 369844
rect 200666 369724 200672 369776
rect 200724 369764 200730 369776
rect 313274 369764 313280 369776
rect 200724 369736 313280 369764
rect 200724 369724 200730 369736
rect 313274 369724 313280 369736
rect 313332 369724 313338 369776
rect 357250 369724 357256 369776
rect 357308 369764 357314 369776
rect 483014 369764 483020 369776
rect 357308 369736 483020 369764
rect 357308 369724 357314 369736
rect 483014 369724 483020 369736
rect 483072 369724 483078 369776
rect 200206 369656 200212 369708
rect 200264 369696 200270 369708
rect 310514 369696 310520 369708
rect 200264 369668 310520 369696
rect 200264 369656 200270 369668
rect 310514 369656 310520 369668
rect 310572 369656 310578 369708
rect 375742 369656 375748 369708
rect 375800 369696 375806 369708
rect 480254 369696 480260 369708
rect 375800 369668 480260 369696
rect 375800 369656 375806 369668
rect 480254 369656 480260 369668
rect 480312 369656 480318 369708
rect 203518 369588 203524 369640
rect 203576 369628 203582 369640
rect 280154 369628 280160 369640
rect 203576 369600 280160 369628
rect 203576 369588 203582 369600
rect 280154 369588 280160 369600
rect 280212 369588 280218 369640
rect 364886 369588 364892 369640
rect 364944 369628 364950 369640
rect 430574 369628 430580 369640
rect 364944 369600 430580 369628
rect 364944 369588 364950 369600
rect 430574 369588 430580 369600
rect 430632 369588 430638 369640
rect 76834 369520 76840 369572
rect 76892 369560 76898 369572
rect 203058 369560 203064 369572
rect 76892 369532 203064 369560
rect 76892 369520 76898 369532
rect 203058 369520 203064 369532
rect 203116 369520 203122 369572
rect 211522 369520 211528 369572
rect 211580 369560 211586 369572
rect 282914 369560 282920 369572
rect 211580 369532 282920 369560
rect 211580 369520 211586 369532
rect 282914 369520 282920 369532
rect 282972 369520 282978 369572
rect 362770 369520 362776 369572
rect 362828 369560 362834 369572
rect 427814 369560 427820 369572
rect 362828 369532 427820 369560
rect 362828 369520 362834 369532
rect 427814 369520 427820 369532
rect 427872 369520 427878 369572
rect 205358 369452 205364 369504
rect 205416 369492 205422 369504
rect 267734 369492 267740 369504
rect 205416 369464 267740 369492
rect 205416 369452 205422 369464
rect 267734 369452 267740 369464
rect 267792 369452 267798 369504
rect 376478 369452 376484 369504
rect 376536 369492 376542 369504
rect 418154 369492 418160 369504
rect 376536 369464 418160 369492
rect 376536 369452 376542 369464
rect 418154 369452 418160 369464
rect 418212 369452 418218 369504
rect 77202 369384 77208 369436
rect 77260 369424 77266 369436
rect 204254 369424 204260 369436
rect 77260 369396 204260 369424
rect 77260 369384 77266 369396
rect 204254 369384 204260 369396
rect 204312 369384 204318 369436
rect 212902 369384 212908 369436
rect 212960 369424 212966 369436
rect 258166 369424 258172 369436
rect 212960 369396 258172 369424
rect 212960 369384 212966 369396
rect 258166 369384 258172 369396
rect 258224 369384 258230 369436
rect 373718 369384 373724 369436
rect 373776 369424 373782 369436
rect 373902 369424 373908 369436
rect 373776 369396 373908 369424
rect 373776 369384 373782 369396
rect 373902 369384 373908 369396
rect 373960 369384 373966 369436
rect 377214 369384 377220 369436
rect 377272 369424 377278 369436
rect 378686 369424 378692 369436
rect 377272 369396 378692 369424
rect 377272 369384 377278 369396
rect 378686 369384 378692 369396
rect 378744 369424 378750 369436
rect 415670 369424 415676 369436
rect 378744 369396 415676 369424
rect 378744 369384 378750 369396
rect 415670 369384 415676 369396
rect 415728 369384 415734 369436
rect 108850 369316 108856 369368
rect 108908 369356 108914 369368
rect 208118 369356 208124 369368
rect 108908 369328 208124 369356
rect 108908 369316 108914 369328
rect 208118 369316 208124 369328
rect 208176 369316 208182 369368
rect 208854 369316 208860 369368
rect 208912 369356 208918 369368
rect 273254 369356 273260 369368
rect 208912 369328 273260 369356
rect 208912 369316 208918 369328
rect 273254 369316 273260 369328
rect 273312 369316 273318 369368
rect 357158 369316 357164 369368
rect 357216 369356 357222 369368
rect 379330 369356 379336 369368
rect 357216 369328 379336 369356
rect 357216 369316 357222 369328
rect 379330 369316 379336 369328
rect 379388 369356 379394 369368
rect 419534 369356 419540 369368
rect 379388 369328 419540 369356
rect 379388 369316 379394 369328
rect 419534 369316 419540 369328
rect 419592 369316 419598 369368
rect 111610 369248 111616 369300
rect 111668 369288 111674 369300
rect 208946 369288 208952 369300
rect 111668 369260 208952 369288
rect 111668 369248 111674 369260
rect 208946 369248 208952 369260
rect 209004 369248 209010 369300
rect 218422 369248 218428 369300
rect 218480 369288 218486 369300
rect 263594 369288 263600 369300
rect 218480 369260 263600 369288
rect 218480 369248 218486 369260
rect 263594 369248 263600 369260
rect 263652 369248 263658 369300
rect 418246 369288 418252 369300
rect 373966 369260 418252 369288
rect 201034 369180 201040 369232
rect 201092 369220 201098 369232
rect 249794 369220 249800 369232
rect 201092 369192 249800 369220
rect 201092 369180 201098 369192
rect 249794 369180 249800 369192
rect 249852 369180 249858 369232
rect 360654 369180 360660 369232
rect 360712 369220 360718 369232
rect 373074 369220 373080 369232
rect 360712 369192 373080 369220
rect 360712 369180 360718 369192
rect 373074 369180 373080 369192
rect 373132 369220 373138 369232
rect 373966 369220 373994 369260
rect 418246 369248 418252 369260
rect 418304 369248 418310 369300
rect 373132 369192 373994 369220
rect 373132 369180 373138 369192
rect 375834 369180 375840 369232
rect 375892 369220 375898 369232
rect 376478 369220 376484 369232
rect 375892 369192 376484 369220
rect 375892 369180 375898 369192
rect 376478 369180 376484 369192
rect 376536 369180 376542 369232
rect 423674 369220 423680 369232
rect 377876 369192 423680 369220
rect 102042 369112 102048 369164
rect 102100 369152 102106 369164
rect 214098 369152 214104 369164
rect 102100 369124 214104 369152
rect 102100 369112 102106 369124
rect 214098 369112 214104 369124
rect 214156 369152 214162 369164
rect 214466 369152 214472 369164
rect 214156 369124 214472 369152
rect 214156 369112 214162 369124
rect 214466 369112 214472 369124
rect 214524 369112 214530 369164
rect 215846 369112 215852 369164
rect 215904 369152 215910 369164
rect 260834 369152 260840 369164
rect 215904 369124 260840 369152
rect 215904 369112 215910 369124
rect 260834 369112 260840 369124
rect 260892 369112 260898 369164
rect 371142 369112 371148 369164
rect 371200 369152 371206 369164
rect 375926 369152 375932 369164
rect 371200 369124 375932 369152
rect 371200 369112 371206 369124
rect 375926 369112 375932 369124
rect 375984 369152 375990 369164
rect 377876 369152 377904 369192
rect 423674 369180 423680 369192
rect 423732 369180 423738 369232
rect 431954 369152 431960 369164
rect 375984 369124 377904 369152
rect 383626 369124 431960 369152
rect 375984 369112 375990 369124
rect 83826 369044 83832 369096
rect 83884 369084 83890 369096
rect 207198 369084 207204 369096
rect 83884 369056 207204 369084
rect 83884 369044 83890 369056
rect 207198 369044 207204 369056
rect 207256 369044 207262 369096
rect 214374 369044 214380 369096
rect 214432 369084 214438 369096
rect 255314 369084 255320 369096
rect 214432 369056 255320 369084
rect 214432 369044 214438 369056
rect 255314 369044 255320 369056
rect 255372 369044 255378 369096
rect 369578 369044 369584 369096
rect 369636 369084 369642 369096
rect 371786 369084 371792 369096
rect 369636 369056 371792 369084
rect 369636 369044 369642 369056
rect 371786 369044 371792 369056
rect 371844 369084 371850 369096
rect 383626 369084 383654 369124
rect 431954 369112 431960 369124
rect 432012 369112 432018 369164
rect 371844 369056 383654 369084
rect 371844 369044 371850 369056
rect 210234 368976 210240 369028
rect 210292 369016 210298 369028
rect 247034 369016 247040 369028
rect 210292 368988 247040 369016
rect 210292 368976 210298 368988
rect 247034 368976 247040 368988
rect 247092 368976 247098 369028
rect 101674 368908 101680 368960
rect 101732 368948 101738 368960
rect 214006 368948 214012 368960
rect 101732 368920 214012 368948
rect 101732 368908 101738 368920
rect 214006 368908 214012 368920
rect 214064 368948 214070 368960
rect 215294 368948 215300 368960
rect 214064 368920 215300 368948
rect 214064 368908 214070 368920
rect 215294 368908 215300 368920
rect 215352 368908 215358 368960
rect 217502 368908 217508 368960
rect 217560 368948 217566 368960
rect 252646 368948 252652 368960
rect 217560 368920 252652 368948
rect 217560 368908 217566 368920
rect 252646 368908 252652 368920
rect 252704 368908 252710 368960
rect 102778 368840 102784 368892
rect 102836 368880 102842 368892
rect 216398 368880 216404 368892
rect 102836 368852 216404 368880
rect 102836 368840 102842 368852
rect 216398 368840 216404 368852
rect 216456 368840 216462 368892
rect 105630 368772 105636 368824
rect 105688 368812 105694 368824
rect 215570 368812 215576 368824
rect 105688 368784 215576 368812
rect 105688 368772 105694 368784
rect 215570 368772 215576 368784
rect 215628 368772 215634 368824
rect 376570 368432 376576 368484
rect 376628 368472 376634 368484
rect 379698 368472 379704 368484
rect 376628 368444 379704 368472
rect 376628 368432 376634 368444
rect 379698 368432 379704 368444
rect 379756 368472 379762 368484
rect 436094 368472 436100 368484
rect 379756 368444 436100 368472
rect 379756 368432 379762 368444
rect 436094 368432 436100 368444
rect 436152 368432 436158 368484
rect 379790 368228 379796 368280
rect 379848 368268 379854 368280
rect 380066 368268 380072 368280
rect 379848 368240 380072 368268
rect 379848 368228 379854 368240
rect 380066 368228 380072 368240
rect 380124 368228 380130 368280
rect 358998 367956 359004 368008
rect 359056 367996 359062 368008
rect 359550 367996 359556 368008
rect 359056 367968 359556 367996
rect 359056 367956 359062 367968
rect 359550 367956 359556 367968
rect 359608 367956 359614 368008
rect 373166 367956 373172 368008
rect 373224 367996 373230 368008
rect 376478 367996 376484 368008
rect 373224 367968 376484 367996
rect 373224 367956 373230 367968
rect 376478 367956 376484 367968
rect 376536 367996 376542 368008
rect 408494 367996 408500 368008
rect 376536 367968 408500 367996
rect 376536 367956 376542 367968
rect 408494 367956 408500 367968
rect 408552 367956 408558 368008
rect 362678 367888 362684 367940
rect 362736 367928 362742 367940
rect 379422 367928 379428 367940
rect 362736 367900 379428 367928
rect 362736 367888 362742 367900
rect 379422 367888 379428 367900
rect 379480 367928 379486 367940
rect 426434 367928 426440 367940
rect 379480 367900 426440 367928
rect 379480 367888 379486 367900
rect 426434 367888 426440 367900
rect 426492 367888 426498 367940
rect 364150 367820 364156 367872
rect 364208 367860 364214 367872
rect 374454 367860 374460 367872
rect 364208 367832 374460 367860
rect 364208 367820 364214 367832
rect 374454 367820 374460 367832
rect 374512 367860 374518 367872
rect 429194 367860 429200 367872
rect 374512 367832 429200 367860
rect 374512 367820 374518 367832
rect 429194 367820 429200 367832
rect 429252 367820 429258 367872
rect 199378 367752 199384 367804
rect 199436 367792 199442 367804
rect 358998 367792 359004 367804
rect 199436 367764 359004 367792
rect 199436 367752 199442 367764
rect 358998 367752 359004 367764
rect 359056 367752 359062 367804
rect 366910 367752 366916 367804
rect 366968 367792 366974 367804
rect 371142 367792 371148 367804
rect 366968 367764 371148 367792
rect 366968 367752 366974 367764
rect 371142 367752 371148 367764
rect 371200 367792 371206 367804
rect 430666 367792 430672 367804
rect 371200 367764 430672 367792
rect 371200 367752 371206 367764
rect 430666 367752 430672 367764
rect 430724 367752 430730 367804
rect 359918 366324 359924 366376
rect 359976 366364 359982 366376
rect 519354 366364 519360 366376
rect 359976 366336 519360 366364
rect 359976 366324 359982 366336
rect 519354 366324 519360 366336
rect 519412 366324 519418 366376
rect 199838 363604 199844 363656
rect 199896 363644 199902 363656
rect 358906 363644 358912 363656
rect 199896 363616 358912 363644
rect 199896 363604 199902 363616
rect 358906 363604 358912 363616
rect 358964 363604 358970 363656
rect 359826 360816 359832 360868
rect 359884 360856 359890 360868
rect 519078 360856 519084 360868
rect 359884 360828 519084 360856
rect 359884 360816 359890 360828
rect 519078 360816 519084 360828
rect 519136 360856 519142 360868
rect 519630 360856 519636 360868
rect 519136 360828 519636 360856
rect 519136 360816 519142 360828
rect 519630 360816 519636 360828
rect 519688 360816 519694 360868
rect 358906 359524 358912 359576
rect 358964 359564 358970 359576
rect 359642 359564 359648 359576
rect 358964 359536 359648 359564
rect 358964 359524 358970 359536
rect 359642 359524 359648 359536
rect 359700 359564 359706 359576
rect 519170 359564 519176 359576
rect 359700 359536 519176 359564
rect 359700 359524 359706 359536
rect 519170 359524 519176 359536
rect 519228 359564 519234 359576
rect 519354 359564 519360 359576
rect 519228 359536 519360 359564
rect 519228 359524 519234 359536
rect 519354 359524 519360 359536
rect 519412 359524 519418 359576
rect 199562 359456 199568 359508
rect 199620 359496 199626 359508
rect 199746 359496 199752 359508
rect 199620 359468 199752 359496
rect 199620 359456 199626 359468
rect 199746 359456 199752 359468
rect 199804 359496 199810 359508
rect 359090 359496 359096 359508
rect 199804 359468 359096 359496
rect 199804 359456 199810 359468
rect 359090 359456 359096 359468
rect 359148 359496 359154 359508
rect 359918 359496 359924 359508
rect 359148 359468 359924 359496
rect 359148 359456 359154 359468
rect 359918 359456 359924 359468
rect 359976 359456 359982 359508
rect 359182 358708 359188 358760
rect 359240 358748 359246 358760
rect 359458 358748 359464 358760
rect 359240 358720 359464 358748
rect 359240 358708 359246 358720
rect 359458 358708 359464 358720
rect 359516 358708 359522 358760
rect 359458 358028 359464 358080
rect 359516 358068 359522 358080
rect 519262 358068 519268 358080
rect 359516 358040 519268 358068
rect 359516 358028 359522 358040
rect 519262 358028 519268 358040
rect 519320 358028 519326 358080
rect 359550 356736 359556 356788
rect 359608 356776 359614 356788
rect 518986 356776 518992 356788
rect 359608 356748 518992 356776
rect 359608 356736 359614 356748
rect 518986 356736 518992 356748
rect 519044 356776 519050 356788
rect 519538 356776 519544 356788
rect 519044 356748 519544 356776
rect 519044 356736 519050 356748
rect 519538 356736 519544 356748
rect 519596 356736 519602 356788
rect 199654 356668 199660 356720
rect 199712 356708 199718 356720
rect 358998 356708 359004 356720
rect 199712 356680 359004 356708
rect 199712 356668 199718 356680
rect 358998 356668 359004 356680
rect 359056 356708 359062 356720
rect 359826 356708 359832 356720
rect 359056 356680 359832 356708
rect 359056 356668 359062 356680
rect 359826 356668 359832 356680
rect 359884 356668 359890 356720
rect 179322 351908 179328 351960
rect 179380 351948 179386 351960
rect 201494 351948 201500 351960
rect 179380 351920 201500 351948
rect 179380 351908 179386 351920
rect 201494 351908 201500 351920
rect 201552 351908 201558 351960
rect 203058 351908 203064 351960
rect 203116 351948 203122 351960
rect 206278 351948 206284 351960
rect 203116 351920 206284 351948
rect 203116 351908 203122 351920
rect 206278 351908 206284 351920
rect 206336 351908 206342 351960
rect 338482 351296 338488 351348
rect 338540 351336 338546 351348
rect 357066 351336 357072 351348
rect 338540 351308 357072 351336
rect 338540 351296 338546 351308
rect 357066 351296 357072 351308
rect 357124 351296 357130 351348
rect 361574 351336 361580 351348
rect 359292 351308 361580 351336
rect 340506 351228 340512 351280
rect 340564 351268 340570 351280
rect 359292 351268 359320 351308
rect 361574 351296 361580 351308
rect 361632 351296 361638 351348
rect 500586 351296 500592 351348
rect 500644 351336 500650 351348
rect 517698 351336 517704 351348
rect 500644 351308 517704 351336
rect 500644 351296 500650 351308
rect 517698 351296 517704 351308
rect 517756 351296 517762 351348
rect 340564 351240 359320 351268
rect 340564 351228 340570 351240
rect 360194 351228 360200 351280
rect 360252 351268 360258 351280
rect 360838 351268 360844 351280
rect 360252 351240 360844 351268
rect 360252 351228 360258 351240
rect 360838 351228 360844 351240
rect 360896 351228 360902 351280
rect 499022 351228 499028 351280
rect 499080 351268 499086 351280
rect 517790 351268 517796 351280
rect 499080 351240 517796 351268
rect 499080 351228 499086 351240
rect 517790 351228 517796 351240
rect 517848 351228 517854 351280
rect 191282 351160 191288 351212
rect 191340 351200 191346 351212
rect 202874 351200 202880 351212
rect 191340 351172 202880 351200
rect 191340 351160 191346 351172
rect 202874 351160 202880 351172
rect 202932 351200 202938 351212
rect 203058 351200 203064 351212
rect 202932 351172 203064 351200
rect 202932 351160 202938 351172
rect 203058 351160 203064 351172
rect 203116 351160 203122 351212
rect 351638 351160 351644 351212
rect 351696 351200 351702 351212
rect 360212 351200 360240 351228
rect 351696 351172 360240 351200
rect 351696 351160 351702 351172
rect 179690 350548 179696 350600
rect 179748 350588 179754 350600
rect 196618 350588 196624 350600
rect 179748 350560 196624 350588
rect 179748 350548 179754 350560
rect 196618 350548 196624 350560
rect 196676 350548 196682 350600
rect 510890 350548 510896 350600
rect 510948 350588 510954 350600
rect 511902 350588 511908 350600
rect 510948 350560 511908 350588
rect 510948 350548 510954 350560
rect 511902 350548 511908 350560
rect 511960 350588 511966 350600
rect 517514 350588 517520 350600
rect 511960 350560 517520 350588
rect 511960 350548 511966 350560
rect 517514 350548 517520 350560
rect 517572 350548 517578 350600
rect 219342 350480 219348 350532
rect 219400 350520 219406 350532
rect 220814 350520 220820 350532
rect 219400 350492 220820 350520
rect 219400 350480 219406 350492
rect 220814 350480 220820 350492
rect 220872 350480 220878 350532
rect 277302 349800 277308 349852
rect 277360 349840 277366 349852
rect 357526 349840 357532 349852
rect 277360 349812 357532 349840
rect 277360 349800 277366 349812
rect 357526 349800 357532 349812
rect 357584 349800 357590 349852
rect 502242 349800 502248 349852
rect 502300 349840 502306 349852
rect 517606 349840 517612 349852
rect 502300 349812 517612 349840
rect 502300 349800 502306 349812
rect 517606 349800 517612 349812
rect 517664 349800 517670 349852
rect 378594 349528 378600 349580
rect 378652 349568 378658 349580
rect 380894 349568 380900 349580
rect 378652 349540 380900 349568
rect 378652 349528 378658 349540
rect 380894 349528 380900 349540
rect 380952 349528 380958 349580
rect 216766 349188 216772 349240
rect 216824 349228 216830 349240
rect 220906 349228 220912 349240
rect 216824 349200 220912 349228
rect 216824 349188 216830 349200
rect 220906 349188 220912 349200
rect 220964 349188 220970 349240
rect 58618 349052 58624 349104
rect 58676 349092 58682 349104
rect 60734 349092 60740 349104
rect 58676 349064 60740 349092
rect 58676 349052 58682 349064
rect 60734 349052 60740 349064
rect 60792 349052 60798 349104
rect 58894 348644 58900 348696
rect 58952 348684 58958 348696
rect 62114 348684 62120 348696
rect 58952 348656 62120 348684
rect 58952 348644 58958 348656
rect 62114 348644 62120 348656
rect 62172 348644 62178 348696
rect 57146 346876 57152 346928
rect 57204 346916 57210 346928
rect 59354 346916 59360 346928
rect 57204 346888 59360 346916
rect 57204 346876 57210 346888
rect 59354 346876 59360 346888
rect 59412 346876 59418 346928
rect 540238 339396 540244 339448
rect 540296 339436 540302 339448
rect 580166 339436 580172 339448
rect 540296 339408 580172 339436
rect 540296 339396 540302 339408
rect 580166 339396 580172 339408
rect 580224 339396 580230 339448
rect 52914 320084 52920 320136
rect 52972 320124 52978 320136
rect 54294 320124 54300 320136
rect 52972 320096 54300 320124
rect 52972 320084 52978 320096
rect 54294 320084 54300 320096
rect 54352 320084 54358 320136
rect 48038 292476 48044 292528
rect 48096 292516 48102 292528
rect 57054 292516 57060 292528
rect 48096 292488 57060 292516
rect 48096 292476 48102 292488
rect 57054 292476 57060 292488
rect 57112 292516 57118 292528
rect 57330 292516 57336 292528
rect 57112 292488 57336 292516
rect 57112 292476 57118 292488
rect 57330 292476 57336 292488
rect 57388 292476 57394 292528
rect 57146 292204 57152 292256
rect 57204 292244 57210 292256
rect 59722 292244 59728 292256
rect 57204 292216 59728 292244
rect 57204 292204 57210 292216
rect 59722 292204 59728 292216
rect 59780 292204 59786 292256
rect 56870 291864 56876 291916
rect 56928 291904 56934 291916
rect 57974 291904 57980 291916
rect 56928 291876 57980 291904
rect 56928 291864 56934 291876
rect 57974 291864 57980 291876
rect 58032 291864 58038 291916
rect 376938 276224 376944 276276
rect 376996 276224 377002 276276
rect 376956 276072 376984 276224
rect 376938 276020 376944 276072
rect 376996 276020 377002 276072
rect 46290 275952 46296 276004
rect 46348 275992 46354 276004
rect 57606 275992 57612 276004
rect 46348 275964 57612 275992
rect 46348 275952 46354 275964
rect 57606 275952 57612 275964
rect 57664 275952 57670 276004
rect 203794 275952 203800 276004
rect 203852 275992 203858 276004
rect 216674 275992 216680 276004
rect 203852 275964 216680 275992
rect 203852 275952 203858 275964
rect 216674 275952 216680 275964
rect 216732 275952 216738 276004
rect 358078 275952 358084 276004
rect 358136 275992 358142 276004
rect 376846 275992 376852 276004
rect 358136 275964 376852 275992
rect 358136 275952 358142 275964
rect 376846 275952 376852 275964
rect 376904 275952 376910 276004
rect 202874 274592 202880 274644
rect 202932 274632 202938 274644
rect 216674 274632 216680 274644
rect 202932 274604 216680 274632
rect 202932 274592 202938 274604
rect 216674 274592 216680 274604
rect 216732 274592 216738 274644
rect 360194 274592 360200 274644
rect 360252 274632 360258 274644
rect 376754 274632 376760 274644
rect 360252 274604 376760 274632
rect 360252 274592 360258 274604
rect 376754 274592 376760 274604
rect 376812 274592 376818 274644
rect 197998 273912 198004 273964
rect 198056 273952 198062 273964
rect 202874 273952 202880 273964
rect 198056 273924 202880 273952
rect 198056 273912 198062 273924
rect 202874 273912 202880 273924
rect 202932 273912 202938 273964
rect 358078 273232 358084 273284
rect 358136 273272 358142 273284
rect 360194 273272 360200 273284
rect 358136 273244 360200 273272
rect 358136 273232 358142 273244
rect 360194 273232 360200 273244
rect 360252 273232 360258 273284
rect 206738 273164 206744 273216
rect 206796 273204 206802 273216
rect 216674 273204 216680 273216
rect 206796 273176 216680 273204
rect 206796 273164 206802 273176
rect 216674 273164 216680 273176
rect 216732 273164 216738 273216
rect 363966 273164 363972 273216
rect 364024 273204 364030 273216
rect 376754 273204 376760 273216
rect 364024 273176 376760 273204
rect 364024 273164 364030 273176
rect 376754 273164 376760 273176
rect 376812 273164 376818 273216
rect 376846 272484 376852 272536
rect 376904 272524 376910 272536
rect 377030 272524 377036 272536
rect 376904 272496 377036 272524
rect 376904 272484 376910 272496
rect 377030 272484 377036 272496
rect 377088 272484 377094 272536
rect 54294 271124 54300 271176
rect 54352 271164 54358 271176
rect 57974 271164 57980 271176
rect 54352 271136 57980 271164
rect 54352 271124 54358 271136
rect 57974 271124 57980 271136
rect 58032 271124 58038 271176
rect 214374 265344 214380 265396
rect 214432 265384 214438 265396
rect 215018 265384 215024 265396
rect 214432 265356 215024 265384
rect 214432 265344 214438 265356
rect 215018 265344 215024 265356
rect 215076 265344 215082 265396
rect 214650 265208 214656 265260
rect 214708 265248 214714 265260
rect 215018 265248 215024 265260
rect 214708 265220 215024 265248
rect 214708 265208 214714 265220
rect 215018 265208 215024 265220
rect 215076 265208 215082 265260
rect 48866 264936 48872 264988
rect 48924 264976 48930 264988
rect 58618 264976 58624 264988
rect 48924 264948 58624 264976
rect 48924 264936 48930 264948
rect 58618 264936 58624 264948
rect 58676 264936 58682 264988
rect 51534 264868 51540 264920
rect 51592 264908 51598 264920
rect 110966 264908 110972 264920
rect 51592 264880 110972 264908
rect 51592 264868 51598 264880
rect 110966 264868 110972 264880
rect 111024 264868 111030 264920
rect 219158 264868 219164 264920
rect 219216 264908 219222 264920
rect 221182 264908 221188 264920
rect 219216 264880 221188 264908
rect 219216 264868 219222 264880
rect 221182 264868 221188 264880
rect 221240 264868 221246 264920
rect 373626 264868 373632 264920
rect 373684 264908 373690 264920
rect 425974 264908 425980 264920
rect 373684 264880 425980 264908
rect 373684 264868 373690 264880
rect 425974 264868 425980 264880
rect 426032 264868 426038 264920
rect 42150 264800 42156 264852
rect 42208 264840 42214 264852
rect 125962 264840 125968 264852
rect 42208 264812 125968 264840
rect 42208 264800 42214 264812
rect 125962 264800 125968 264812
rect 126020 264800 126026 264852
rect 218606 264800 218612 264852
rect 218664 264840 218670 264852
rect 221090 264840 221096 264852
rect 218664 264812 221096 264840
rect 218664 264800 218670 264812
rect 221090 264800 221096 264812
rect 221148 264800 221154 264852
rect 368198 264800 368204 264852
rect 368256 264840 368262 264852
rect 421098 264840 421104 264852
rect 368256 264812 421104 264840
rect 368256 264800 368262 264812
rect 421098 264800 421104 264812
rect 421156 264800 421162 264852
rect 45002 264732 45008 264784
rect 45060 264772 45066 264784
rect 130930 264772 130936 264784
rect 45060 264744 130936 264772
rect 45060 264732 45066 264744
rect 130930 264732 130936 264744
rect 130988 264732 130994 264784
rect 208026 264732 208032 264784
rect 208084 264772 208090 264784
rect 214650 264772 214656 264784
rect 208084 264744 214656 264772
rect 208084 264732 208090 264744
rect 214650 264732 214656 264744
rect 214708 264732 214714 264784
rect 218514 264732 218520 264784
rect 218572 264772 218578 264784
rect 220998 264772 221004 264784
rect 218572 264744 221004 264772
rect 218572 264732 218578 264744
rect 220998 264732 221004 264744
rect 221056 264732 221062 264784
rect 373074 264732 373080 264784
rect 373132 264772 373138 264784
rect 374454 264772 374460 264784
rect 373132 264744 374460 264772
rect 373132 264732 373138 264744
rect 374454 264732 374460 264744
rect 374512 264772 374518 264784
rect 429746 264772 429752 264784
rect 374512 264744 429752 264772
rect 374512 264732 374518 264744
rect 429746 264732 429752 264744
rect 429804 264732 429810 264784
rect 43530 264664 43536 264716
rect 43588 264704 43594 264716
rect 128354 264704 128360 264716
rect 43588 264676 128360 264704
rect 43588 264664 43594 264676
rect 128354 264664 128360 264676
rect 128412 264664 128418 264716
rect 207842 264664 207848 264716
rect 207900 264704 207906 264716
rect 250438 264704 250444 264716
rect 207900 264676 250444 264704
rect 207900 264664 207906 264676
rect 250438 264664 250444 264676
rect 250496 264664 250502 264716
rect 362586 264664 362592 264716
rect 362644 264704 362650 264716
rect 418430 264704 418436 264716
rect 362644 264676 418436 264704
rect 362644 264664 362650 264676
rect 418430 264664 418436 264676
rect 418488 264664 418494 264716
rect 45186 264596 45192 264648
rect 45244 264636 45250 264648
rect 133414 264636 133420 264648
rect 45244 264608 133420 264636
rect 45244 264596 45250 264608
rect 133414 264596 133420 264608
rect 133472 264596 133478 264648
rect 217226 264596 217232 264648
rect 217284 264636 217290 264648
rect 220906 264636 220912 264648
rect 217284 264608 220912 264636
rect 217284 264596 217290 264608
rect 220906 264596 220912 264608
rect 220964 264596 220970 264648
rect 224218 264596 224224 264648
rect 224276 264636 224282 264648
rect 274174 264636 274180 264648
rect 224276 264608 274180 264636
rect 224276 264596 224282 264608
rect 274174 264596 274180 264608
rect 274232 264596 274238 264648
rect 365530 264596 365536 264648
rect 365588 264636 365594 264648
rect 468478 264636 468484 264648
rect 365588 264608 468484 264636
rect 365588 264596 365594 264608
rect 468478 264596 468484 264608
rect 468536 264596 468542 264648
rect 45094 264528 45100 264580
rect 45152 264568 45158 264580
rect 135898 264568 135904 264580
rect 45152 264540 135904 264568
rect 45152 264528 45158 264540
rect 135898 264528 135904 264540
rect 135956 264528 135962 264580
rect 214834 264528 214840 264580
rect 214892 264568 214898 264580
rect 280798 264568 280804 264580
rect 214892 264540 280804 264568
rect 214892 264528 214898 264540
rect 280798 264528 280804 264540
rect 280856 264528 280862 264580
rect 375006 264528 375012 264580
rect 375064 264568 375070 264580
rect 480898 264568 480904 264580
rect 375064 264540 480904 264568
rect 375064 264528 375070 264540
rect 480898 264528 480904 264540
rect 480956 264528 480962 264580
rect 46198 264460 46204 264512
rect 46256 264500 46262 264512
rect 138474 264500 138480 264512
rect 46256 264472 138480 264500
rect 46256 264460 46262 264472
rect 138474 264460 138480 264472
rect 138532 264460 138538 264512
rect 216214 264460 216220 264512
rect 216272 264500 216278 264512
rect 285950 264500 285956 264512
rect 216272 264472 285956 264500
rect 216272 264460 216278 264472
rect 285950 264460 285956 264472
rect 286008 264460 286014 264512
rect 366818 264460 366824 264512
rect 366876 264500 366882 264512
rect 473446 264500 473452 264512
rect 366876 264472 473452 264500
rect 366876 264460 366882 264472
rect 473446 264460 473452 264472
rect 473504 264460 473510 264512
rect 48130 264392 48136 264444
rect 48188 264432 48194 264444
rect 143534 264432 143540 264444
rect 48188 264404 143540 264432
rect 48188 264392 48194 264404
rect 143534 264392 143540 264404
rect 143592 264392 143598 264444
rect 210786 264392 210792 264444
rect 210844 264432 210850 264444
rect 283374 264432 283380 264444
rect 210844 264404 283380 264432
rect 210844 264392 210850 264404
rect 283374 264392 283380 264404
rect 283432 264392 283438 264444
rect 363874 264392 363880 264444
rect 363932 264432 363938 264444
rect 470962 264432 470968 264444
rect 363932 264404 470968 264432
rect 363932 264392 363938 264404
rect 470962 264392 470968 264404
rect 471020 264392 471026 264444
rect 43438 264324 43444 264376
rect 43496 264364 43502 264376
rect 140866 264364 140872 264376
rect 43496 264336 140872 264364
rect 43496 264324 43502 264336
rect 140866 264324 140872 264336
rect 140924 264324 140930 264376
rect 209406 264324 209412 264376
rect 209464 264364 209470 264376
rect 290918 264364 290924 264376
rect 209464 264336 290924 264364
rect 209464 264324 209470 264336
rect 290918 264324 290924 264336
rect 290976 264324 290982 264376
rect 372338 264324 372344 264376
rect 372396 264364 372402 264376
rect 483382 264364 483388 264376
rect 372396 264336 483388 264364
rect 372396 264324 372402 264336
rect 483382 264324 483388 264336
rect 483440 264324 483446 264376
rect 45278 264256 45284 264308
rect 45336 264296 45342 264308
rect 145926 264296 145932 264308
rect 45336 264268 145932 264296
rect 45336 264256 45342 264268
rect 145926 264256 145932 264268
rect 145984 264256 145990 264308
rect 203702 264256 203708 264308
rect 203760 264296 203766 264308
rect 288158 264296 288164 264308
rect 203760 264268 288164 264296
rect 203760 264256 203766 264268
rect 288158 264256 288164 264268
rect 288216 264256 288222 264308
rect 369486 264256 369492 264308
rect 369544 264296 369550 264308
rect 485958 264296 485964 264308
rect 369544 264268 485964 264296
rect 369544 264256 369550 264268
rect 485958 264256 485964 264268
rect 486016 264256 486022 264308
rect 45370 264188 45376 264240
rect 45428 264228 45434 264240
rect 148502 264228 148508 264240
rect 45428 264200 148508 264228
rect 45428 264188 45434 264200
rect 148502 264188 148508 264200
rect 148560 264188 148566 264240
rect 200942 264188 200948 264240
rect 201000 264228 201006 264240
rect 293402 264228 293408 264240
rect 201000 264200 293408 264228
rect 201000 264188 201006 264200
rect 293402 264188 293408 264200
rect 293460 264188 293466 264240
rect 356882 264188 356888 264240
rect 356940 264228 356946 264240
rect 475838 264228 475844 264240
rect 356940 264200 475844 264228
rect 356940 264188 356946 264200
rect 475838 264188 475844 264200
rect 475896 264188 475902 264240
rect 46382 264120 46388 264172
rect 46440 264160 46446 264172
rect 62206 264160 62212 264172
rect 46440 264132 62212 264160
rect 46440 264120 46446 264132
rect 62206 264120 62212 264132
rect 62264 264120 62270 264172
rect 212994 264120 213000 264172
rect 213052 264160 213058 264172
rect 224218 264160 224224 264172
rect 213052 264132 224224 264160
rect 213052 264120 213058 264132
rect 224218 264120 224224 264132
rect 224276 264120 224282 264172
rect 370958 264120 370964 264172
rect 371016 264160 371022 264172
rect 423490 264160 423496 264172
rect 371016 264132 423496 264160
rect 371016 264120 371022 264132
rect 423490 264120 423496 264132
rect 423548 264120 423554 264172
rect 46474 264052 46480 264104
rect 46532 264092 46538 264104
rect 62114 264092 62120 264104
rect 46532 264064 62120 264092
rect 46532 264052 46538 264064
rect 62114 264052 62120 264064
rect 62172 264052 62178 264104
rect 214650 264052 214656 264104
rect 214708 264092 214714 264104
rect 220814 264092 220820 264104
rect 214708 264064 220820 264092
rect 214708 264052 214714 264064
rect 220814 264052 220820 264064
rect 220872 264052 220878 264104
rect 62206 263712 62212 263764
rect 62264 263752 62270 263764
rect 89990 263752 89996 263764
rect 62264 263724 89996 263752
rect 62264 263712 62270 263724
rect 89990 263712 89996 263724
rect 90048 263712 90054 263764
rect 58894 263644 58900 263696
rect 58952 263684 58958 263696
rect 62298 263684 62304 263696
rect 58952 263656 62304 263684
rect 58952 263644 58958 263656
rect 62298 263644 62304 263656
rect 62356 263684 62362 263696
rect 92382 263684 92388 263696
rect 62356 263656 92388 263684
rect 62356 263644 62362 263656
rect 92382 263644 92388 263656
rect 92440 263644 92446 263696
rect 211614 263644 211620 263696
rect 211672 263684 211678 263696
rect 214282 263684 214288 263696
rect 211672 263656 214288 263684
rect 211672 263644 211678 263656
rect 214282 263644 214288 263656
rect 214340 263684 214346 263696
rect 214340 263656 219434 263684
rect 214340 263644 214346 263656
rect 62114 263576 62120 263628
rect 62172 263616 62178 263628
rect 91278 263616 91284 263628
rect 62172 263588 91284 263616
rect 62172 263576 62178 263588
rect 91278 263576 91284 263588
rect 91336 263576 91342 263628
rect 212350 263576 212356 263628
rect 212408 263616 212414 263628
rect 212994 263616 213000 263628
rect 212408 263588 213000 263616
rect 212408 263576 212414 263588
rect 212994 263576 213000 263588
rect 213052 263576 213058 263628
rect 219406 263616 219434 263656
rect 373902 263644 373908 263696
rect 373960 263684 373966 263696
rect 374362 263684 374368 263696
rect 373960 263656 374368 263684
rect 373960 263644 373966 263656
rect 374362 263644 374368 263656
rect 374420 263684 374426 263696
rect 433334 263684 433340 263696
rect 374420 263656 433340 263684
rect 374420 263644 374426 263656
rect 433334 263644 433340 263656
rect 433392 263644 433398 263696
rect 273254 263616 273260 263628
rect 219406 263588 273260 263616
rect 273254 263576 273260 263588
rect 273312 263576 273318 263628
rect 279234 263576 279240 263628
rect 279292 263616 279298 263628
rect 357710 263616 357716 263628
rect 279292 263588 357716 263616
rect 279292 263576 279298 263588
rect 357710 263576 357716 263588
rect 357768 263616 357774 263628
rect 359274 263616 359280 263628
rect 357768 263588 359280 263616
rect 357768 263576 357774 263588
rect 359274 263576 359280 263588
rect 359332 263576 359338 263628
rect 371786 263576 371792 263628
rect 371844 263616 371850 263628
rect 373626 263616 373632 263628
rect 371844 263588 373632 263616
rect 371844 263576 371850 263588
rect 373626 263576 373632 263588
rect 373684 263616 373690 263628
rect 432230 263616 432236 263628
rect 373684 263588 432236 263616
rect 373684 263576 373690 263588
rect 432230 263576 432236 263588
rect 432288 263576 432294 263628
rect 54478 263508 54484 263560
rect 54536 263548 54542 263560
rect 120902 263548 120908 263560
rect 54536 263520 120908 263548
rect 54536 263508 54542 263520
rect 120902 263508 120908 263520
rect 120960 263508 120966 263560
rect 155954 263508 155960 263560
rect 156012 263548 156018 263560
rect 204346 263548 204352 263560
rect 156012 263520 204352 263548
rect 156012 263508 156018 263520
rect 204346 263508 204352 263520
rect 204404 263508 204410 263560
rect 210694 263508 210700 263560
rect 210752 263548 210758 263560
rect 308398 263548 308404 263560
rect 210752 263520 308404 263548
rect 210752 263508 210758 263520
rect 308398 263508 308404 263520
rect 308456 263508 308462 263560
rect 362494 263508 362500 263560
rect 362552 263548 362558 263560
rect 453390 263548 453396 263560
rect 362552 263520 453396 263548
rect 362552 263508 362558 263520
rect 453390 263508 453396 263520
rect 453448 263508 453454 263560
rect 57790 263440 57796 263492
rect 57848 263480 57854 263492
rect 123478 263480 123484 263492
rect 57848 263452 123484 263480
rect 57848 263440 57854 263452
rect 123478 263440 123484 263452
rect 123536 263440 123542 263492
rect 158530 263440 158536 263492
rect 158588 263480 158594 263492
rect 205634 263480 205640 263492
rect 158588 263452 205640 263480
rect 158588 263440 158594 263452
rect 205634 263440 205640 263452
rect 205692 263440 205698 263492
rect 212258 263440 212264 263492
rect 212316 263480 212322 263492
rect 305822 263480 305828 263492
rect 212316 263452 305828 263480
rect 212316 263440 212322 263452
rect 305822 263440 305828 263452
rect 305880 263440 305886 263492
rect 368106 263440 368112 263492
rect 368164 263480 368170 263492
rect 455782 263480 455788 263492
rect 368164 263452 455788 263480
rect 368164 263440 368170 263452
rect 455782 263440 455788 263452
rect 455840 263440 455846 263492
rect 53098 263372 53104 263424
rect 53156 263412 53162 263424
rect 115934 263412 115940 263424
rect 53156 263384 115940 263412
rect 53156 263372 53162 263384
rect 115934 263372 115940 263384
rect 115992 263372 115998 263424
rect 150986 263372 150992 263424
rect 151044 263412 151050 263424
rect 197630 263412 197636 263424
rect 151044 263384 197636 263412
rect 151044 263372 151050 263384
rect 197630 263372 197636 263384
rect 197688 263372 197694 263424
rect 205082 263372 205088 263424
rect 205140 263412 205146 263424
rect 268286 263412 268292 263424
rect 205140 263384 268292 263412
rect 205140 263372 205146 263384
rect 268286 263372 268292 263384
rect 268344 263372 268350 263424
rect 370866 263372 370872 263424
rect 370924 263412 370930 263424
rect 450998 263412 451004 263424
rect 370924 263384 451004 263412
rect 370924 263372 370930 263384
rect 450998 263372 451004 263384
rect 451056 263372 451062 263424
rect 54570 263304 54576 263356
rect 54628 263344 54634 263356
rect 118050 263344 118056 263356
rect 54628 263316 118056 263344
rect 54628 263304 54634 263316
rect 118050 263304 118056 263316
rect 118108 263304 118114 263356
rect 161106 263304 161112 263356
rect 161164 263344 161170 263356
rect 207106 263344 207112 263356
rect 161164 263316 207112 263344
rect 161164 263304 161170 263316
rect 207106 263304 207112 263316
rect 207164 263304 207170 263356
rect 214742 263304 214748 263356
rect 214800 263344 214806 263356
rect 276106 263344 276112 263356
rect 214800 263316 276112 263344
rect 214800 263304 214806 263316
rect 276106 263304 276112 263316
rect 276164 263304 276170 263356
rect 364058 263304 364064 263356
rect 364116 263344 364122 263356
rect 443454 263344 443460 263356
rect 364116 263316 443460 263344
rect 364116 263304 364122 263316
rect 443454 263304 443460 263316
rect 443512 263304 443518 263356
rect 53006 263236 53012 263288
rect 53064 263276 53070 263288
rect 113358 263276 113364 263288
rect 53064 263248 113364 263276
rect 53064 263236 53070 263248
rect 113358 263236 113364 263248
rect 113416 263236 113422 263288
rect 166074 263236 166080 263288
rect 166132 263276 166138 263288
rect 210050 263276 210056 263288
rect 166132 263248 210056 263276
rect 166132 263236 166138 263248
rect 210050 263236 210056 263248
rect 210108 263236 210114 263288
rect 210602 263236 210608 263288
rect 210660 263276 210666 263288
rect 270862 263276 270868 263288
rect 210660 263248 270868 263276
rect 210660 263236 210666 263248
rect 270862 263236 270868 263248
rect 270920 263236 270926 263288
rect 361298 263236 361304 263288
rect 361356 263276 361362 263288
rect 438394 263276 438400 263288
rect 361356 263248 438400 263276
rect 361356 263236 361362 263248
rect 438394 263236 438400 263248
rect 438452 263236 438458 263288
rect 53374 263168 53380 263220
rect 53432 263208 53438 263220
rect 108206 263208 108212 263220
rect 53432 263180 108212 263208
rect 53432 263168 53438 263180
rect 108206 263168 108212 263180
rect 108264 263168 108270 263220
rect 163498 263168 163504 263220
rect 163556 263208 163562 263220
rect 197722 263208 197728 263220
rect 163556 263180 197728 263208
rect 163556 263168 163562 263180
rect 197722 263168 197728 263180
rect 197780 263168 197786 263220
rect 209314 263168 209320 263220
rect 209372 263208 209378 263220
rect 265894 263208 265900 263220
rect 209372 263180 265900 263208
rect 209372 263168 209378 263180
rect 265894 263168 265900 263180
rect 265952 263168 265958 263220
rect 372246 263168 372252 263220
rect 372304 263208 372310 263220
rect 448238 263208 448244 263220
rect 372304 263180 448244 263208
rect 372304 263168 372310 263180
rect 448238 263168 448244 263180
rect 448296 263168 448302 263220
rect 51626 263100 51632 263152
rect 51684 263140 51690 263152
rect 105630 263140 105636 263152
rect 51684 263112 105636 263140
rect 51684 263100 51690 263112
rect 105630 263100 105636 263112
rect 105688 263100 105694 263152
rect 200850 263100 200856 263152
rect 200908 263140 200914 263152
rect 256142 263140 256148 263152
rect 200908 263112 256148 263140
rect 200908 263100 200914 263112
rect 256142 263100 256148 263112
rect 256200 263100 256206 263152
rect 365346 263100 365352 263152
rect 365404 263140 365410 263152
rect 435910 263140 435916 263152
rect 365404 263112 435916 263140
rect 365404 263100 365410 263112
rect 435910 263100 435916 263112
rect 435968 263100 435974 263152
rect 51810 263032 51816 263084
rect 51868 263072 51874 263084
rect 103514 263072 103520 263084
rect 51868 263044 103520 263072
rect 51868 263032 51874 263044
rect 103514 263032 103520 263044
rect 103572 263032 103578 263084
rect 206554 263032 206560 263084
rect 206612 263072 206618 263084
rect 260926 263072 260932 263084
rect 206612 263044 260932 263072
rect 206612 263032 206618 263044
rect 260926 263032 260932 263044
rect 260984 263032 260990 263084
rect 373534 263032 373540 263084
rect 373592 263072 373598 263084
rect 440878 263072 440884 263084
rect 373592 263044 440884 263072
rect 373592 263032 373598 263044
rect 440878 263032 440884 263044
rect 440936 263032 440942 263084
rect 503530 263032 503536 263084
rect 503588 263072 503594 263084
rect 517606 263072 517612 263084
rect 503588 263044 517612 263072
rect 503588 263032 503594 263044
rect 517606 263032 517612 263044
rect 517664 263032 517670 263084
rect 50246 262964 50252 263016
rect 50304 263004 50310 263016
rect 101030 263004 101036 263016
rect 50304 262976 101036 263004
rect 50304 262964 50310 262976
rect 101030 262964 101036 262976
rect 101088 262964 101094 263016
rect 183370 262964 183376 263016
rect 183428 263004 183434 263016
rect 201586 263004 201592 263016
rect 183428 262976 201592 263004
rect 183428 262964 183434 262976
rect 201586 262964 201592 262976
rect 201644 262964 201650 263016
rect 218974 262964 218980 263016
rect 219032 263004 219038 263016
rect 273346 263004 273352 263016
rect 219032 262976 273352 263004
rect 219032 262964 219038 262976
rect 273346 262964 273352 262976
rect 273404 262964 273410 263016
rect 343542 262964 343548 263016
rect 343600 263004 343606 263016
rect 357434 263004 357440 263016
rect 343600 262976 357440 263004
rect 343600 262964 343606 262976
rect 357434 262964 357440 262976
rect 357492 262964 357498 263016
rect 369302 262964 369308 263016
rect 369360 263004 369366 263016
rect 433518 263004 433524 263016
rect 369360 262976 433524 263004
rect 369360 262964 369366 262976
rect 433518 262964 433524 262976
rect 433576 262964 433582 263016
rect 50338 262896 50344 262948
rect 50396 262936 50402 262948
rect 98086 262936 98092 262948
rect 50396 262908 98092 262936
rect 50396 262896 50402 262908
rect 98086 262896 98092 262908
rect 98144 262896 98150 262948
rect 183462 262896 183468 262948
rect 183520 262936 183526 262948
rect 202966 262936 202972 262948
rect 183520 262908 202972 262936
rect 183520 262896 183526 262908
rect 202966 262896 202972 262908
rect 203024 262896 203030 262948
rect 212166 262896 212172 262948
rect 212224 262936 212230 262948
rect 263594 262936 263600 262948
rect 212224 262908 263600 262936
rect 212224 262896 212230 262908
rect 263594 262896 263600 262908
rect 263652 262896 263658 262948
rect 369394 262896 369400 262948
rect 369452 262936 369458 262948
rect 410702 262936 410708 262948
rect 369452 262908 410708 262936
rect 369452 262896 369458 262908
rect 410702 262896 410708 262908
rect 410760 262896 410766 262948
rect 503622 262896 503628 262948
rect 503680 262936 503686 262948
rect 517882 262936 517888 262948
rect 503680 262908 517888 262936
rect 503680 262896 503686 262908
rect 517882 262896 517888 262908
rect 517940 262896 517946 262948
rect 50430 262828 50436 262880
rect 50488 262868 50494 262880
rect 96062 262868 96068 262880
rect 50488 262840 96068 262868
rect 50488 262828 50494 262840
rect 96062 262828 96068 262840
rect 96120 262828 96126 262880
rect 114370 262828 114376 262880
rect 114428 262868 114434 262880
rect 196894 262868 196900 262880
rect 114428 262840 196900 262868
rect 114428 262828 114434 262840
rect 196894 262828 196900 262840
rect 196952 262828 196958 262880
rect 202230 262828 202236 262880
rect 202288 262868 202294 262880
rect 253566 262868 253572 262880
rect 202288 262840 253572 262868
rect 202288 262828 202294 262840
rect 253566 262828 253572 262840
rect 253624 262828 253630 262880
rect 343450 262828 343456 262880
rect 343508 262868 343514 262880
rect 360286 262868 360292 262880
rect 343508 262840 360292 262868
rect 343508 262828 343514 262840
rect 360286 262828 360292 262840
rect 360344 262828 360350 262880
rect 374822 262828 374828 262880
rect 374880 262868 374886 262880
rect 413646 262868 413652 262880
rect 374880 262840 413652 262868
rect 374880 262828 374886 262840
rect 413646 262828 413652 262840
rect 413704 262828 413710 262880
rect 49142 262760 49148 262812
rect 49200 262800 49206 262812
rect 93578 262800 93584 262812
rect 49200 262772 93584 262800
rect 49200 262760 49206 262772
rect 93578 262760 93584 262772
rect 93636 262760 93642 262812
rect 207934 262760 207940 262812
rect 207992 262800 207998 262812
rect 258350 262800 258356 262812
rect 207992 262772 258356 262800
rect 207992 262760 207998 262772
rect 258350 262760 258356 262772
rect 258408 262760 258414 262812
rect 379054 262760 379060 262812
rect 379112 262800 379118 262812
rect 415762 262800 415768 262812
rect 379112 262772 415768 262800
rect 379112 262760 379118 262772
rect 415762 262760 415768 262772
rect 415820 262760 415826 262812
rect 55766 262692 55772 262744
rect 55824 262732 55830 262744
rect 90726 262732 90732 262744
rect 55824 262704 90732 262732
rect 55824 262692 55830 262704
rect 90726 262692 90732 262704
rect 90784 262692 90790 262744
rect 215018 262692 215024 262744
rect 215076 262732 215082 262744
rect 247678 262732 247684 262744
rect 215076 262704 247684 262732
rect 215076 262692 215082 262704
rect 247678 262692 247684 262704
rect 247736 262692 247742 262744
rect 374914 262692 374920 262744
rect 374972 262732 374978 262744
rect 408310 262732 408316 262744
rect 374972 262704 408316 262732
rect 374972 262692 374978 262704
rect 408310 262692 408316 262704
rect 408368 262692 408374 262744
rect 54662 262624 54668 262676
rect 54720 262664 54726 262676
rect 88334 262664 88340 262676
rect 54720 262636 88340 262664
rect 54720 262624 54726 262636
rect 88334 262624 88340 262636
rect 88392 262624 88398 262676
rect 96522 262624 96528 262676
rect 96580 262664 96586 262676
rect 101766 262664 101772 262676
rect 96580 262636 101772 262664
rect 96580 262624 96586 262636
rect 101766 262624 101772 262636
rect 101824 262624 101830 262676
rect 210326 262624 210332 262676
rect 210384 262664 210390 262676
rect 213270 262664 213276 262676
rect 210384 262636 213276 262664
rect 210384 262624 210390 262636
rect 213270 262624 213276 262636
rect 213328 262624 213334 262676
rect 100018 262420 100024 262472
rect 100076 262460 100082 262472
rect 116210 262460 116216 262472
rect 100076 262432 116216 262460
rect 100076 262420 100082 262432
rect 116210 262420 116216 262432
rect 116268 262420 116274 262472
rect 511902 262420 511908 262472
rect 511960 262460 511966 262472
rect 517514 262460 517520 262472
rect 511960 262432 517520 262460
rect 511960 262420 511966 262432
rect 517514 262420 517520 262432
rect 517572 262420 517578 262472
rect 89714 262352 89720 262404
rect 89772 262392 89778 262404
rect 109310 262392 109316 262404
rect 89772 262364 109316 262392
rect 89772 262352 89778 262364
rect 109310 262352 109316 262364
rect 109368 262352 109374 262404
rect 213270 262216 213276 262268
rect 213328 262256 213334 262268
rect 272058 262256 272064 262268
rect 213328 262228 272064 262256
rect 213328 262216 213334 262228
rect 272058 262216 272064 262228
rect 272116 262216 272122 262268
rect 378686 262216 378692 262268
rect 378744 262256 378750 262268
rect 379974 262256 379980 262268
rect 378744 262228 379980 262256
rect 378744 262216 378750 262228
rect 379974 262216 379980 262228
rect 380032 262256 380038 262268
rect 415854 262256 415860 262268
rect 380032 262228 415860 262256
rect 380032 262216 380038 262228
rect 415854 262216 415860 262228
rect 415912 262216 415918 262268
rect 425698 262216 425704 262268
rect 425756 262256 425762 262268
rect 428274 262256 428280 262268
rect 425756 262228 428280 262256
rect 425756 262216 425762 262228
rect 428274 262216 428280 262228
rect 428332 262216 428338 262268
rect 206646 262148 206652 262200
rect 206704 262188 206710 262200
rect 325786 262188 325792 262200
rect 206704 262160 325792 262188
rect 206704 262148 206710 262160
rect 325786 262148 325792 262160
rect 325844 262148 325850 262200
rect 365438 262148 365444 262200
rect 365496 262188 365502 262200
rect 430942 262188 430948 262200
rect 365496 262160 430948 262188
rect 365496 262148 365502 262160
rect 430942 262148 430948 262160
rect 431000 262148 431006 262200
rect 205174 262080 205180 262132
rect 205232 262120 205238 262132
rect 323026 262120 323032 262132
rect 205232 262092 323032 262120
rect 205232 262080 205238 262092
rect 323026 262080 323032 262092
rect 323084 262080 323090 262132
rect 374914 262080 374920 262132
rect 374972 262120 374978 262132
rect 375834 262120 375840 262132
rect 374972 262092 375840 262120
rect 374972 262080 374978 262092
rect 375834 262080 375840 262092
rect 375892 262080 375898 262132
rect 376294 262080 376300 262132
rect 376352 262120 376358 262132
rect 428182 262120 428188 262132
rect 376352 262092 428188 262120
rect 376352 262080 376358 262092
rect 428182 262080 428188 262092
rect 428240 262080 428246 262132
rect 211706 262012 211712 262064
rect 211764 262052 211770 262064
rect 212902 262052 212908 262064
rect 211764 262024 212908 262052
rect 211764 262012 211770 262024
rect 212902 262012 212908 262024
rect 212960 262012 212966 262064
rect 373166 262012 373172 262064
rect 373224 262052 373230 262064
rect 376386 262052 376392 262064
rect 373224 262024 376392 262052
rect 373224 262012 373230 262024
rect 376386 262012 376392 262024
rect 376444 262012 376450 262064
rect 378594 262012 378600 262064
rect 378652 262052 378658 262064
rect 379238 262052 379244 262064
rect 378652 262024 379244 262052
rect 378652 262012 378658 262024
rect 379238 262012 379244 262024
rect 379296 262052 379302 262064
rect 426434 262052 426440 262064
rect 379296 262024 426440 262052
rect 379296 262012 379302 262024
rect 426434 262012 426440 262024
rect 426492 262012 426498 262064
rect 372982 261944 372988 261996
rect 373040 261984 373046 261996
rect 376294 261984 376300 261996
rect 373040 261956 376300 261984
rect 373040 261944 373046 261956
rect 376294 261944 376300 261956
rect 376352 261944 376358 261996
rect 379606 261944 379612 261996
rect 379664 261984 379670 261996
rect 396166 261984 396172 261996
rect 379664 261956 396172 261984
rect 379664 261944 379670 261956
rect 396166 261944 396172 261956
rect 396224 261944 396230 261996
rect 212902 261536 212908 261588
rect 212960 261576 212966 261588
rect 269758 261576 269764 261588
rect 212960 261548 269764 261576
rect 212960 261536 212966 261548
rect 269758 261536 269764 261548
rect 269816 261536 269822 261588
rect 375834 261536 375840 261588
rect 375892 261576 375898 261588
rect 393406 261576 393412 261588
rect 375892 261548 393412 261576
rect 375892 261536 375898 261548
rect 393406 261536 393412 261548
rect 393464 261536 393470 261588
rect 208946 261468 208952 261520
rect 209004 261508 209010 261520
rect 212810 261508 212816 261520
rect 209004 261480 212816 261508
rect 209004 261468 209010 261480
rect 212810 261468 212816 261480
rect 212868 261508 212874 261520
rect 271230 261508 271236 261520
rect 212868 261480 271236 261508
rect 212868 261468 212874 261480
rect 271230 261468 271236 261480
rect 271288 261468 271294 261520
rect 380342 261468 380348 261520
rect 380400 261508 380406 261520
rect 425238 261508 425244 261520
rect 380400 261480 425244 261508
rect 380400 261468 380406 261480
rect 425238 261468 425244 261480
rect 425296 261468 425302 261520
rect 379330 260992 379336 261044
rect 379388 261032 379394 261044
rect 389174 261032 389180 261044
rect 379388 261004 389180 261032
rect 379388 260992 379394 261004
rect 389174 260992 389180 261004
rect 389232 260992 389238 261044
rect 376294 260924 376300 260976
rect 376352 260964 376358 260976
rect 388438 260964 388444 260976
rect 376352 260936 388444 260964
rect 376352 260924 376358 260936
rect 388438 260924 388444 260936
rect 388496 260924 388502 260976
rect 52822 260856 52828 260908
rect 52880 260896 52886 260908
rect 57974 260896 57980 260908
rect 52880 260868 57980 260896
rect 52880 260856 52886 260868
rect 57974 260856 57980 260868
rect 58032 260896 58038 260908
rect 58032 260868 59308 260896
rect 58032 260856 58038 260868
rect 59280 260760 59308 260868
rect 214300 260868 214972 260896
rect 59722 260788 59728 260840
rect 59780 260828 59786 260840
rect 118694 260828 118700 260840
rect 59780 260800 118700 260828
rect 59780 260788 59786 260800
rect 118694 260788 118700 260800
rect 118752 260788 118758 260840
rect 213546 260788 213552 260840
rect 213604 260828 213610 260840
rect 214300 260828 214328 260868
rect 213604 260800 214328 260828
rect 213604 260788 213610 260800
rect 214374 260788 214380 260840
rect 214432 260828 214438 260840
rect 214834 260828 214840 260840
rect 214432 260800 214840 260828
rect 214432 260788 214438 260800
rect 214834 260788 214840 260800
rect 214892 260788 214898 260840
rect 214944 260828 214972 260868
rect 376386 260856 376392 260908
rect 376444 260896 376450 260908
rect 390554 260896 390560 260908
rect 376444 260868 390560 260896
rect 376444 260856 376450 260868
rect 390554 260856 390560 260868
rect 390612 260856 390618 260908
rect 244366 260828 244372 260840
rect 214944 260800 244372 260828
rect 244366 260788 244372 260800
rect 244424 260788 244430 260840
rect 375006 260788 375012 260840
rect 375064 260828 375070 260840
rect 375190 260828 375196 260840
rect 375064 260800 375196 260828
rect 375064 260788 375070 260800
rect 375190 260788 375196 260800
rect 375248 260788 375254 260840
rect 375926 260788 375932 260840
rect 375984 260828 375990 260840
rect 377030 260828 377036 260840
rect 375984 260800 377036 260828
rect 375984 260788 375990 260800
rect 377030 260788 377036 260800
rect 377088 260788 377094 260840
rect 435174 260828 435180 260840
rect 383626 260800 435180 260828
rect 100754 260760 100760 260772
rect 59280 260732 100760 260760
rect 100754 260720 100760 260732
rect 100812 260720 100818 260772
rect 213086 260720 213092 260772
rect 213144 260760 213150 260772
rect 214742 260760 214748 260772
rect 213144 260732 214748 260760
rect 213144 260720 213150 260732
rect 214742 260720 214748 260732
rect 214800 260720 214806 260772
rect 214852 260760 214880 260788
rect 243078 260760 243084 260772
rect 214852 260732 243084 260760
rect 243078 260720 243084 260732
rect 243136 260720 243142 260772
rect 375208 260760 375236 260788
rect 383626 260760 383654 260800
rect 435174 260788 435180 260800
rect 435232 260788 435238 260840
rect 375208 260732 383654 260760
rect 388438 260720 388444 260772
rect 388496 260760 388502 260772
rect 421742 260760 421748 260772
rect 388496 260732 421748 260760
rect 388496 260720 388502 260732
rect 421742 260720 421748 260732
rect 421800 260720 421806 260772
rect 50522 260652 50528 260704
rect 50580 260692 50586 260704
rect 84194 260692 84200 260704
rect 50580 260664 84200 260692
rect 50580 260652 50586 260664
rect 84194 260652 84200 260664
rect 84252 260652 84258 260704
rect 389174 260652 389180 260704
rect 389232 260692 389238 260704
rect 419810 260692 419816 260704
rect 389232 260664 419816 260692
rect 389232 260652 389238 260664
rect 419810 260652 419816 260664
rect 419868 260652 419874 260704
rect 51718 260584 51724 260636
rect 51776 260624 51782 260636
rect 84746 260624 84752 260636
rect 51776 260596 84752 260624
rect 51776 260584 51782 260596
rect 84746 260584 84752 260596
rect 84804 260584 84810 260636
rect 390554 260584 390560 260636
rect 390612 260624 390618 260636
rect 419350 260624 419356 260636
rect 390612 260596 419356 260624
rect 390612 260584 390618 260596
rect 419350 260584 419356 260596
rect 419408 260584 419414 260636
rect 53190 260516 53196 260568
rect 53248 260556 53254 260568
rect 54570 260556 54576 260568
rect 53248 260528 54576 260556
rect 53248 260516 53254 260528
rect 54570 260516 54576 260528
rect 54628 260556 54634 260568
rect 87598 260556 87604 260568
rect 54628 260528 87604 260556
rect 54628 260516 54634 260528
rect 87598 260516 87604 260528
rect 87656 260516 87662 260568
rect 393406 260516 393412 260568
rect 393464 260556 393470 260568
rect 418154 260556 418160 260568
rect 393464 260528 418160 260556
rect 393464 260516 393470 260528
rect 418154 260516 418160 260528
rect 418212 260516 418218 260568
rect 55766 260448 55772 260500
rect 55824 260488 55830 260500
rect 88610 260488 88616 260500
rect 55824 260460 88616 260488
rect 55824 260448 55830 260460
rect 88610 260448 88616 260460
rect 88668 260448 88674 260500
rect 49050 260380 49056 260432
rect 49108 260420 49114 260432
rect 89714 260420 89720 260432
rect 49108 260392 89720 260420
rect 49108 260380 49114 260392
rect 89714 260380 89720 260392
rect 89772 260380 89778 260432
rect 57974 260312 57980 260364
rect 58032 260352 58038 260364
rect 102318 260352 102324 260364
rect 58032 260324 102324 260352
rect 58032 260312 58038 260324
rect 102318 260312 102324 260324
rect 102376 260312 102382 260364
rect 52914 260244 52920 260296
rect 52972 260284 52978 260296
rect 54294 260284 54300 260296
rect 52972 260256 54300 260284
rect 52972 260244 52978 260256
rect 54294 260244 54300 260256
rect 54352 260284 54358 260296
rect 99466 260284 99472 260296
rect 54352 260256 99472 260284
rect 54352 260244 54358 260256
rect 99466 260244 99472 260256
rect 99524 260244 99530 260296
rect 45462 260176 45468 260228
rect 45520 260216 45526 260228
rect 49050 260216 49056 260228
rect 45520 260188 49056 260216
rect 45520 260176 45526 260188
rect 49050 260176 49056 260188
rect 49108 260176 49114 260228
rect 51626 260176 51632 260228
rect 51684 260216 51690 260228
rect 105078 260216 105084 260228
rect 51684 260188 105084 260216
rect 51684 260176 51690 260188
rect 105078 260176 105084 260188
rect 105136 260176 105142 260228
rect 377030 260176 377036 260228
rect 377088 260216 377094 260228
rect 423950 260216 423956 260228
rect 377088 260188 423956 260216
rect 377088 260176 377094 260188
rect 423950 260176 423956 260188
rect 424008 260176 424014 260228
rect 42242 260108 42248 260160
rect 42300 260148 42306 260160
rect 46198 260148 46204 260160
rect 42300 260120 46204 260148
rect 42300 260108 42306 260120
rect 46198 260108 46204 260120
rect 46256 260148 46262 260160
rect 108022 260148 108028 260160
rect 46256 260120 108028 260148
rect 46256 260108 46262 260120
rect 108022 260108 108028 260120
rect 108080 260108 108086 260160
rect 214742 260108 214748 260160
rect 214800 260148 214806 260160
rect 235994 260148 236000 260160
rect 214800 260120 236000 260148
rect 214800 260108 214806 260120
rect 235994 260108 236000 260120
rect 236052 260108 236058 260160
rect 379606 260108 379612 260160
rect 379664 260148 379670 260160
rect 427446 260148 427452 260160
rect 379664 260120 427452 260148
rect 379664 260108 379670 260120
rect 427446 260108 427452 260120
rect 427504 260108 427510 260160
rect 53282 260040 53288 260092
rect 53340 260080 53346 260092
rect 85942 260080 85948 260092
rect 53340 260052 85948 260080
rect 53340 260040 53346 260052
rect 85942 260040 85948 260052
rect 86000 260040 86006 260092
rect 54386 259972 54392 260024
rect 54444 260012 54450 260024
rect 64874 260012 64880 260024
rect 54444 259984 64880 260012
rect 54444 259972 54450 259984
rect 64874 259972 64880 259984
rect 64932 259972 64938 260024
rect 43714 259360 43720 259412
rect 43772 259400 43778 259412
rect 57974 259400 57980 259412
rect 43772 259372 57980 259400
rect 43772 259360 43778 259372
rect 57974 259360 57980 259372
rect 58032 259360 58038 259412
rect 46658 259292 46664 259344
rect 46716 259332 46722 259344
rect 55766 259332 55772 259344
rect 46716 259304 55772 259332
rect 46716 259292 46722 259304
rect 55766 259292 55772 259304
rect 55824 259292 55830 259344
rect 43622 259224 43628 259276
rect 43680 259264 43686 259276
rect 51626 259264 51632 259276
rect 43680 259236 51632 259264
rect 43680 259224 43686 259236
rect 51626 259224 51632 259236
rect 51684 259224 51690 259276
rect 372430 244196 372436 244248
rect 372488 244236 372494 244248
rect 374546 244236 374552 244248
rect 372488 244208 374552 244236
rect 372488 244196 372494 244208
rect 374546 244196 374552 244208
rect 374604 244196 374610 244248
rect 440142 244196 440148 244248
rect 440200 244236 440206 244248
rect 516686 244236 516692 244248
rect 440200 244208 516692 244236
rect 440200 244196 440206 244208
rect 516686 244196 516692 244208
rect 516744 244196 516750 244248
rect 371050 243652 371056 243704
rect 371108 243692 371114 243704
rect 373534 243692 373540 243704
rect 371108 243664 373540 243692
rect 371108 243652 371114 243664
rect 373534 243652 373540 243664
rect 373592 243692 373598 243704
rect 398834 243692 398840 243704
rect 373592 243664 398840 243692
rect 373592 243652 373598 243664
rect 398834 243652 398840 243664
rect 398892 243652 398898 243704
rect 374546 243584 374552 243636
rect 374604 243624 374610 243636
rect 374822 243624 374828 243636
rect 374604 243596 374828 243624
rect 374604 243584 374610 243596
rect 374822 243584 374828 243596
rect 374880 243624 374886 243636
rect 401594 243624 401600 243636
rect 374880 243596 401600 243624
rect 374880 243584 374886 243596
rect 401594 243584 401600 243596
rect 401652 243584 401658 243636
rect 368382 243516 368388 243568
rect 368440 243556 368446 243568
rect 373442 243556 373448 243568
rect 368440 243528 373448 243556
rect 368440 243516 368446 243528
rect 373442 243516 373448 243528
rect 373500 243556 373506 243568
rect 400214 243556 400220 243568
rect 373500 243528 400220 243556
rect 373500 243516 373506 243528
rect 400214 243516 400220 243528
rect 400272 243516 400278 243568
rect 356882 242632 356888 242684
rect 356940 242672 356946 242684
rect 361574 242672 361580 242684
rect 356940 242644 361580 242672
rect 356940 242632 356946 242644
rect 361574 242632 361580 242644
rect 361632 242632 361638 242684
rect 196710 242088 196716 242140
rect 196768 242128 196774 242140
rect 201494 242128 201500 242140
rect 196768 242100 201500 242128
rect 196768 242088 196774 242100
rect 201494 242088 201500 242100
rect 201552 242088 201558 242140
rect 54386 241544 54392 241596
rect 54444 241584 54450 241596
rect 64874 241584 64880 241596
rect 54444 241556 64880 241584
rect 54444 241544 54450 241556
rect 64874 241544 64880 241556
rect 64932 241584 64938 241596
rect 64932 241556 66208 241584
rect 64932 241544 64938 241556
rect 53006 241476 53012 241528
rect 53064 241516 53070 241528
rect 66070 241516 66076 241528
rect 53064 241488 66076 241516
rect 53064 241476 53070 241488
rect 66070 241476 66076 241488
rect 66128 241476 66134 241528
rect 46106 241408 46112 241460
rect 46164 241448 46170 241460
rect 46290 241448 46296 241460
rect 46164 241420 46296 241448
rect 46164 241408 46170 241420
rect 46290 241408 46296 241420
rect 46348 241408 46354 241460
rect 47854 241408 47860 241460
rect 47912 241448 47918 241460
rect 48038 241448 48044 241460
rect 47912 241420 48044 241448
rect 47912 241408 47918 241420
rect 48038 241408 48044 241420
rect 48096 241448 48102 241460
rect 66180 241448 66208 241556
rect 357250 241476 357256 241528
rect 357308 241516 357314 241528
rect 360194 241516 360200 241528
rect 357308 241488 360200 241516
rect 357308 241476 357314 241488
rect 360194 241476 360200 241488
rect 360252 241476 360258 241528
rect 99374 241448 99380 241460
rect 48096 241420 55214 241448
rect 66180 241420 99380 241448
rect 48096 241408 48102 241420
rect 47486 241340 47492 241392
rect 47544 241380 47550 241392
rect 48130 241380 48136 241392
rect 47544 241352 48136 241380
rect 47544 241340 47550 241352
rect 48130 241340 48136 241352
rect 48188 241340 48194 241392
rect 55186 241380 55214 241420
rect 99374 241408 99380 241420
rect 99432 241408 99438 241460
rect 210970 241408 210976 241460
rect 211028 241448 211034 241460
rect 214282 241448 214288 241460
rect 211028 241420 214288 241448
rect 211028 241408 211034 241420
rect 214282 241408 214288 241420
rect 214340 241408 214346 241460
rect 214650 241408 214656 241460
rect 214708 241448 214714 241460
rect 216766 241448 216772 241460
rect 214708 241420 216772 241448
rect 214708 241408 214714 241420
rect 216766 241408 216772 241420
rect 216824 241448 216830 241460
rect 240134 241448 240140 241460
rect 216824 241420 240140 241448
rect 216824 241408 216830 241420
rect 240134 241408 240140 241420
rect 240192 241408 240198 241460
rect 275922 241408 275928 241460
rect 275980 241448 275986 241460
rect 356606 241448 356612 241460
rect 275980 241420 356612 241448
rect 275980 241408 275986 241420
rect 356606 241408 356612 241420
rect 356664 241408 356670 241460
rect 374454 241408 374460 241460
rect 374512 241448 374518 241460
rect 375190 241448 375196 241460
rect 374512 241420 375196 241448
rect 374512 241408 374518 241420
rect 375190 241408 375196 241420
rect 375248 241408 375254 241460
rect 375742 241408 375748 241460
rect 375800 241448 375806 241460
rect 376478 241448 376484 241460
rect 375800 241420 376484 241448
rect 375800 241408 375806 241420
rect 376478 241408 376484 241420
rect 376536 241448 376542 241460
rect 376536 241420 377996 241448
rect 376536 241408 376542 241420
rect 81434 241380 81440 241392
rect 55186 241352 81440 241380
rect 81434 241340 81440 241352
rect 81492 241340 81498 241392
rect 219526 241340 219532 241392
rect 219584 241380 219590 241392
rect 221182 241380 221188 241392
rect 219584 241352 221188 241380
rect 219584 241340 219590 241352
rect 221182 241340 221188 241352
rect 221240 241380 221246 241392
rect 253934 241380 253940 241392
rect 221240 241352 253940 241380
rect 221240 241340 221246 241352
rect 253934 241340 253940 241352
rect 253992 241340 253998 241392
rect 277302 241340 277308 241392
rect 277360 241380 277366 241392
rect 356974 241380 356980 241392
rect 277360 241352 356980 241380
rect 277360 241340 277366 241352
rect 356974 241340 356980 241352
rect 357032 241340 357038 241392
rect 46290 241272 46296 241324
rect 46348 241312 46354 241324
rect 78674 241312 78680 241324
rect 46348 241284 78680 241312
rect 46348 241272 46354 241284
rect 78674 241272 78680 241284
rect 78732 241272 78738 241324
rect 212994 241272 213000 241324
rect 213052 241312 213058 241324
rect 214926 241312 214932 241324
rect 213052 241284 214932 241312
rect 213052 241272 213058 241284
rect 214926 241272 214932 241284
rect 214984 241312 214990 241324
rect 247126 241312 247132 241324
rect 214984 241284 247132 241312
rect 214984 241272 214990 241284
rect 247126 241272 247132 241284
rect 247184 241272 247190 241324
rect 278682 241272 278688 241324
rect 278740 241312 278746 241324
rect 357526 241312 357532 241324
rect 278740 241284 357532 241312
rect 278740 241272 278746 241284
rect 357526 241272 357532 241284
rect 357584 241272 357590 241324
rect 376478 241272 376484 241324
rect 376536 241312 376542 241324
rect 377490 241312 377496 241324
rect 376536 241284 377496 241312
rect 376536 241272 376542 241284
rect 377490 241272 377496 241284
rect 377548 241272 377554 241324
rect 377968 241312 377996 241420
rect 378594 241408 378600 241460
rect 378652 241448 378658 241460
rect 379882 241448 379888 241460
rect 378652 241420 379888 241448
rect 378652 241408 378658 241420
rect 379882 241408 379888 241420
rect 379940 241448 379946 241460
rect 412726 241448 412732 241460
rect 379940 241420 412732 241448
rect 379940 241408 379946 241420
rect 412726 241408 412732 241420
rect 412784 241408 412790 241460
rect 438762 241408 438768 241460
rect 438820 241448 438826 241460
rect 516594 241448 516600 241460
rect 438820 241420 516600 241448
rect 438820 241408 438826 241420
rect 516594 241408 516600 241420
rect 516652 241408 516658 241460
rect 378042 241340 378048 241392
rect 378100 241380 378106 241392
rect 378686 241380 378692 241392
rect 378100 241352 378692 241380
rect 378100 241340 378106 241352
rect 378686 241340 378692 241352
rect 378744 241340 378750 241392
rect 408494 241380 408500 241392
rect 378796 241352 408500 241380
rect 378796 241312 378824 241352
rect 408494 241340 408500 241352
rect 408552 241340 408558 241392
rect 377968 241284 378824 241312
rect 379422 241272 379428 241324
rect 379480 241312 379486 241324
rect 407206 241312 407212 241324
rect 379480 241284 407212 241312
rect 379480 241272 379486 241284
rect 407206 241272 407212 241284
rect 407264 241272 407270 241324
rect 47578 241204 47584 241256
rect 47636 241244 47642 241256
rect 80054 241244 80060 241256
rect 47636 241216 80060 241244
rect 47636 241204 47642 241216
rect 80054 241204 80060 241216
rect 80112 241204 80118 241256
rect 219618 241204 219624 241256
rect 219676 241244 219682 241256
rect 220262 241244 220268 241256
rect 219676 241216 220268 241244
rect 219676 241204 219682 241216
rect 220262 241204 220268 241216
rect 220320 241244 220326 241256
rect 251174 241244 251180 241256
rect 220320 241216 251180 241244
rect 220320 241204 220326 241216
rect 251174 241204 251180 241216
rect 251232 241204 251238 241256
rect 339402 241204 339408 241256
rect 339460 241244 339466 241256
rect 357250 241244 357256 241256
rect 339460 241216 357256 241244
rect 339460 241204 339466 241216
rect 357250 241204 357256 241216
rect 357308 241204 357314 241256
rect 377582 241204 377588 241256
rect 377640 241244 377646 241256
rect 379790 241244 379796 241256
rect 377640 241216 379796 241244
rect 377640 241204 377646 241216
rect 379790 241204 379796 241216
rect 379848 241244 379854 241256
rect 411254 241244 411260 241256
rect 379848 241216 411260 241244
rect 379848 241204 379854 241216
rect 411254 241204 411260 241216
rect 411312 241204 411318 241256
rect 48130 241136 48136 241188
rect 48188 241176 48194 241188
rect 77294 241176 77300 241188
rect 48188 241148 77300 241176
rect 48188 241136 48194 241148
rect 77294 241136 77300 241148
rect 77352 241136 77358 241188
rect 219894 241136 219900 241188
rect 219952 241176 219958 241188
rect 220630 241176 220636 241188
rect 219952 241148 220636 241176
rect 219952 241136 219958 241148
rect 220630 241136 220636 241148
rect 220688 241176 220694 241188
rect 251266 241176 251272 241188
rect 220688 241148 251272 241176
rect 220688 241136 220694 241148
rect 251266 241136 251272 241148
rect 251324 241136 251330 241188
rect 373810 241136 373816 241188
rect 373868 241176 373874 241188
rect 404354 241176 404360 241188
rect 373868 241148 404360 241176
rect 373868 241136 373874 241148
rect 404354 241136 404360 241148
rect 404412 241136 404418 241188
rect 66254 241068 66260 241120
rect 66312 241108 66318 241120
rect 96614 241108 96620 241120
rect 66312 241080 96620 241108
rect 66312 241068 66318 241080
rect 96614 241068 96620 241080
rect 96672 241068 96678 241120
rect 219802 241068 219808 241120
rect 219860 241108 219866 241120
rect 220078 241108 220084 241120
rect 219860 241080 220084 241108
rect 219860 241068 219866 241080
rect 220078 241068 220084 241080
rect 220136 241108 220142 241120
rect 249794 241108 249800 241120
rect 220136 241080 249800 241108
rect 220136 241068 220142 241080
rect 249794 241068 249800 241080
rect 249852 241068 249858 241120
rect 377674 241068 377680 241120
rect 377732 241108 377738 241120
rect 379698 241108 379704 241120
rect 377732 241080 379704 241108
rect 377732 241068 377738 241080
rect 379698 241068 379704 241080
rect 379756 241108 379762 241120
rect 409874 241108 409880 241120
rect 379756 241080 409880 241108
rect 379756 241068 379762 241080
rect 409874 241068 409880 241080
rect 409932 241068 409938 241120
rect 180150 241000 180156 241052
rect 180208 241040 180214 241052
rect 196618 241040 196624 241052
rect 180208 241012 196624 241040
rect 180208 241000 180214 241012
rect 196618 241000 196624 241012
rect 196676 241000 196682 241052
rect 220722 241000 220728 241052
rect 220780 241040 220786 241052
rect 248414 241040 248420 241052
rect 220780 241012 248420 241040
rect 220780 241000 220786 241012
rect 248414 241000 248420 241012
rect 248472 241000 248478 241052
rect 376662 241000 376668 241052
rect 376720 241040 376726 241052
rect 402974 241040 402980 241052
rect 376720 241012 402980 241040
rect 376720 241000 376726 241012
rect 402974 241000 402980 241012
rect 403032 241000 403038 241052
rect 183370 240932 183376 240984
rect 183428 240972 183434 240984
rect 200114 240972 200120 240984
rect 183428 240944 200120 240972
rect 183428 240932 183434 240944
rect 200114 240932 200120 240944
rect 200172 240932 200178 240984
rect 210878 240932 210884 240984
rect 210936 240972 210942 240984
rect 237374 240972 237380 240984
rect 210936 240944 237380 240972
rect 210936 240932 210942 240944
rect 237374 240932 237380 240944
rect 237432 240932 237438 240984
rect 377490 240932 377496 240984
rect 377548 240972 377554 240984
rect 403066 240972 403072 240984
rect 377548 240944 403072 240972
rect 377548 240932 377554 240944
rect 403066 240932 403072 240944
rect 403124 240932 403130 240984
rect 503622 240932 503628 240984
rect 503680 240972 503686 240984
rect 517882 240972 517888 240984
rect 503680 240944 517888 240972
rect 503680 240932 503686 240944
rect 517882 240932 517888 240944
rect 517940 240932 517946 240984
rect 179322 240864 179328 240916
rect 179380 240904 179386 240916
rect 196710 240904 196716 240916
rect 179380 240876 196716 240904
rect 179380 240864 179386 240876
rect 196710 240864 196716 240876
rect 196768 240864 196774 240916
rect 213362 240864 213368 240916
rect 213420 240904 213426 240916
rect 218974 240904 218980 240916
rect 213420 240876 218980 240904
rect 213420 240864 213426 240876
rect 218974 240864 218980 240876
rect 219032 240904 219038 240916
rect 245654 240904 245660 240916
rect 219032 240876 245660 240904
rect 219032 240864 219038 240876
rect 245654 240864 245660 240876
rect 245712 240864 245718 240916
rect 343450 240864 343456 240916
rect 343508 240904 343514 240916
rect 359458 240904 359464 240916
rect 343508 240876 359464 240904
rect 343508 240864 343514 240876
rect 359458 240864 359464 240876
rect 359516 240864 359522 240916
rect 372522 240864 372528 240916
rect 372580 240904 372586 240916
rect 379054 240904 379060 240916
rect 372580 240876 379060 240904
rect 372580 240864 372586 240876
rect 379054 240864 379060 240876
rect 379112 240904 379118 240916
rect 405734 240904 405740 240916
rect 379112 240876 405740 240904
rect 379112 240864 379118 240876
rect 405734 240864 405740 240876
rect 405792 240864 405798 240916
rect 500770 240864 500776 240916
rect 500828 240904 500834 240916
rect 517698 240904 517704 240916
rect 500828 240876 517704 240904
rect 500828 240864 500834 240876
rect 517698 240864 517704 240876
rect 517756 240864 517762 240916
rect 183462 240796 183468 240848
rect 183520 240836 183526 240848
rect 201494 240836 201500 240848
rect 183520 240808 201500 240836
rect 183520 240796 183526 240808
rect 201494 240796 201500 240808
rect 201552 240796 201558 240848
rect 214282 240796 214288 240848
rect 214340 240836 214346 240848
rect 244274 240836 244280 240848
rect 214340 240808 244280 240836
rect 214340 240796 214346 240808
rect 244274 240796 244280 240808
rect 244332 240796 244338 240848
rect 340046 240796 340052 240848
rect 340104 240836 340110 240848
rect 356882 240836 356888 240848
rect 340104 240808 356888 240836
rect 340104 240796 340110 240808
rect 356882 240796 356888 240808
rect 356940 240796 356946 240848
rect 375098 240796 375104 240848
rect 375156 240836 375162 240848
rect 375156 240808 378640 240836
rect 375156 240796 375162 240808
rect 67542 240728 67548 240780
rect 67600 240768 67606 240780
rect 97994 240768 98000 240780
rect 67600 240740 98000 240768
rect 67600 240728 67606 240740
rect 97994 240728 98000 240740
rect 98052 240728 98058 240780
rect 209498 240728 209504 240780
rect 209556 240768 209562 240780
rect 210786 240768 210792 240780
rect 209556 240740 210792 240768
rect 209556 240728 209562 240740
rect 210786 240728 210792 240740
rect 210844 240768 210850 240780
rect 241514 240768 241520 240780
rect 210844 240740 241520 240768
rect 210844 240728 210850 240740
rect 241514 240728 241520 240740
rect 241572 240728 241578 240780
rect 351546 240728 351552 240780
rect 351604 240768 351610 240780
rect 358078 240768 358084 240780
rect 351604 240740 358084 240768
rect 351604 240728 351610 240740
rect 358078 240728 358084 240740
rect 358136 240728 358142 240780
rect 375650 240728 375656 240780
rect 375708 240768 375714 240780
rect 376662 240768 376668 240780
rect 375708 240740 376668 240768
rect 375708 240728 375714 240740
rect 376662 240728 376668 240740
rect 376720 240728 376726 240780
rect 378612 240768 378640 240808
rect 378686 240796 378692 240848
rect 378744 240836 378750 240848
rect 411346 240836 411352 240848
rect 378744 240808 411352 240836
rect 378744 240796 378750 240808
rect 411346 240796 411352 240808
rect 411404 240796 411410 240848
rect 499022 240796 499028 240848
rect 499080 240836 499086 240848
rect 517790 240836 517796 240848
rect 499080 240808 517796 240836
rect 499080 240796 499086 240808
rect 517790 240796 517796 240808
rect 517848 240796 517854 240848
rect 379422 240768 379428 240780
rect 378612 240740 379428 240768
rect 379422 240728 379428 240740
rect 379480 240728 379486 240780
rect 379882 240728 379888 240780
rect 379940 240768 379946 240780
rect 414014 240768 414020 240780
rect 379940 240740 414020 240768
rect 379940 240728 379946 240740
rect 414014 240728 414020 240740
rect 414072 240728 414078 240780
rect 218330 240660 218336 240712
rect 218388 240700 218394 240712
rect 219342 240700 219348 240712
rect 218388 240672 219348 240700
rect 218388 240660 218394 240672
rect 219342 240660 219348 240672
rect 219400 240700 219406 240712
rect 252646 240700 252652 240712
rect 219400 240672 252652 240700
rect 219400 240660 219406 240672
rect 252646 240660 252652 240672
rect 252704 240660 252710 240712
rect 369670 240660 369676 240712
rect 369728 240700 369734 240712
rect 372522 240700 372528 240712
rect 369728 240672 372528 240700
rect 369728 240660 369734 240672
rect 372522 240660 372528 240672
rect 372580 240700 372586 240712
rect 397454 240700 397460 240712
rect 372580 240672 397460 240700
rect 372580 240660 372586 240672
rect 397454 240660 397460 240672
rect 397512 240660 397518 240712
rect 238754 240632 238760 240644
rect 219406 240604 238760 240632
rect 213546 240524 213552 240576
rect 213604 240564 213610 240576
rect 216306 240564 216312 240576
rect 213604 240536 216312 240564
rect 213604 240524 213610 240536
rect 216306 240524 216312 240536
rect 216364 240564 216370 240576
rect 219406 240564 219434 240604
rect 238754 240592 238760 240604
rect 238812 240592 238818 240644
rect 374546 240592 374552 240644
rect 374604 240632 374610 240644
rect 396166 240632 396172 240644
rect 374604 240604 396172 240632
rect 374604 240592 374610 240604
rect 396166 240592 396172 240604
rect 396224 240592 396230 240644
rect 511902 240592 511908 240644
rect 511960 240632 511966 240644
rect 517514 240632 517520 240644
rect 511960 240604 517520 240632
rect 511960 240592 511966 240604
rect 517514 240592 517520 240604
rect 517572 240592 517578 240644
rect 216364 240536 219434 240564
rect 216364 240524 216370 240536
rect 375190 240456 375196 240508
rect 375248 240496 375254 240508
rect 396074 240496 396080 240508
rect 375248 240468 396080 240496
rect 375248 240456 375254 240468
rect 396074 240456 396080 240468
rect 396132 240456 396138 240508
rect 216306 240388 216312 240440
rect 216364 240428 216370 240440
rect 219710 240428 219716 240440
rect 216364 240400 219716 240428
rect 216364 240388 216370 240400
rect 219710 240388 219716 240400
rect 219768 240428 219774 240440
rect 220722 240428 220728 240440
rect 219768 240400 220728 240428
rect 219768 240388 219774 240400
rect 220722 240388 220728 240400
rect 220780 240388 220786 240440
rect 217594 240252 217600 240304
rect 217652 240292 217658 240304
rect 220262 240292 220268 240304
rect 217652 240264 220268 240292
rect 217652 240252 217658 240264
rect 220262 240252 220268 240264
rect 220320 240252 220326 240304
rect 190914 240184 190920 240236
rect 190972 240224 190978 240236
rect 197998 240224 198004 240236
rect 190972 240196 198004 240224
rect 190972 240184 190978 240196
rect 197998 240184 198004 240196
rect 198056 240184 198062 240236
rect 219342 240184 219348 240236
rect 219400 240224 219406 240236
rect 220630 240224 220636 240236
rect 219400 240196 220636 240224
rect 219400 240184 219406 240196
rect 220630 240184 220636 240196
rect 220688 240184 220694 240236
rect 50614 240048 50620 240100
rect 50672 240088 50678 240100
rect 53098 240088 53104 240100
rect 50672 240060 53104 240088
rect 50672 240048 50678 240060
rect 53098 240048 53104 240060
rect 53156 240048 53162 240100
rect 58986 240048 58992 240100
rect 59044 240088 59050 240100
rect 62298 240088 62304 240100
rect 59044 240060 62304 240088
rect 59044 240048 59050 240060
rect 62298 240048 62304 240060
rect 62356 240048 62362 240100
rect 214926 240048 214932 240100
rect 214984 240088 214990 240100
rect 215294 240088 215300 240100
rect 214984 240060 215300 240088
rect 214984 240048 214990 240060
rect 215294 240048 215300 240060
rect 215352 240048 215358 240100
rect 219894 240048 219900 240100
rect 219952 240088 219958 240100
rect 221090 240088 221096 240100
rect 219952 240060 221096 240088
rect 219952 240048 219958 240060
rect 221090 240048 221096 240060
rect 221148 240048 221154 240100
rect 222102 240048 222108 240100
rect 222160 240088 222166 240100
rect 267734 240088 267740 240100
rect 222160 240060 267740 240088
rect 222160 240048 222166 240060
rect 267734 240048 267740 240060
rect 267792 240048 267798 240100
rect 371142 240048 371148 240100
rect 371200 240088 371206 240100
rect 373166 240088 373172 240100
rect 371200 240060 373172 240088
rect 371200 240048 371206 240060
rect 373166 240048 373172 240060
rect 373224 240048 373230 240100
rect 376570 240048 376576 240100
rect 376628 240088 376634 240100
rect 436094 240088 436100 240100
rect 376628 240060 436100 240088
rect 376628 240048 376634 240060
rect 436094 240048 436100 240060
rect 436152 240048 436158 240100
rect 58802 239980 58808 240032
rect 58860 240020 58866 240032
rect 62206 240020 62212 240032
rect 58860 239992 62212 240020
rect 58860 239980 58866 239992
rect 62206 239980 62212 239992
rect 62264 239980 62270 240032
rect 213638 239980 213644 240032
rect 213696 240020 213702 240032
rect 215662 240020 215668 240032
rect 213696 239992 215668 240020
rect 213696 239980 213702 239992
rect 215662 239980 215668 239992
rect 215720 239980 215726 240032
rect 218606 239980 218612 240032
rect 218664 240020 218670 240032
rect 219250 240020 219256 240032
rect 218664 239992 219256 240020
rect 218664 239980 218670 239992
rect 219250 239980 219256 239992
rect 219308 240020 219314 240032
rect 264974 240020 264980 240032
rect 219308 239992 264980 240020
rect 219308 239980 219314 239992
rect 264974 239980 264980 239992
rect 265032 239980 265038 240032
rect 375282 239980 375288 240032
rect 375340 240020 375346 240032
rect 434714 240020 434720 240032
rect 375340 239992 434720 240020
rect 375340 239980 375346 239992
rect 434714 239980 434720 239992
rect 434772 239980 434778 240032
rect 55674 239912 55680 239964
rect 55732 239952 55738 239964
rect 60734 239952 60740 239964
rect 55732 239924 60740 239952
rect 55732 239912 55738 239924
rect 60734 239912 60740 239924
rect 60792 239912 60798 239964
rect 216398 239912 216404 239964
rect 216456 239952 216462 239964
rect 262214 239952 262220 239964
rect 216456 239924 262220 239952
rect 216456 239912 216462 239924
rect 262214 239912 262220 239924
rect 262272 239912 262278 239964
rect 378042 239912 378048 239964
rect 378100 239952 378106 239964
rect 423674 239952 423680 239964
rect 378100 239924 423680 239952
rect 378100 239912 378106 239924
rect 423674 239912 423680 239924
rect 423732 239912 423738 239964
rect 219802 239844 219808 239896
rect 219860 239884 219866 239896
rect 220814 239884 220820 239896
rect 219860 239856 220820 239884
rect 219860 239844 219866 239856
rect 220814 239844 220820 239856
rect 220872 239844 220878 239896
rect 221090 239844 221096 239896
rect 221148 239884 221154 239896
rect 266446 239884 266452 239896
rect 221148 239856 266452 239884
rect 221148 239844 221154 239856
rect 266446 239844 266452 239856
rect 266504 239844 266510 239896
rect 369762 239844 369768 239896
rect 369820 239884 369826 239896
rect 379698 239884 379704 239896
rect 369820 239856 379704 239884
rect 369820 239844 369826 239856
rect 379698 239844 379704 239856
rect 379756 239884 379762 239896
rect 425698 239884 425704 239896
rect 379756 239856 425704 239884
rect 379756 239844 379762 239856
rect 425698 239844 425704 239856
rect 425756 239844 425762 239896
rect 53098 239776 53104 239828
rect 53156 239816 53162 239828
rect 67542 239816 67548 239828
rect 53156 239788 67548 239816
rect 53156 239776 53162 239788
rect 67542 239776 67548 239788
rect 67600 239776 67606 239828
rect 217226 239776 217232 239828
rect 217284 239816 217290 239828
rect 217962 239816 217968 239828
rect 217284 239788 217968 239816
rect 217284 239776 217290 239788
rect 217962 239776 217968 239788
rect 218020 239776 218026 239828
rect 219158 239776 219164 239828
rect 219216 239816 219222 239828
rect 220722 239816 220728 239828
rect 219216 239788 220728 239816
rect 219216 239776 219222 239788
rect 220722 239776 220728 239788
rect 220780 239776 220786 239828
rect 220832 239816 220860 239844
rect 222102 239816 222108 239828
rect 220832 239788 222108 239816
rect 222102 239776 222108 239788
rect 222160 239776 222166 239828
rect 222194 239776 222200 239828
rect 222252 239816 222258 239828
rect 266354 239816 266360 239828
rect 222252 239788 266360 239816
rect 222252 239776 222258 239788
rect 266354 239776 266360 239788
rect 266412 239776 266418 239828
rect 57146 239708 57152 239760
rect 57204 239748 57210 239760
rect 82078 239748 82084 239760
rect 57204 239720 82084 239748
rect 57204 239708 57210 239720
rect 82078 239708 82084 239720
rect 82136 239708 82142 239760
rect 215294 239708 215300 239760
rect 215352 239748 215358 239760
rect 259546 239748 259552 239760
rect 215352 239720 259552 239748
rect 215352 239708 215358 239720
rect 259546 239708 259552 239720
rect 259604 239708 259610 239760
rect 53834 239640 53840 239692
rect 53892 239680 53898 239692
rect 100018 239680 100024 239692
rect 53892 239652 100024 239680
rect 53892 239640 53898 239652
rect 100018 239640 100024 239652
rect 100076 239640 100082 239692
rect 219618 239640 219624 239692
rect 219676 239680 219682 239692
rect 220906 239680 220912 239692
rect 219676 239652 220912 239680
rect 219676 239640 219682 239652
rect 220906 239640 220912 239652
rect 220964 239680 220970 239692
rect 263594 239680 263600 239692
rect 220964 239652 263600 239680
rect 220964 239640 220970 239652
rect 263594 239640 263600 239652
rect 263652 239640 263658 239692
rect 60642 239572 60648 239624
rect 60700 239612 60706 239624
rect 107654 239612 107660 239624
rect 60700 239584 107660 239612
rect 60700 239572 60706 239584
rect 107654 239572 107660 239584
rect 107712 239572 107718 239624
rect 217042 239572 217048 239624
rect 217100 239612 217106 239624
rect 219066 239612 219072 239624
rect 217100 239584 219072 239612
rect 217100 239572 217106 239584
rect 219066 239572 219072 239584
rect 219124 239612 219130 239624
rect 258166 239612 258172 239624
rect 219124 239584 258172 239612
rect 219124 239572 219130 239584
rect 258166 239572 258172 239584
rect 258224 239572 258230 239624
rect 58894 239504 58900 239556
rect 58952 239544 58958 239556
rect 107746 239544 107752 239556
rect 58952 239516 107752 239544
rect 58952 239504 58958 239516
rect 107746 239504 107752 239516
rect 107804 239504 107810 239556
rect 215662 239504 215668 239556
rect 215720 239544 215726 239556
rect 256694 239544 256700 239556
rect 215720 239516 256700 239544
rect 215720 239504 215726 239516
rect 256694 239504 256700 239516
rect 256752 239504 256758 239556
rect 50798 239436 50804 239488
rect 50856 239476 50862 239488
rect 110414 239476 110420 239488
rect 50856 239448 110420 239476
rect 50856 239436 50862 239448
rect 110414 239436 110420 239448
rect 110472 239436 110478 239488
rect 218514 239436 218520 239488
rect 218572 239476 218578 239488
rect 259454 239476 259460 239488
rect 218572 239448 259460 239476
rect 218572 239436 218578 239448
rect 259454 239436 259460 239448
rect 259512 239436 259518 239488
rect 51810 239368 51816 239420
rect 51868 239408 51874 239420
rect 113174 239408 113180 239420
rect 51868 239380 113180 239408
rect 51868 239368 51874 239380
rect 113174 239368 113180 239380
rect 113232 239368 113238 239420
rect 216214 239368 216220 239420
rect 216272 239408 216278 239420
rect 260834 239408 260840 239420
rect 216272 239380 260840 239408
rect 216272 239368 216278 239380
rect 260834 239368 260840 239380
rect 260892 239368 260898 239420
rect 373166 239368 373172 239420
rect 373224 239408 373230 239420
rect 430666 239408 430672 239420
rect 373224 239380 430672 239408
rect 373224 239368 373230 239380
rect 430666 239368 430672 239380
rect 430724 239368 430730 239420
rect 217962 239300 217968 239352
rect 218020 239340 218026 239352
rect 255314 239340 255320 239352
rect 218020 239312 255320 239340
rect 218020 239300 218026 239312
rect 255314 239300 255320 239312
rect 255372 239300 255378 239352
rect 57238 239232 57244 239284
rect 57296 239272 57302 239284
rect 62114 239272 62120 239284
rect 57296 239244 62120 239272
rect 57296 239232 57302 239244
rect 62114 239232 62120 239244
rect 62172 239232 62178 239284
rect 220814 239232 220820 239284
rect 220872 239272 220878 239284
rect 222102 239272 222108 239284
rect 220872 239244 222108 239272
rect 220872 239232 220878 239244
rect 222102 239232 222108 239244
rect 222160 239232 222166 239284
rect 375926 239232 375932 239284
rect 375984 239272 375990 239284
rect 376570 239272 376576 239284
rect 375984 239244 376576 239272
rect 375984 239232 375990 239244
rect 376570 239232 376576 239244
rect 376628 239232 376634 239284
rect 372430 238756 372436 238808
rect 372488 238796 372494 238808
rect 375282 238796 375288 238808
rect 372488 238768 375288 238796
rect 372488 238756 372494 238768
rect 375282 238756 375288 238768
rect 375340 238756 375346 238808
rect 46842 238688 46848 238740
rect 46900 238728 46906 238740
rect 50798 238728 50804 238740
rect 46900 238700 50804 238728
rect 46900 238688 46906 238700
rect 50798 238688 50804 238700
rect 50856 238688 50862 238740
rect 214466 238688 214472 238740
rect 214524 238728 214530 238740
rect 216214 238728 216220 238740
rect 214524 238700 216220 238728
rect 214524 238688 214530 238700
rect 216214 238688 216220 238700
rect 216272 238688 216278 238740
rect 42334 238620 42340 238672
rect 42392 238660 42398 238672
rect 42392 238632 45554 238660
rect 42392 238620 42398 238632
rect 45526 238524 45554 238632
rect 46750 238620 46756 238672
rect 46808 238660 46814 238672
rect 51810 238660 51816 238672
rect 46808 238632 51816 238660
rect 46808 238620 46814 238632
rect 51810 238620 51816 238632
rect 51868 238620 51874 238672
rect 215202 238620 215208 238672
rect 215260 238660 215266 238672
rect 218514 238660 218520 238672
rect 215260 238632 218520 238660
rect 215260 238620 215266 238632
rect 218514 238620 218520 238632
rect 218572 238620 218578 238672
rect 47946 238552 47952 238604
rect 48004 238592 48010 238604
rect 60642 238592 60648 238604
rect 48004 238564 60648 238592
rect 48004 238552 48010 238564
rect 60642 238552 60648 238564
rect 60700 238552 60706 238604
rect 53834 238524 53840 238536
rect 45526 238496 53840 238524
rect 53834 238484 53840 238496
rect 53892 238484 53898 238536
rect 43806 238416 43812 238468
rect 43864 238456 43870 238468
rect 57146 238456 57152 238468
rect 43864 238428 57152 238456
rect 43864 238416 43870 238428
rect 57146 238416 57152 238428
rect 57204 238416 57210 238468
rect 50338 237396 50344 237448
rect 50396 237436 50402 237448
rect 50798 237436 50804 237448
rect 50396 237408 50804 237436
rect 50396 237396 50402 237408
rect 50798 237396 50804 237408
rect 50856 237396 50862 237448
rect 51534 237396 51540 237448
rect 51592 237436 51598 237448
rect 51810 237436 51816 237448
rect 51592 237408 51816 237436
rect 51592 237396 51598 237408
rect 51810 237396 51816 237408
rect 51868 237396 51874 237448
rect 53834 237396 53840 237448
rect 53892 237436 53898 237448
rect 54478 237436 54484 237448
rect 53892 237408 54484 237436
rect 53892 237396 53898 237408
rect 54478 237396 54484 237408
rect 54536 237396 54542 237448
rect 56962 235968 56968 236020
rect 57020 236008 57026 236020
rect 59722 236008 59728 236020
rect 57020 235980 59728 236008
rect 57020 235968 57026 235980
rect 59722 235968 59728 235980
rect 59780 235968 59786 236020
rect 2866 169668 2872 169720
rect 2924 169708 2930 169720
rect 4798 169708 4804 169720
rect 2924 169680 4804 169708
rect 2924 169668 2930 169680
rect 4798 169668 4804 169680
rect 4856 169668 4862 169720
rect 207750 165520 207756 165572
rect 207808 165560 207814 165572
rect 216674 165560 216680 165572
rect 207808 165532 216680 165560
rect 207808 165520 207814 165532
rect 216674 165520 216680 165532
rect 216732 165520 216738 165572
rect 362402 165520 362408 165572
rect 362460 165560 362466 165572
rect 376938 165560 376944 165572
rect 362460 165532 376944 165560
rect 362460 165520 362466 165532
rect 376938 165520 376944 165532
rect 376996 165520 377002 165572
rect 377766 165112 377772 165164
rect 377824 165152 377830 165164
rect 377950 165152 377956 165164
rect 377824 165124 377956 165152
rect 377824 165112 377830 165124
rect 377950 165112 377956 165124
rect 378008 165112 378014 165164
rect 203610 164160 203616 164212
rect 203668 164200 203674 164212
rect 217042 164200 217048 164212
rect 203668 164172 217048 164200
rect 203668 164160 203674 164172
rect 217042 164160 217048 164172
rect 217100 164160 217106 164212
rect 367830 164160 367836 164212
rect 367888 164200 367894 164212
rect 376754 164200 376760 164212
rect 367888 164172 376760 164200
rect 367888 164160 367894 164172
rect 376754 164160 376760 164172
rect 376812 164160 376818 164212
rect 197998 163480 198004 163532
rect 198056 163520 198062 163532
rect 216674 163520 216680 163532
rect 198056 163492 216680 163520
rect 198056 163480 198062 163492
rect 216674 163480 216680 163492
rect 216732 163480 216738 163532
rect 358078 163480 358084 163532
rect 358136 163520 358142 163532
rect 376938 163520 376944 163532
rect 358136 163492 376944 163520
rect 358136 163480 358142 163492
rect 376938 163480 376944 163492
rect 376996 163480 377002 163532
rect 377766 156612 377772 156664
rect 377824 156652 377830 156664
rect 377950 156652 377956 156664
rect 377824 156624 377956 156652
rect 377824 156612 377830 156624
rect 377950 156612 377956 156624
rect 378008 156612 378014 156664
rect 42426 154640 42432 154692
rect 42484 154680 42490 154692
rect 163314 154680 163320 154692
rect 42484 154652 163320 154680
rect 42484 154640 42490 154652
rect 163314 154640 163320 154652
rect 163372 154640 163378 154692
rect 43898 154572 43904 154624
rect 43956 154612 43962 154624
rect 165890 154612 165896 154624
rect 43956 154584 165896 154612
rect 43956 154572 43962 154584
rect 165890 154572 165896 154584
rect 165948 154572 165954 154624
rect 50338 154504 50344 154556
rect 50396 154544 50402 154556
rect 51810 154544 51816 154556
rect 50396 154516 51816 154544
rect 50396 154504 50402 154516
rect 51810 154504 51816 154516
rect 51868 154504 51874 154556
rect 56962 154504 56968 154556
rect 57020 154544 57026 154556
rect 59354 154544 59360 154556
rect 57020 154516 59360 154544
rect 57020 154504 57026 154516
rect 59354 154504 59360 154516
rect 59412 154504 59418 154556
rect 358262 154504 358268 154556
rect 358320 154544 358326 154556
rect 418430 154544 418436 154556
rect 358320 154516 418436 154544
rect 358320 154504 358326 154516
rect 418430 154504 418436 154516
rect 418488 154504 418494 154556
rect 50706 154436 50712 154488
rect 50764 154476 50770 154488
rect 96062 154476 96068 154488
rect 50764 154448 96068 154476
rect 50764 154436 50770 154448
rect 96062 154436 96068 154448
rect 96120 154436 96126 154488
rect 358354 154436 358360 154488
rect 358412 154476 358418 154488
rect 421006 154476 421012 154488
rect 358412 154448 421012 154476
rect 358412 154436 358418 154448
rect 421006 154436 421012 154448
rect 421064 154436 421070 154488
rect 49510 154368 49516 154420
rect 49568 154408 49574 154420
rect 98454 154408 98460 154420
rect 49568 154380 98460 154408
rect 49568 154368 49574 154380
rect 98454 154368 98460 154380
rect 98512 154368 98518 154420
rect 357618 154368 357624 154420
rect 357676 154408 357682 154420
rect 360286 154408 360292 154420
rect 357676 154380 360292 154408
rect 357676 154368 357682 154380
rect 360286 154368 360292 154380
rect 360344 154368 360350 154420
rect 362310 154368 362316 154420
rect 362368 154408 362374 154420
rect 425974 154408 425980 154420
rect 362368 154380 425980 154408
rect 362368 154368 362374 154380
rect 425974 154368 425980 154380
rect 426032 154368 426038 154420
rect 438854 154368 438860 154420
rect 438912 154408 438918 154420
rect 516594 154408 516600 154420
rect 438912 154380 516600 154408
rect 438912 154368 438918 154380
rect 516594 154368 516600 154380
rect 516652 154368 516658 154420
rect 52086 154300 52092 154352
rect 52144 154340 52150 154352
rect 101030 154340 101036 154352
rect 52144 154312 101036 154340
rect 52144 154300 52150 154312
rect 101030 154300 101036 154312
rect 101088 154300 101094 154352
rect 365254 154300 365260 154352
rect 365312 154340 365318 154352
rect 443454 154340 443460 154352
rect 365312 154312 443460 154340
rect 365312 154300 365318 154312
rect 443454 154300 443460 154312
rect 443512 154300 443518 154352
rect 53558 154232 53564 154284
rect 53616 154272 53622 154284
rect 105814 154272 105820 154284
rect 53616 154244 105820 154272
rect 53616 154232 53622 154244
rect 105814 154232 105820 154244
rect 105872 154232 105878 154284
rect 206462 154232 206468 154284
rect 206520 154272 206526 154284
rect 261018 154272 261024 154284
rect 206520 154244 261024 154272
rect 206520 154232 206526 154244
rect 261018 154232 261024 154244
rect 261076 154232 261082 154284
rect 372154 154232 372160 154284
rect 372212 154272 372218 154284
rect 475838 154272 475844 154284
rect 372212 154244 475844 154272
rect 372212 154232 372218 154244
rect 475838 154232 475844 154244
rect 475896 154232 475902 154284
rect 56318 154164 56324 154216
rect 56376 154204 56382 154216
rect 138382 154204 138388 154216
rect 56376 154176 138388 154204
rect 56376 154164 56382 154176
rect 138382 154164 138388 154176
rect 138440 154164 138446 154216
rect 202138 154164 202144 154216
rect 202196 154204 202202 154216
rect 273530 154204 273536 154216
rect 202196 154176 273536 154204
rect 202196 154164 202202 154176
rect 273530 154164 273536 154176
rect 273588 154164 273594 154216
rect 373350 154164 373356 154216
rect 373408 154204 373414 154216
rect 478414 154204 478420 154216
rect 373408 154176 478420 154204
rect 373408 154164 373414 154176
rect 478414 154164 478420 154176
rect 478472 154164 478478 154216
rect 52178 154096 52184 154148
rect 52236 154136 52242 154148
rect 108206 154136 108212 154148
rect 52236 154108 108212 154136
rect 52236 154096 52242 154108
rect 108206 154096 108212 154108
rect 108264 154096 108270 154148
rect 113358 154096 113364 154148
rect 113416 154136 113422 154148
rect 114462 154136 114468 154148
rect 113416 154108 114468 154136
rect 113416 154096 113422 154108
rect 114462 154096 114468 154108
rect 114520 154136 114526 154148
rect 196802 154136 196808 154148
rect 114520 154108 196808 154136
rect 114520 154096 114526 154108
rect 196802 154096 196808 154108
rect 196860 154096 196866 154148
rect 204990 154096 204996 154148
rect 205048 154136 205054 154148
rect 293310 154136 293316 154148
rect 205048 154108 293316 154136
rect 205048 154096 205054 154108
rect 293310 154096 293316 154108
rect 293368 154096 293374 154148
rect 366634 154096 366640 154148
rect 366692 154136 366698 154148
rect 473446 154136 473452 154148
rect 366692 154108 473452 154136
rect 366692 154096 366698 154108
rect 473446 154096 473452 154108
rect 473504 154096 473510 154148
rect 59262 154028 59268 154080
rect 59320 154068 59326 154080
rect 143534 154068 143540 154080
rect 59320 154040 143540 154068
rect 59320 154028 59326 154040
rect 143534 154028 143540 154040
rect 143592 154028 143598 154080
rect 198090 154028 198096 154080
rect 198148 154068 198154 154080
rect 288158 154068 288164 154080
rect 198148 154040 288164 154068
rect 198148 154028 198154 154040
rect 288158 154028 288164 154040
rect 288216 154028 288222 154080
rect 369210 154028 369216 154080
rect 369268 154068 369274 154080
rect 480806 154068 480812 154080
rect 369268 154040 480812 154068
rect 369268 154028 369274 154040
rect 480806 154028 480812 154040
rect 480864 154028 480870 154080
rect 46382 153960 46388 154012
rect 46440 154000 46446 154012
rect 52178 154000 52184 154012
rect 46440 153972 52184 154000
rect 46440 153960 46446 153972
rect 52178 153960 52184 153972
rect 52236 153960 52242 154012
rect 59906 153960 59912 154012
rect 59964 154000 59970 154012
rect 145926 154000 145932 154012
rect 59964 153972 145932 154000
rect 59964 153960 59970 153972
rect 145926 153960 145932 153972
rect 145984 153960 145990 154012
rect 206370 153960 206376 154012
rect 206428 154000 206434 154012
rect 298462 154000 298468 154012
rect 206428 153972 298468 154000
rect 206428 153960 206434 153972
rect 298462 153960 298468 153972
rect 298520 153960 298526 154012
rect 356790 153960 356796 154012
rect 356848 154000 356854 154012
rect 470870 154000 470876 154012
rect 356848 153972 470876 154000
rect 356848 153960 356854 153972
rect 470870 153960 470876 153972
rect 470928 153960 470934 154012
rect 510522 153960 510528 154012
rect 510580 154000 510586 154012
rect 517514 154000 517520 154012
rect 510580 153972 517520 154000
rect 510580 153960 510586 153972
rect 517514 153960 517520 153972
rect 517572 153960 517578 154012
rect 59998 153892 60004 153944
rect 60056 153932 60062 153944
rect 150894 153932 150900 153944
rect 60056 153904 150900 153932
rect 60056 153892 60062 153904
rect 150894 153892 150900 153904
rect 150952 153892 150958 153944
rect 210510 153892 210516 153944
rect 210568 153932 210574 153944
rect 303430 153932 303436 153944
rect 210568 153904 303436 153932
rect 210568 153892 210574 153904
rect 303430 153892 303436 153904
rect 303488 153892 303494 153944
rect 368014 153892 368020 153944
rect 368072 153932 368078 153944
rect 483198 153932 483204 153944
rect 368072 153904 483204 153932
rect 368072 153892 368078 153904
rect 483198 153892 483204 153904
rect 483256 153892 483262 153944
rect 59170 153824 59176 153876
rect 59228 153864 59234 153876
rect 153286 153864 153292 153876
rect 59228 153836 153292 153864
rect 59228 153824 59234 153836
rect 153286 153824 153292 153836
rect 153344 153824 153350 153876
rect 209222 153824 209228 153876
rect 209280 153864 209286 153876
rect 308398 153864 308404 153876
rect 209280 153836 308404 153864
rect 209280 153824 209286 153836
rect 308398 153824 308404 153836
rect 308456 153824 308462 153876
rect 370774 153824 370780 153876
rect 370832 153864 370838 153876
rect 485958 153864 485964 153876
rect 370832 153836 485964 153864
rect 370832 153824 370838 153836
rect 485958 153824 485964 153836
rect 486016 153824 486022 153876
rect 366542 153756 366548 153808
rect 366600 153796 366606 153808
rect 423398 153796 423404 153808
rect 366600 153768 423404 153796
rect 366600 153756 366606 153768
rect 423398 153756 423404 153768
rect 423456 153756 423462 153808
rect 51810 153348 51816 153400
rect 51868 153388 51874 153400
rect 111150 153388 111156 153400
rect 51868 153360 111156 153388
rect 51868 153348 51874 153360
rect 111150 153348 111156 153360
rect 111208 153348 111214 153400
rect 59354 153280 59360 153332
rect 59412 153320 59418 153332
rect 118694 153320 118700 153332
rect 59412 153292 118700 153320
rect 59412 153280 59418 153292
rect 118694 153280 118700 153292
rect 118752 153280 118758 153332
rect 52178 153212 52184 153264
rect 52236 153252 52242 153264
rect 114738 153252 114744 153264
rect 52236 153224 114744 153252
rect 52236 153212 52242 153224
rect 114738 153212 114744 153224
rect 114796 153212 114802 153264
rect 197354 153212 197360 153264
rect 197412 153252 197418 153264
rect 201494 153252 201500 153264
rect 197412 153224 201500 153252
rect 197412 153212 197418 153224
rect 201494 153212 201500 153224
rect 201552 153212 201558 153264
rect 373626 153212 373632 153264
rect 373684 153252 373690 153264
rect 373810 153252 373816 153264
rect 373684 153224 373816 153252
rect 373684 153212 373690 153224
rect 373810 153212 373816 153224
rect 373868 153252 373874 153264
rect 431954 153252 431960 153264
rect 373868 153224 431960 153252
rect 373868 153212 373874 153224
rect 431954 153212 431960 153224
rect 432012 153212 432018 153264
rect 51902 153144 51908 153196
rect 51960 153184 51966 153196
rect 155954 153184 155960 153196
rect 51960 153156 155960 153184
rect 51960 153144 51966 153156
rect 155954 153144 155960 153156
rect 156012 153144 156018 153196
rect 210418 153144 210424 153196
rect 210476 153184 210482 153196
rect 300854 153184 300860 153196
rect 210476 153156 300860 153184
rect 210476 153144 210482 153156
rect 300854 153144 300860 153156
rect 300912 153144 300918 153196
rect 361114 153144 361120 153196
rect 361172 153184 361178 153196
rect 455414 153184 455420 153196
rect 361172 153156 455420 153184
rect 361172 153144 361178 153156
rect 455414 153144 455420 153156
rect 455472 153144 455478 153196
rect 56134 153076 56140 153128
rect 56192 153116 56198 153128
rect 135254 153116 135260 153128
rect 56192 153088 135260 153116
rect 56192 153076 56198 153088
rect 135254 153076 135260 153088
rect 135312 153076 135318 153128
rect 209038 153076 209044 153128
rect 209096 153116 209102 153128
rect 285674 153116 285680 153128
rect 209096 153088 285680 153116
rect 209096 153076 209102 153088
rect 285674 153076 285680 153088
rect 285732 153076 285738 153128
rect 358446 153076 358452 153128
rect 358504 153116 358510 153128
rect 447134 153116 447140 153128
rect 358504 153088 447140 153116
rect 358504 153076 358510 153088
rect 447134 153076 447140 153088
rect 447192 153076 447198 153128
rect 55950 153008 55956 153060
rect 56008 153048 56014 153060
rect 132770 153048 132776 153060
rect 56008 153020 132776 153048
rect 56008 153008 56014 153020
rect 132770 153008 132776 153020
rect 132828 153008 132834 153060
rect 215938 153008 215944 153060
rect 215996 153048 216002 153060
rect 289814 153048 289820 153060
rect 215996 153020 289820 153048
rect 215996 153008 216002 153020
rect 289814 153008 289820 153020
rect 289872 153008 289878 153060
rect 376110 153008 376116 153060
rect 376168 153048 376174 153060
rect 458174 153048 458180 153060
rect 376168 153020 458180 153048
rect 376168 153008 376174 153020
rect 458174 153008 458180 153020
rect 458232 153008 458238 153060
rect 54846 152940 54852 152992
rect 54904 152980 54910 152992
rect 129734 152980 129740 152992
rect 54904 152952 129740 152980
rect 54904 152940 54910 152952
rect 129734 152940 129740 152952
rect 129792 152940 129798 152992
rect 211982 152940 211988 152992
rect 212040 152980 212046 152992
rect 277946 152980 277952 152992
rect 212040 152952 277952 152980
rect 212040 152940 212046 152952
rect 277946 152940 277952 152952
rect 278004 152940 278010 152992
rect 373258 152940 373264 152992
rect 373316 152980 373322 152992
rect 452654 152980 452660 152992
rect 373316 152952 452660 152980
rect 373316 152940 373322 152952
rect 452654 152940 452660 152952
rect 452712 152940 452718 152992
rect 56410 152872 56416 152924
rect 56468 152912 56474 152924
rect 128354 152912 128360 152924
rect 56468 152884 128360 152912
rect 56468 152872 56474 152884
rect 128354 152872 128360 152884
rect 128412 152872 128418 152924
rect 216122 152872 216128 152924
rect 216180 152912 216186 152924
rect 280246 152912 280252 152924
rect 216180 152884 280252 152912
rect 216180 152872 216186 152884
rect 280246 152872 280252 152884
rect 280304 152872 280310 152924
rect 369118 152872 369124 152924
rect 369176 152912 369182 152924
rect 445754 152912 445760 152924
rect 369176 152884 445760 152912
rect 369176 152872 369182 152884
rect 445754 152872 445760 152884
rect 445812 152872 445818 152924
rect 54754 152804 54760 152856
rect 54812 152844 54818 152856
rect 125594 152844 125600 152856
rect 54812 152816 125600 152844
rect 54812 152804 54818 152816
rect 125594 152804 125600 152816
rect 125652 152804 125658 152856
rect 218882 152804 218888 152856
rect 218940 152844 218946 152856
rect 282914 152844 282920 152856
rect 218940 152816 282920 152844
rect 218940 152804 218946 152816
rect 282914 152804 282920 152816
rect 282972 152804 282978 152856
rect 363782 152804 363788 152856
rect 363840 152844 363846 152856
rect 440326 152844 440332 152856
rect 363840 152816 440332 152844
rect 363840 152804 363846 152816
rect 440326 152804 440332 152816
rect 440384 152804 440390 152856
rect 56042 152736 56048 152788
rect 56100 152776 56106 152788
rect 122834 152776 122840 152788
rect 56100 152748 122840 152776
rect 56100 152736 56106 152748
rect 122834 152736 122840 152748
rect 122892 152736 122898 152788
rect 209130 152736 209136 152788
rect 209188 152776 209194 152788
rect 268010 152776 268016 152788
rect 209188 152748 268016 152776
rect 209188 152736 209194 152748
rect 268010 152736 268016 152748
rect 268068 152736 268074 152788
rect 374638 152736 374644 152788
rect 374696 152776 374702 152788
rect 449894 152776 449900 152788
rect 374696 152748 449900 152776
rect 374696 152736 374702 152748
rect 449894 152736 449900 152748
rect 449952 152736 449958 152788
rect 54938 152668 54944 152720
rect 54996 152708 55002 152720
rect 120074 152708 120080 152720
rect 54996 152680 120080 152708
rect 54996 152668 55002 152680
rect 120074 152668 120080 152680
rect 120132 152668 120138 152720
rect 200758 152668 200764 152720
rect 200816 152708 200822 152720
rect 255958 152708 255964 152720
rect 200816 152680 255964 152708
rect 200816 152668 200822 152680
rect 255958 152668 255964 152680
rect 256016 152668 256022 152720
rect 365162 152668 365168 152720
rect 365220 152708 365226 152720
rect 434806 152708 434812 152720
rect 365220 152680 434812 152708
rect 365220 152668 365226 152680
rect 434806 152668 434812 152680
rect 434864 152668 434870 152720
rect 53466 152600 53472 152652
rect 53524 152640 53530 152652
rect 117498 152640 117504 152652
rect 53524 152612 117504 152640
rect 53524 152600 53530 152612
rect 117498 152600 117504 152612
rect 117556 152600 117562 152652
rect 183462 152600 183468 152652
rect 183520 152640 183526 152652
rect 197354 152640 197360 152652
rect 183520 152612 197360 152640
rect 183520 152600 183526 152612
rect 197354 152600 197360 152612
rect 197412 152600 197418 152652
rect 216030 152600 216036 152652
rect 216088 152640 216094 152652
rect 265066 152640 265072 152652
rect 216088 152612 265072 152640
rect 216088 152600 216094 152612
rect 265066 152600 265072 152612
rect 265124 152600 265130 152652
rect 343542 152600 343548 152652
rect 343600 152640 343606 152652
rect 357618 152640 357624 152652
rect 343600 152612 357624 152640
rect 343600 152600 343606 152612
rect 357618 152600 357624 152612
rect 357676 152600 357682 152652
rect 371970 152600 371976 152652
rect 372028 152640 372034 152652
rect 437474 152640 437480 152652
rect 372028 152612 437480 152640
rect 372028 152600 372034 152612
rect 437474 152600 437480 152612
rect 437532 152600 437538 152652
rect 503622 152600 503628 152652
rect 503680 152640 503686 152652
rect 517606 152640 517612 152652
rect 503680 152612 517612 152640
rect 503680 152600 503686 152612
rect 517606 152600 517612 152612
rect 517664 152600 517670 152652
rect 51994 152532 52000 152584
rect 52052 152572 52058 152584
rect 113174 152572 113180 152584
rect 52052 152544 113180 152572
rect 52052 152532 52058 152544
rect 113174 152532 113180 152544
rect 113232 152532 113238 152584
rect 204898 152532 204904 152584
rect 204956 152572 204962 152584
rect 253566 152572 253572 152584
rect 204956 152544 253572 152572
rect 204956 152532 204962 152544
rect 253566 152532 253572 152544
rect 253624 152532 253630 152584
rect 370682 152532 370688 152584
rect 370740 152572 370746 152584
rect 433334 152572 433340 152584
rect 370740 152544 433340 152572
rect 370740 152532 370746 152544
rect 433334 152532 433340 152544
rect 433392 152532 433398 152584
rect 55858 152464 55864 152516
rect 55916 152504 55922 152516
rect 115934 152504 115940 152516
rect 55916 152476 115940 152504
rect 55916 152464 55922 152476
rect 115934 152464 115940 152476
rect 115992 152464 115998 152516
rect 183462 152464 183468 152516
rect 183520 152504 183526 152516
rect 200114 152504 200120 152516
rect 183520 152476 200120 152504
rect 183520 152464 183526 152476
rect 200114 152464 200120 152476
rect 200172 152464 200178 152516
rect 213178 152464 213184 152516
rect 213236 152504 213242 152516
rect 258258 152504 258264 152516
rect 213236 152476 258264 152504
rect 213236 152464 213242 152476
rect 258258 152464 258264 152476
rect 258316 152464 258322 152516
rect 343542 152464 343548 152516
rect 343600 152504 343606 152516
rect 359458 152504 359464 152516
rect 343600 152476 359464 152504
rect 343600 152464 343606 152476
rect 359458 152464 359464 152476
rect 359516 152464 359522 152516
rect 376202 152464 376208 152516
rect 376260 152504 376266 152516
rect 415670 152504 415676 152516
rect 376260 152476 415676 152504
rect 376260 152464 376266 152476
rect 415670 152464 415676 152476
rect 415728 152464 415734 152516
rect 503622 152464 503628 152516
rect 503680 152504 503686 152516
rect 517882 152504 517888 152516
rect 503680 152476 517888 152504
rect 503680 152464 503686 152476
rect 517882 152464 517888 152476
rect 517940 152464 517946 152516
rect 50890 152396 50896 152448
rect 50948 152436 50954 152448
rect 103514 152436 103520 152448
rect 50948 152408 103520 152436
rect 50948 152396 50954 152408
rect 103514 152396 103520 152408
rect 103572 152396 103578 152448
rect 214558 152396 214564 152448
rect 214616 152436 214622 152448
rect 250254 152436 250260 152448
rect 214616 152408 250260 152436
rect 214616 152396 214622 152408
rect 250254 152396 250260 152408
rect 250312 152396 250318 152448
rect 374730 152396 374736 152448
rect 374788 152436 374794 152448
rect 413094 152436 413100 152448
rect 374788 152408 413100 152436
rect 374788 152396 374794 152408
rect 413094 152396 413100 152408
rect 413152 152396 413158 152448
rect 49234 152328 49240 152380
rect 49292 152368 49298 152380
rect 89714 152368 89720 152380
rect 49292 152340 89720 152368
rect 49292 152328 49298 152340
rect 89714 152328 89720 152340
rect 89772 152328 89778 152380
rect 97258 152328 97264 152380
rect 97316 152368 97322 152380
rect 100754 152368 100760 152380
rect 97316 152340 100760 152368
rect 97316 152328 97322 152340
rect 100754 152328 100760 152340
rect 100812 152328 100818 152380
rect 218790 152328 218796 152380
rect 218848 152368 218854 152380
rect 247126 152368 247132 152380
rect 218848 152340 247132 152368
rect 218848 152328 218854 152340
rect 247126 152328 247132 152340
rect 247184 152328 247190 152380
rect 372062 152328 372068 152380
rect 372120 152368 372126 152380
rect 409874 152368 409880 152380
rect 372120 152340 409880 152368
rect 372120 152328 372126 152340
rect 409874 152328 409880 152340
rect 409932 152328 409938 152380
rect 55030 152260 55036 152312
rect 55088 152300 55094 152312
rect 88334 152300 88340 152312
rect 55088 152272 88340 152300
rect 55088 152260 55094 152272
rect 88334 152260 88340 152272
rect 88392 152260 88398 152312
rect 378870 152260 378876 152312
rect 378928 152300 378934 152312
rect 407114 152300 407120 152312
rect 378928 152272 407120 152300
rect 378928 152260 378934 152272
rect 407114 152260 407120 152272
rect 407172 152260 407178 152312
rect 98638 151852 98644 151904
rect 98696 151892 98702 151904
rect 104894 151892 104900 151904
rect 98696 151864 104900 151892
rect 98696 151852 98702 151864
rect 104894 151852 104900 151864
rect 104952 151852 104958 151904
rect 212258 151784 212264 151836
rect 212316 151824 212322 151836
rect 219434 151824 219440 151836
rect 212316 151796 219440 151824
rect 212316 151784 212322 151796
rect 219434 151784 219440 151796
rect 219492 151784 219498 151836
rect 55674 151716 55680 151768
rect 55732 151756 55738 151768
rect 57790 151756 57796 151768
rect 55732 151728 57796 151756
rect 55732 151716 55738 151728
rect 57790 151716 57796 151728
rect 57848 151756 57854 151768
rect 117406 151756 117412 151768
rect 57848 151728 117412 151756
rect 57848 151716 57854 151728
rect 117406 151716 117412 151728
rect 117464 151716 117470 151768
rect 212074 151716 212080 151768
rect 212132 151756 212138 151768
rect 320174 151756 320180 151768
rect 212132 151728 320180 151756
rect 212132 151716 212138 151728
rect 320174 151716 320180 151728
rect 320232 151716 320238 151768
rect 375926 151716 375932 151768
rect 375984 151756 375990 151768
rect 436186 151756 436192 151768
rect 375984 151728 436192 151756
rect 375984 151716 375990 151728
rect 436186 151716 436192 151728
rect 436244 151716 436250 151768
rect 53650 151648 53656 151700
rect 53708 151688 53714 151700
rect 110414 151688 110420 151700
rect 53708 151660 110420 151688
rect 53708 151648 53714 151660
rect 110414 151648 110420 151660
rect 110472 151648 110478 151700
rect 219434 151648 219440 151700
rect 219492 151688 219498 151700
rect 219802 151688 219808 151700
rect 219492 151660 219808 151688
rect 219492 151648 219498 151660
rect 219802 151648 219808 151660
rect 219860 151688 219866 151700
rect 267734 151688 267740 151700
rect 219860 151660 267740 151688
rect 219860 151648 219866 151660
rect 267734 151648 267740 151660
rect 267792 151648 267798 151700
rect 277394 151648 277400 151700
rect 277452 151688 277458 151700
rect 278038 151688 278044 151700
rect 277452 151660 278044 151688
rect 277452 151648 277458 151660
rect 278038 151648 278044 151660
rect 278096 151688 278102 151700
rect 356974 151688 356980 151700
rect 278096 151660 356980 151688
rect 278096 151648 278102 151660
rect 356974 151648 356980 151660
rect 357032 151648 357038 151700
rect 379238 151648 379244 151700
rect 379296 151688 379302 151700
rect 426526 151688 426532 151700
rect 379296 151660 426532 151688
rect 379296 151648 379302 151660
rect 426526 151648 426532 151660
rect 426584 151648 426590 151700
rect 54386 151580 54392 151632
rect 54444 151620 54450 151632
rect 54938 151620 54944 151632
rect 54444 151592 54944 151620
rect 54444 151580 54450 151592
rect 54938 151580 54944 151592
rect 54996 151620 55002 151632
rect 97994 151620 98000 151632
rect 54996 151592 98000 151620
rect 54996 151580 55002 151592
rect 97994 151580 98000 151592
rect 98052 151580 98058 151632
rect 219894 151580 219900 151632
rect 219952 151620 219958 151632
rect 266354 151620 266360 151632
rect 219952 151592 266360 151620
rect 219952 151580 219958 151592
rect 266354 151580 266360 151592
rect 266412 151580 266418 151632
rect 375834 151580 375840 151632
rect 375892 151620 375898 151632
rect 375892 151592 380204 151620
rect 375892 151580 375898 151592
rect 218606 151512 218612 151564
rect 218664 151552 218670 151564
rect 219250 151552 219256 151564
rect 218664 151524 219256 151552
rect 218664 151512 218670 151524
rect 219250 151512 219256 151524
rect 219308 151552 219314 151564
rect 264974 151552 264980 151564
rect 219308 151524 264980 151552
rect 219308 151512 219314 151524
rect 264974 151512 264980 151524
rect 265032 151512 265038 151564
rect 376386 151512 376392 151564
rect 376444 151552 376450 151564
rect 380066 151552 380072 151564
rect 376444 151524 380072 151552
rect 376444 151512 376450 151524
rect 380066 151512 380072 151524
rect 380124 151512 380130 151564
rect 380176 151552 380204 151592
rect 380802 151580 380808 151632
rect 380860 151620 380866 151632
rect 427814 151620 427820 151632
rect 380860 151592 427820 151620
rect 380860 151580 380866 151592
rect 427814 151580 427820 151592
rect 427872 151580 427878 151632
rect 422294 151552 422300 151564
rect 380176 151524 422300 151552
rect 422294 151512 422300 151524
rect 422352 151512 422358 151564
rect 216398 151444 216404 151496
rect 216456 151484 216462 151496
rect 262214 151484 262220 151496
rect 216456 151456 262220 151484
rect 216456 151444 216462 151456
rect 262214 151444 262220 151456
rect 262272 151444 262278 151496
rect 425054 151484 425060 151496
rect 379808 151456 425060 151484
rect 53098 151376 53104 151428
rect 53156 151416 53162 151428
rect 57054 151416 57060 151428
rect 53156 151388 57060 151416
rect 53156 151376 53162 151388
rect 57054 151376 57060 151388
rect 57112 151416 57118 151428
rect 96614 151416 96620 151428
rect 57112 151388 96620 151416
rect 57112 151376 57118 151388
rect 96614 151376 96620 151388
rect 96672 151376 96678 151428
rect 214926 151376 214932 151428
rect 214984 151416 214990 151428
rect 259454 151416 259460 151428
rect 214984 151388 259460 151416
rect 214984 151376 214990 151388
rect 259454 151376 259460 151388
rect 259512 151376 259518 151428
rect 379808 151360 379836 151456
rect 425054 151444 425060 151456
rect 425112 151444 425118 151496
rect 420914 151416 420920 151428
rect 379900 151388 420920 151416
rect 59998 151308 60004 151360
rect 60056 151348 60062 151360
rect 106366 151348 106372 151360
rect 60056 151320 106372 151348
rect 60056 151308 60062 151320
rect 106366 151308 106372 151320
rect 106424 151308 106430 151360
rect 216214 151308 216220 151360
rect 216272 151348 216278 151360
rect 261202 151348 261208 151360
rect 216272 151320 261208 151348
rect 216272 151308 216278 151320
rect 261202 151308 261208 151320
rect 261260 151308 261266 151360
rect 379514 151308 379520 151360
rect 379572 151348 379578 151360
rect 379790 151348 379796 151360
rect 379572 151320 379796 151348
rect 379572 151308 379578 151320
rect 379790 151308 379796 151320
rect 379848 151308 379854 151360
rect 52822 151240 52828 151292
rect 52880 151280 52886 151292
rect 54846 151280 54852 151292
rect 52880 151252 54852 151280
rect 52880 151240 52886 151252
rect 54846 151240 54852 151252
rect 54904 151280 54910 151292
rect 100846 151280 100852 151292
rect 54904 151252 100852 151280
rect 54904 151240 54910 151252
rect 100846 151240 100852 151252
rect 100904 151240 100910 151292
rect 219618 151240 219624 151292
rect 219676 151280 219682 151292
rect 263594 151280 263600 151292
rect 219676 151252 263600 151280
rect 219676 151240 219682 151252
rect 263594 151240 263600 151252
rect 263652 151240 263658 151292
rect 376294 151240 376300 151292
rect 376352 151280 376358 151292
rect 379900 151280 379928 151388
rect 420914 151376 420920 151388
rect 420972 151376 420978 151428
rect 380158 151308 380164 151360
rect 380216 151348 380222 151360
rect 418246 151348 418252 151360
rect 380216 151320 418252 151348
rect 380216 151308 380222 151320
rect 418246 151308 418252 151320
rect 418304 151308 418310 151360
rect 376352 151252 379928 151280
rect 376352 151240 376358 151252
rect 380066 151240 380072 151292
rect 380124 151280 380130 151292
rect 418154 151280 418160 151292
rect 380124 151252 418160 151280
rect 380124 151240 380130 151252
rect 418154 151240 418160 151252
rect 418212 151240 418218 151292
rect 59262 151172 59268 151224
rect 59320 151212 59326 151224
rect 106274 151212 106280 151224
rect 59320 151184 106280 151212
rect 59320 151172 59326 151184
rect 106274 151172 106280 151184
rect 106332 151172 106338 151224
rect 217134 151172 217140 151224
rect 217192 151212 217198 151224
rect 258074 151212 258080 151224
rect 217192 151184 258080 151212
rect 217192 151172 217198 151184
rect 258074 151172 258080 151184
rect 258132 151172 258138 151224
rect 379698 151172 379704 151224
rect 379756 151212 379762 151224
rect 423674 151212 423680 151224
rect 379756 151184 423680 151212
rect 379756 151172 379762 151184
rect 423674 151172 423680 151184
rect 423732 151172 423738 151224
rect 49050 151104 49056 151156
rect 49108 151144 49114 151156
rect 55030 151144 55036 151156
rect 49108 151116 55036 151144
rect 49108 151104 49114 151116
rect 55030 151104 55036 151116
rect 55088 151144 55094 151156
rect 109126 151144 109132 151156
rect 55088 151116 109132 151144
rect 55088 151104 55094 151116
rect 109126 151104 109132 151116
rect 109184 151104 109190 151156
rect 219158 151104 219164 151156
rect 219216 151144 219222 151156
rect 219802 151144 219808 151156
rect 219216 151116 219808 151144
rect 219216 151104 219222 151116
rect 219802 151104 219808 151116
rect 219860 151144 219866 151156
rect 266446 151144 266452 151156
rect 219860 151116 266452 151144
rect 219860 151104 219866 151116
rect 266446 151104 266452 151116
rect 266504 151104 266510 151156
rect 373166 151104 373172 151156
rect 373224 151144 373230 151156
rect 375282 151144 375288 151156
rect 373224 151116 375288 151144
rect 373224 151104 373230 151116
rect 375282 151104 375288 151116
rect 375340 151144 375346 151156
rect 430574 151144 430580 151156
rect 375340 151116 430580 151144
rect 375340 151104 375346 151116
rect 430574 151104 430580 151116
rect 430632 151104 430638 151156
rect 46474 151036 46480 151088
rect 46532 151076 46538 151088
rect 51902 151076 51908 151088
rect 46532 151048 51908 151076
rect 46532 151036 46538 151048
rect 51902 151036 51908 151048
rect 51960 151076 51966 151088
rect 111794 151076 111800 151088
rect 51960 151048 111800 151076
rect 51960 151036 51966 151048
rect 111794 151036 111800 151048
rect 111852 151036 111858 151088
rect 213270 151036 213276 151088
rect 213328 151076 213334 151088
rect 216490 151076 216496 151088
rect 213328 151048 216496 151076
rect 213328 151036 213334 151048
rect 216490 151036 216496 151048
rect 216548 151076 216554 151088
rect 271874 151076 271880 151088
rect 216548 151048 271880 151076
rect 216548 151036 216554 151048
rect 271874 151036 271880 151048
rect 271932 151036 271938 151088
rect 372430 151036 372436 151088
rect 372488 151076 372494 151088
rect 374454 151076 374460 151088
rect 372488 151048 374460 151076
rect 372488 151036 372494 151048
rect 374454 151036 374460 151048
rect 374512 151076 374518 151088
rect 433978 151076 433984 151088
rect 374512 151048 433984 151076
rect 374512 151036 374518 151048
rect 433978 151036 433984 151048
rect 434036 151036 434042 151088
rect 218514 150968 218520 151020
rect 218572 151008 218578 151020
rect 218882 151008 218888 151020
rect 218572 150980 218888 151008
rect 218572 150968 218578 150980
rect 218882 150968 218888 150980
rect 218940 151008 218946 151020
rect 259546 151008 259552 151020
rect 218940 150980 259552 151008
rect 218940 150968 218946 150980
rect 259546 150968 259552 150980
rect 259604 150968 259610 151020
rect 379330 150968 379336 151020
rect 379388 151008 379394 151020
rect 419534 151008 419540 151020
rect 379388 150980 419540 151008
rect 379388 150968 379394 150980
rect 419534 150968 419540 150980
rect 419592 150968 419598 151020
rect 374546 150900 374552 150952
rect 374604 150940 374610 150952
rect 396074 150940 396080 150952
rect 374604 150912 396080 150940
rect 374604 150900 374610 150912
rect 396074 150900 396080 150912
rect 396132 150900 396138 150952
rect 375190 150832 375196 150884
rect 375248 150872 375254 150884
rect 396166 150872 396172 150884
rect 375248 150844 396172 150872
rect 375248 150832 375254 150844
rect 396166 150832 396172 150844
rect 396224 150832 396230 150884
rect 374914 150764 374920 150816
rect 374972 150804 374978 150816
rect 380158 150804 380164 150816
rect 374972 150776 380164 150804
rect 374972 150764 374978 150776
rect 380158 150764 380164 150776
rect 380216 150764 380222 150816
rect 58618 150628 58624 150680
rect 58676 150668 58682 150680
rect 59998 150668 60004 150680
rect 58676 150640 60004 150668
rect 58676 150628 58682 150640
rect 59998 150628 60004 150640
rect 60056 150628 60062 150680
rect 375926 150492 375932 150544
rect 375984 150532 375990 150544
rect 376662 150532 376668 150544
rect 375984 150504 376668 150532
rect 375984 150492 375990 150504
rect 376662 150492 376668 150504
rect 376720 150492 376726 150544
rect 377030 150492 377036 150544
rect 377088 150532 377094 150544
rect 379698 150532 379704 150544
rect 377088 150504 379704 150532
rect 377088 150492 377094 150504
rect 379698 150492 379704 150504
rect 379756 150492 379762 150544
rect 214190 150424 214196 150476
rect 214248 150464 214254 150476
rect 214926 150464 214932 150476
rect 214248 150436 214932 150464
rect 214248 150424 214254 150436
rect 214926 150424 214932 150436
rect 214984 150424 214990 150476
rect 216122 150424 216128 150476
rect 216180 150464 216186 150476
rect 216398 150464 216404 150476
rect 216180 150436 216404 150464
rect 216180 150424 216186 150436
rect 216398 150424 216404 150436
rect 216456 150424 216462 150476
rect 376202 150424 376208 150476
rect 376260 150464 376266 150476
rect 376386 150464 376392 150476
rect 376260 150436 376392 150464
rect 376260 150424 376266 150436
rect 376386 150424 376392 150436
rect 376444 150424 376450 150476
rect 379238 150424 379244 150476
rect 379296 150464 379302 150476
rect 379422 150464 379428 150476
rect 379296 150436 379428 150464
rect 379296 150424 379302 150436
rect 379422 150424 379428 150436
rect 379480 150424 379486 150476
rect 47946 150356 47952 150408
rect 48004 150396 48010 150408
rect 58618 150396 58624 150408
rect 48004 150368 58624 150396
rect 48004 150356 48010 150368
rect 58618 150356 58624 150368
rect 58676 150396 58682 150408
rect 59262 150396 59268 150408
rect 58676 150368 59268 150396
rect 58676 150356 58682 150368
rect 59262 150356 59268 150368
rect 59320 150356 59326 150408
rect 214742 150356 214748 150408
rect 214800 150396 214806 150408
rect 236086 150396 236092 150408
rect 214800 150368 236092 150396
rect 214800 150356 214806 150368
rect 236086 150356 236092 150368
rect 236144 150356 236150 150408
rect 212810 149676 212816 149728
rect 212868 149716 212874 149728
rect 214926 149716 214932 149728
rect 212868 149688 214932 149716
rect 212868 149676 212874 149688
rect 214926 149676 214932 149688
rect 214984 149716 214990 149728
rect 270494 149716 270500 149728
rect 214984 149688 270500 149716
rect 214984 149676 214990 149688
rect 270494 149676 270500 149688
rect 270552 149676 270558 149728
rect 52178 147064 52184 147076
rect 52104 147036 52184 147064
rect 52104 146872 52132 147036
rect 52178 147024 52184 147036
rect 52236 147024 52242 147076
rect 52086 146820 52092 146872
rect 52144 146820 52150 146872
rect 51810 146752 51816 146804
rect 51868 146792 51874 146804
rect 52178 146792 52184 146804
rect 51868 146764 52184 146792
rect 51868 146752 51874 146764
rect 52178 146752 52184 146764
rect 52236 146752 52242 146804
rect 213288 133912 213684 133940
rect 54478 133832 54484 133884
rect 54536 133872 54542 133884
rect 117314 133872 117320 133884
rect 54536 133844 117320 133872
rect 54536 133832 54542 133844
rect 117314 133832 117320 133844
rect 117372 133832 117378 133884
rect 212350 133832 212356 133884
rect 212408 133872 212414 133884
rect 213288 133872 213316 133912
rect 212408 133844 213316 133872
rect 212408 133832 212414 133844
rect 213362 133832 213368 133884
rect 213420 133872 213426 133884
rect 213546 133872 213552 133884
rect 213420 133844 213552 133872
rect 213420 133832 213426 133844
rect 213546 133832 213552 133844
rect 213604 133832 213610 133884
rect 213656 133872 213684 133912
rect 273254 133872 273260 133884
rect 213656 133844 273260 133872
rect 273254 133832 273260 133844
rect 273312 133832 273318 133884
rect 378594 133832 378600 133884
rect 378652 133872 378658 133884
rect 379146 133872 379152 133884
rect 378652 133844 379152 133872
rect 378652 133832 378658 133844
rect 379146 133832 379152 133844
rect 379204 133832 379210 133884
rect 436094 133872 436100 133884
rect 379256 133844 436100 133872
rect 48038 133764 48044 133816
rect 48096 133804 48102 133816
rect 53650 133804 53656 133816
rect 48096 133776 53656 133804
rect 48096 133764 48102 133776
rect 53650 133764 53656 133776
rect 53708 133764 53714 133816
rect 56318 133764 56324 133816
rect 56376 133804 56382 133816
rect 56962 133804 56968 133816
rect 56376 133776 56968 133804
rect 56376 133764 56382 133776
rect 56962 133764 56968 133776
rect 57020 133804 57026 133816
rect 103606 133804 103612 133816
rect 57020 133776 103612 133804
rect 57020 133764 57026 133776
rect 103606 133764 103612 133776
rect 103664 133764 103670 133816
rect 47762 133696 47768 133748
rect 47820 133736 47826 133748
rect 53466 133736 53472 133748
rect 47820 133708 53472 133736
rect 47820 133696 47826 133708
rect 53466 133696 53472 133708
rect 53524 133736 53530 133748
rect 213564 133736 213592 133832
rect 214650 133764 214656 133816
rect 214708 133804 214714 133816
rect 240134 133804 240140 133816
rect 214708 133776 240140 133804
rect 214708 133764 214714 133776
rect 240134 133764 240140 133776
rect 240192 133764 240198 133816
rect 375006 133764 375012 133816
rect 375064 133804 375070 133816
rect 379256 133804 379284 133844
rect 436094 133832 436100 133844
rect 436152 133832 436158 133884
rect 375064 133776 379284 133804
rect 375064 133764 375070 133776
rect 379330 133764 379336 133816
rect 379388 133804 379394 133816
rect 434714 133804 434720 133816
rect 379388 133776 434720 133804
rect 379388 133764 379394 133776
rect 434714 133764 434720 133776
rect 434772 133764 434778 133816
rect 238754 133736 238760 133748
rect 53524 133708 60734 133736
rect 213564 133708 238760 133736
rect 53524 133696 53530 133708
rect 46290 133628 46296 133680
rect 46348 133668 46354 133680
rect 46348 133640 51074 133668
rect 46348 133628 46354 133640
rect 51046 133464 51074 133640
rect 54478 133492 54484 133544
rect 54536 133532 54542 133544
rect 54754 133532 54760 133544
rect 54536 133504 54760 133532
rect 54536 133492 54542 133504
rect 54754 133492 54760 133504
rect 54812 133492 54818 133544
rect 60706 133532 60734 133708
rect 238754 133696 238760 133708
rect 238812 133696 238818 133748
rect 379146 133696 379152 133748
rect 379204 133736 379210 133748
rect 412726 133736 412732 133748
rect 379204 133708 412732 133736
rect 379204 133696 379210 133708
rect 412726 133696 412732 133708
rect 412784 133696 412790 133748
rect 210786 133628 210792 133680
rect 210844 133668 210850 133680
rect 215018 133668 215024 133680
rect 210844 133640 215024 133668
rect 210844 133628 210850 133640
rect 215018 133628 215024 133640
rect 215076 133628 215082 133680
rect 374822 133628 374828 133680
rect 374880 133668 374886 133680
rect 401594 133668 401600 133680
rect 374880 133640 401600 133668
rect 374880 133628 374886 133640
rect 401594 133628 401600 133640
rect 401652 133628 401658 133680
rect 372430 133560 372436 133612
rect 372488 133600 372494 133612
rect 373442 133600 373448 133612
rect 372488 133572 373448 133600
rect 372488 133560 372494 133572
rect 373442 133560 373448 133572
rect 373500 133600 373506 133612
rect 400214 133600 400220 133612
rect 373500 133572 400220 133600
rect 373500 133560 373506 133572
rect 400214 133560 400220 133572
rect 400272 133560 400278 133612
rect 80054 133532 80060 133544
rect 60706 133504 80060 133532
rect 80054 133492 80060 133504
rect 80112 133492 80118 133544
rect 377674 133492 377680 133544
rect 377732 133532 377738 133544
rect 379330 133532 379336 133544
rect 377732 133504 379336 133532
rect 377732 133492 377738 133504
rect 379330 133492 379336 133504
rect 379388 133492 379394 133544
rect 51902 133464 51908 133476
rect 51046 133436 51908 133464
rect 51902 133424 51908 133436
rect 51960 133464 51966 133476
rect 78674 133464 78680 133476
rect 51960 133436 78680 133464
rect 51960 133424 51966 133436
rect 78674 133424 78680 133436
rect 78732 133424 78738 133476
rect 213638 133424 213644 133476
rect 213696 133464 213702 133476
rect 214650 133464 214656 133476
rect 213696 133436 214656 133464
rect 213696 133424 213702 133436
rect 214650 133424 214656 133436
rect 214708 133424 214714 133476
rect 53650 133356 53656 133408
rect 53708 133396 53714 133408
rect 81434 133396 81440 133408
rect 53708 133368 81440 133396
rect 53708 133356 53714 133368
rect 81434 133356 81440 133368
rect 81492 133356 81498 133408
rect 46198 133288 46204 133340
rect 46256 133328 46262 133340
rect 59906 133328 59912 133340
rect 46256 133300 59912 133328
rect 46256 133288 46262 133300
rect 59906 133288 59912 133300
rect 59964 133328 59970 133340
rect 109034 133328 109040 133340
rect 59964 133300 109040 133328
rect 59964 133288 59970 133300
rect 109034 133288 109040 133300
rect 109092 133288 109098 133340
rect 51534 133220 51540 133272
rect 51592 133260 51598 133272
rect 53558 133260 53564 133272
rect 51592 133232 53564 133260
rect 51592 133220 51598 133232
rect 53558 133220 53564 133232
rect 53616 133260 53622 133272
rect 114554 133260 114560 133272
rect 53616 133232 114560 133260
rect 53616 133220 53622 133232
rect 114554 133220 114560 133232
rect 114612 133220 114618 133272
rect 215018 133220 215024 133272
rect 215076 133260 215082 133272
rect 241514 133260 241520 133272
rect 215076 133232 241520 133260
rect 215076 133220 215082 133232
rect 241514 133220 241520 133232
rect 241572 133220 241578 133272
rect 53282 133152 53288 133204
rect 53340 133192 53346 133204
rect 114646 133192 114652 133204
rect 53340 133164 114652 133192
rect 53340 133152 53346 133164
rect 114646 133152 114652 133164
rect 114704 133152 114710 133204
rect 216490 133152 216496 133204
rect 216548 133192 216554 133204
rect 278038 133192 278044 133204
rect 216548 133164 278044 133192
rect 216548 133152 216554 133164
rect 278038 133152 278044 133164
rect 278096 133152 278102 133204
rect 280062 133152 280068 133204
rect 280120 133192 280126 133204
rect 306374 133192 306380 133204
rect 280120 133164 306380 133192
rect 280120 133152 280126 133164
rect 306374 133152 306380 133164
rect 306432 133152 306438 133204
rect 373534 133152 373540 133204
rect 373592 133192 373598 133204
rect 375190 133192 375196 133204
rect 373592 133164 375196 133192
rect 373592 133152 373598 133164
rect 375190 133152 375196 133164
rect 375248 133192 375254 133204
rect 398834 133192 398840 133204
rect 375248 133164 398840 133192
rect 375248 133152 375254 133164
rect 398834 133152 398840 133164
rect 398892 133152 398898 133204
rect 373902 132472 373908 132524
rect 373960 132512 373966 132524
rect 374822 132512 374828 132524
rect 373960 132484 374828 132512
rect 373960 132472 373966 132484
rect 374822 132472 374828 132484
rect 374880 132472 374886 132524
rect 306374 131792 306380 131844
rect 306432 131832 306438 131844
rect 356974 131832 356980 131844
rect 306432 131804 356980 131832
rect 306432 131792 306438 131804
rect 356974 131792 356980 131804
rect 357032 131792 357038 131844
rect 356974 131588 356980 131640
rect 357032 131628 357038 131640
rect 357710 131628 357716 131640
rect 357032 131600 357716 131628
rect 357032 131588 357038 131600
rect 357710 131588 357716 131600
rect 357768 131588 357774 131640
rect 191742 131112 191748 131164
rect 191800 131152 191806 131164
rect 197998 131152 198004 131164
rect 191800 131124 198004 131152
rect 191800 131112 191806 131124
rect 197998 131112 198004 131124
rect 198056 131112 198062 131164
rect 213546 131112 213552 131164
rect 213604 131152 213610 131164
rect 274726 131152 274732 131164
rect 213604 131124 274732 131152
rect 213604 131112 213610 131124
rect 274726 131112 274732 131124
rect 274784 131112 274790 131164
rect 55766 131044 55772 131096
rect 55824 131084 55830 131096
rect 56410 131084 56416 131096
rect 55824 131056 56416 131084
rect 55824 131044 55830 131056
rect 56410 131044 56416 131056
rect 56468 131044 56474 131096
rect 56962 131044 56968 131096
rect 57020 131084 57026 131096
rect 57238 131084 57244 131096
rect 57020 131056 57244 131084
rect 57020 131044 57026 131056
rect 57238 131044 57244 131056
rect 57296 131044 57302 131096
rect 59814 131044 59820 131096
rect 59872 131084 59878 131096
rect 93854 131084 93860 131096
rect 59872 131056 93860 131084
rect 59872 131044 59878 131056
rect 93854 131044 93860 131056
rect 93912 131044 93918 131096
rect 179046 131044 179052 131096
rect 179104 131084 179110 131096
rect 196710 131084 196716 131096
rect 179104 131056 196716 131084
rect 179104 131044 179110 131056
rect 196710 131044 196716 131056
rect 196768 131044 196774 131096
rect 216030 131044 216036 131096
rect 216088 131084 216094 131096
rect 218974 131084 218980 131096
rect 216088 131056 218980 131084
rect 216088 131044 216094 131056
rect 218974 131044 218980 131056
rect 219032 131084 219038 131096
rect 245654 131084 245660 131096
rect 219032 131056 245660 131084
rect 219032 131044 219038 131056
rect 245654 131044 245660 131056
rect 245712 131044 245718 131096
rect 338482 131044 338488 131096
rect 338540 131084 338546 131096
rect 360194 131084 360200 131096
rect 338540 131056 360200 131084
rect 338540 131044 338546 131056
rect 360194 131044 360200 131056
rect 360252 131044 360258 131096
rect 379974 131044 379980 131096
rect 380032 131084 380038 131096
rect 415394 131084 415400 131096
rect 380032 131056 415400 131084
rect 380032 131044 380038 131056
rect 415394 131044 415400 131056
rect 415452 131044 415458 131096
rect 57256 131016 57284 131044
rect 91094 131016 91100 131028
rect 57256 130988 91100 131016
rect 91094 130976 91100 130988
rect 91152 130976 91158 131028
rect 179782 130976 179788 131028
rect 179840 131016 179846 131028
rect 196618 131016 196624 131028
rect 179840 130988 196624 131016
rect 179840 130976 179846 130988
rect 196618 130976 196624 130988
rect 196676 130976 196682 131028
rect 219526 130976 219532 131028
rect 219584 131016 219590 131028
rect 253934 131016 253940 131028
rect 219584 130988 253940 131016
rect 219584 130976 219590 130988
rect 253934 130976 253940 130988
rect 253992 130976 253998 131028
rect 340598 130976 340604 131028
rect 340656 131016 340662 131028
rect 356882 131016 356888 131028
rect 340656 130988 356888 131016
rect 340656 130976 340662 130988
rect 356882 130976 356888 130988
rect 356940 130976 356946 131028
rect 377582 130976 377588 131028
rect 377640 131016 377646 131028
rect 411254 131016 411260 131028
rect 377640 130988 411260 131016
rect 377640 130976 377646 130988
rect 411254 130976 411260 130988
rect 411312 130976 411318 131028
rect 500218 130976 500224 131028
rect 500276 131016 500282 131028
rect 517698 131016 517704 131028
rect 500276 130988 517704 131016
rect 500276 130976 500282 130988
rect 517698 130976 517704 130988
rect 517756 130976 517762 131028
rect 56410 130908 56416 130960
rect 56468 130948 56474 130960
rect 88426 130948 88432 130960
rect 56468 130920 88432 130948
rect 56468 130908 56474 130920
rect 88426 130908 88432 130920
rect 88484 130908 88490 130960
rect 218330 130908 218336 130960
rect 218388 130948 218394 130960
rect 218790 130948 218796 130960
rect 218388 130920 218796 130948
rect 218388 130908 218394 130920
rect 218790 130908 218796 130920
rect 218848 130948 218854 130960
rect 252554 130948 252560 130960
rect 218848 130920 252560 130948
rect 218848 130908 218854 130920
rect 252554 130908 252560 130920
rect 252612 130908 252618 130960
rect 379330 130908 379336 130960
rect 379388 130948 379394 130960
rect 411346 130948 411352 130960
rect 379388 130920 411352 130948
rect 379388 130908 379394 130920
rect 411346 130908 411352 130920
rect 411404 130908 411410 130960
rect 498746 130908 498752 130960
rect 498804 130948 498810 130960
rect 517790 130948 517796 130960
rect 498804 130920 517796 130948
rect 498804 130908 498810 130920
rect 517790 130908 517796 130920
rect 517848 130908 517854 130960
rect 51718 130840 51724 130892
rect 51776 130880 51782 130892
rect 84194 130880 84200 130892
rect 51776 130852 84200 130880
rect 51776 130840 51782 130852
rect 84194 130840 84200 130852
rect 84252 130840 84258 130892
rect 217594 130840 217600 130892
rect 217652 130880 217658 130892
rect 251266 130880 251272 130892
rect 217652 130852 251272 130880
rect 217652 130840 217658 130852
rect 251266 130840 251272 130852
rect 251324 130840 251330 130892
rect 377674 130840 377680 130892
rect 377732 130880 377738 130892
rect 409966 130880 409972 130892
rect 377732 130852 409972 130880
rect 377732 130840 377738 130852
rect 409966 130840 409972 130852
rect 410024 130840 410030 130892
rect 53374 130772 53380 130824
rect 53432 130812 53438 130824
rect 85574 130812 85580 130824
rect 53432 130784 85580 130812
rect 53432 130772 53438 130784
rect 85574 130772 85580 130784
rect 85632 130772 85638 130824
rect 218974 130772 218980 130824
rect 219032 130812 219038 130824
rect 219342 130812 219348 130824
rect 219032 130784 219348 130812
rect 219032 130772 219038 130784
rect 219342 130772 219348 130784
rect 219400 130812 219406 130824
rect 251174 130812 251180 130824
rect 219400 130784 251180 130812
rect 219400 130772 219406 130784
rect 251174 130772 251180 130784
rect 251232 130772 251238 130824
rect 376478 130772 376484 130824
rect 376536 130812 376542 130824
rect 376536 130784 379652 130812
rect 376536 130772 376542 130784
rect 48958 130704 48964 130756
rect 49016 130744 49022 130756
rect 55950 130744 55956 130756
rect 49016 130716 55956 130744
rect 49016 130704 49022 130716
rect 55950 130704 55956 130716
rect 56008 130704 56014 130756
rect 59078 130704 59084 130756
rect 59136 130744 59142 130756
rect 91186 130744 91192 130756
rect 59136 130716 91192 130744
rect 59136 130704 59142 130716
rect 91186 130704 91192 130716
rect 91244 130704 91250 130756
rect 216306 130704 216312 130756
rect 216364 130744 216370 130756
rect 248414 130744 248420 130756
rect 216364 130716 248420 130744
rect 216364 130704 216370 130716
rect 248414 130704 248420 130716
rect 248472 130704 248478 130756
rect 379624 130744 379652 130784
rect 380066 130772 380072 130824
rect 380124 130812 380130 130824
rect 408494 130812 408500 130824
rect 380124 130784 408500 130812
rect 380124 130772 380130 130784
rect 408494 130772 408500 130784
rect 408552 130772 408558 130824
rect 402974 130744 402980 130756
rect 379624 130716 402980 130744
rect 402974 130704 402980 130716
rect 403032 130704 403038 130756
rect 58894 130636 58900 130688
rect 58952 130676 58958 130688
rect 59262 130676 59268 130688
rect 58952 130648 59268 130676
rect 58952 130636 58958 130648
rect 59262 130636 59268 130648
rect 59320 130676 59326 130688
rect 89806 130676 89812 130688
rect 59320 130648 89812 130676
rect 59320 130636 59326 130648
rect 89806 130636 89812 130648
rect 89864 130636 89870 130688
rect 214650 130636 214656 130688
rect 214708 130676 214714 130688
rect 244366 130676 244372 130688
rect 214708 130648 244372 130676
rect 214708 130636 214714 130648
rect 244366 130636 244372 130648
rect 244424 130636 244430 130688
rect 379054 130636 379060 130688
rect 379112 130676 379118 130688
rect 405734 130676 405740 130688
rect 379112 130648 405740 130676
rect 379112 130636 379118 130648
rect 405734 130636 405740 130648
rect 405792 130636 405798 130688
rect 55950 130568 55956 130620
rect 56008 130608 56014 130620
rect 82814 130608 82820 130620
rect 56008 130580 82820 130608
rect 56008 130568 56014 130580
rect 82814 130568 82820 130580
rect 82872 130568 82878 130620
rect 214466 130568 214472 130620
rect 214524 130608 214530 130620
rect 242894 130608 242900 130620
rect 214524 130580 242900 130608
rect 214524 130568 214530 130580
rect 242894 130568 242900 130580
rect 242952 130568 242958 130620
rect 378686 130568 378692 130620
rect 378744 130608 378750 130620
rect 379330 130608 379336 130620
rect 378744 130580 379336 130608
rect 378744 130568 378750 130580
rect 379330 130568 379336 130580
rect 379388 130568 379394 130620
rect 380250 130568 380256 130620
rect 380308 130608 380314 130620
rect 403066 130608 403072 130620
rect 380308 130580 403072 130608
rect 380308 130568 380314 130580
rect 403066 130568 403072 130580
rect 403124 130568 403130 130620
rect 54478 130500 54484 130552
rect 54536 130540 54542 130552
rect 84286 130540 84292 130552
rect 54536 130512 84292 130540
rect 54536 130500 54542 130512
rect 84286 130500 84292 130512
rect 84344 130500 84350 130552
rect 212994 130500 213000 130552
rect 213052 130540 213058 130552
rect 219066 130540 219072 130552
rect 213052 130512 219072 130540
rect 213052 130500 213058 130512
rect 219066 130500 219072 130512
rect 219124 130540 219130 130552
rect 247034 130540 247040 130552
rect 219124 130512 247040 130540
rect 219124 130500 219130 130512
rect 247034 130500 247040 130512
rect 247092 130500 247098 130552
rect 375742 130500 375748 130552
rect 375800 130540 375806 130552
rect 380066 130540 380072 130552
rect 375800 130512 380072 130540
rect 375800 130500 375806 130512
rect 380066 130500 380072 130512
rect 380124 130500 380130 130552
rect 380158 130500 380164 130552
rect 380216 130540 380222 130552
rect 407206 130540 407212 130552
rect 380216 130512 407212 130540
rect 380216 130500 380222 130512
rect 407206 130500 407212 130512
rect 407264 130500 407270 130552
rect 55858 130432 55864 130484
rect 55916 130472 55922 130484
rect 86954 130472 86960 130484
rect 55916 130444 86960 130472
rect 55916 130432 55922 130444
rect 86954 130432 86960 130444
rect 87012 130432 87018 130484
rect 183462 130432 183468 130484
rect 183520 130472 183526 130484
rect 197446 130472 197452 130484
rect 183520 130444 197452 130472
rect 183520 130432 183526 130444
rect 197446 130432 197452 130444
rect 197504 130432 197510 130484
rect 214282 130432 214288 130484
rect 214340 130472 214346 130484
rect 214650 130472 214656 130484
rect 214340 130444 214656 130472
rect 214340 130432 214346 130444
rect 214650 130432 214656 130444
rect 214708 130432 214714 130484
rect 215938 130432 215944 130484
rect 215996 130472 216002 130484
rect 244274 130472 244280 130484
rect 215996 130444 244280 130472
rect 215996 130432 216002 130444
rect 244274 130432 244280 130444
rect 244332 130432 244338 130484
rect 278682 130432 278688 130484
rect 278740 130472 278746 130484
rect 302234 130472 302240 130484
rect 278740 130444 302240 130472
rect 278740 130432 278746 130444
rect 302234 130432 302240 130444
rect 302292 130432 302298 130484
rect 343542 130432 343548 130484
rect 343600 130472 343606 130484
rect 357434 130472 357440 130484
rect 343600 130444 357440 130472
rect 343600 130432 343606 130444
rect 357434 130432 357440 130444
rect 357492 130432 357498 130484
rect 373718 130432 373724 130484
rect 373776 130472 373782 130484
rect 374730 130472 374736 130484
rect 373776 130444 374736 130472
rect 373776 130432 373782 130444
rect 374730 130432 374736 130444
rect 374788 130472 374794 130484
rect 404354 130472 404360 130484
rect 374788 130444 404360 130472
rect 374788 130432 374794 130444
rect 404354 130432 404360 130444
rect 404412 130432 404418 130484
rect 440142 130432 440148 130484
rect 440200 130472 440206 130484
rect 466454 130472 466460 130484
rect 440200 130444 466460 130472
rect 440200 130432 440206 130444
rect 466454 130432 466460 130444
rect 466512 130432 466518 130484
rect 503622 130432 503628 130484
rect 503680 130472 503686 130484
rect 517606 130472 517612 130484
rect 503680 130444 517612 130472
rect 503680 130432 503686 130444
rect 517606 130432 517612 130444
rect 517664 130432 517670 130484
rect 48866 130364 48872 130416
rect 48924 130404 48930 130416
rect 59170 130404 59176 130416
rect 48924 130376 59176 130404
rect 48924 130364 48930 130376
rect 59170 130364 59176 130376
rect 59228 130404 59234 130416
rect 92474 130404 92480 130416
rect 59228 130376 92480 130404
rect 59228 130364 59234 130376
rect 92474 130364 92480 130376
rect 92532 130364 92538 130416
rect 197998 130364 198004 130416
rect 198056 130404 198062 130416
rect 214558 130404 214564 130416
rect 198056 130376 214564 130404
rect 198056 130364 198062 130376
rect 214558 130364 214564 130376
rect 214616 130364 214622 130416
rect 215662 130364 215668 130416
rect 215720 130404 215726 130416
rect 218514 130404 218520 130416
rect 215720 130376 218520 130404
rect 215720 130364 215726 130376
rect 218514 130364 218520 130376
rect 218572 130404 218578 130416
rect 256694 130404 256700 130416
rect 218572 130376 256700 130404
rect 218572 130364 218578 130376
rect 256694 130364 256700 130376
rect 256752 130364 256758 130416
rect 274726 130364 274732 130416
rect 274784 130404 274790 130416
rect 300762 130404 300768 130416
rect 274784 130376 300768 130404
rect 274784 130364 274790 130376
rect 300762 130364 300768 130376
rect 300820 130364 300826 130416
rect 351730 130364 351736 130416
rect 351788 130404 351794 130416
rect 358078 130404 358084 130416
rect 351788 130376 358084 130404
rect 351788 130364 351794 130376
rect 358078 130364 358084 130376
rect 358136 130404 358142 130416
rect 358722 130404 358728 130416
rect 358136 130376 358728 130404
rect 358136 130364 358142 130376
rect 358722 130364 358728 130376
rect 358780 130404 358786 130416
rect 510614 130404 510620 130416
rect 358780 130376 510620 130404
rect 358780 130364 358786 130376
rect 510614 130364 510620 130376
rect 510672 130364 510678 130416
rect 48130 130296 48136 130348
rect 48188 130336 48194 130348
rect 51626 130336 51632 130348
rect 48188 130308 51632 130336
rect 48188 130296 48194 130308
rect 51626 130296 51632 130308
rect 51684 130336 51690 130348
rect 77294 130336 77300 130348
rect 51684 130308 77300 130336
rect 51684 130296 51690 130308
rect 77294 130296 77300 130308
rect 77352 130296 77358 130348
rect 215754 130296 215760 130348
rect 215812 130336 215818 130348
rect 235994 130336 236000 130348
rect 215812 130308 236000 130336
rect 215812 130296 215818 130308
rect 235994 130296 236000 130308
rect 236052 130296 236058 130348
rect 372522 130296 372528 130348
rect 372580 130336 372586 130348
rect 374822 130336 374828 130348
rect 372580 130308 374828 130336
rect 372580 130296 372586 130308
rect 374822 130296 374828 130308
rect 374880 130336 374886 130348
rect 397454 130336 397460 130348
rect 374880 130308 397460 130336
rect 374880 130296 374886 130308
rect 397454 130296 397460 130308
rect 397512 130296 397518 130348
rect 46566 130228 46572 130280
rect 46624 130268 46630 130280
rect 54202 130268 54208 130280
rect 46624 130240 54208 130268
rect 46624 130228 46630 130240
rect 54202 130228 54208 130240
rect 54260 130268 54266 130280
rect 76006 130268 76012 130280
rect 54260 130240 76012 130268
rect 54260 130228 54266 130240
rect 76006 130228 76012 130240
rect 76064 130228 76070 130280
rect 218606 130228 218612 130280
rect 218664 130268 218670 130280
rect 236086 130268 236092 130280
rect 218664 130240 236092 130268
rect 218664 130228 218670 130240
rect 236086 130228 236092 130240
rect 236144 130228 236150 130280
rect 378686 130228 378692 130280
rect 378744 130268 378750 130280
rect 396166 130268 396172 130280
rect 378744 130240 396172 130268
rect 378744 130228 378750 130240
rect 396166 130228 396172 130240
rect 396224 130228 396230 130280
rect 48222 130160 48228 130212
rect 48280 130200 48286 130212
rect 54662 130200 54668 130212
rect 48280 130172 54668 130200
rect 48280 130160 48286 130172
rect 54662 130160 54668 130172
rect 54720 130200 54726 130212
rect 75914 130200 75920 130212
rect 54720 130172 75920 130200
rect 54720 130160 54726 130172
rect 75914 130160 75920 130172
rect 75972 130160 75978 130212
rect 217226 130160 217232 130212
rect 217284 130200 217290 130212
rect 255314 130200 255320 130212
rect 217284 130172 255320 130200
rect 217284 130160 217290 130172
rect 255314 130160 255320 130172
rect 255372 130160 255378 130212
rect 378594 130160 378600 130212
rect 378652 130200 378658 130212
rect 396074 130200 396080 130212
rect 378652 130172 396080 130200
rect 378652 130160 378658 130172
rect 396074 130160 396080 130172
rect 396132 130160 396138 130212
rect 375098 130092 375104 130144
rect 375156 130132 375162 130144
rect 378870 130132 378876 130144
rect 375156 130104 378876 130132
rect 375156 130092 375162 130104
rect 378870 130092 378876 130104
rect 378928 130132 378934 130144
rect 380158 130132 380164 130144
rect 378928 130104 380164 130132
rect 378928 130092 378934 130104
rect 380158 130092 380164 130104
rect 380216 130092 380222 130144
rect 375650 130024 375656 130076
rect 375708 130064 375714 130076
rect 380250 130064 380256 130076
rect 375708 130036 380256 130064
rect 375708 130024 375714 130036
rect 380250 130024 380256 130036
rect 380308 130024 380314 130076
rect 376386 129820 376392 129872
rect 376444 129860 376450 129872
rect 379054 129860 379060 129872
rect 376444 129832 379060 129860
rect 376444 129820 376450 129832
rect 379054 129820 379060 129832
rect 379112 129820 379118 129872
rect 219526 129752 219532 129804
rect 219584 129792 219590 129804
rect 219710 129792 219716 129804
rect 219584 129764 219716 129792
rect 219584 129752 219590 129764
rect 219710 129752 219716 129764
rect 219768 129752 219774 129804
rect 374638 129752 374644 129804
rect 374696 129792 374702 129804
rect 375650 129792 375656 129804
rect 374696 129764 375656 129792
rect 374696 129752 374702 129764
rect 375650 129752 375656 129764
rect 375708 129752 375714 129804
rect 375926 129752 375932 129804
rect 375984 129792 375990 129804
rect 376478 129792 376484 129804
rect 375984 129764 376484 129792
rect 375984 129752 375990 129764
rect 376478 129752 376484 129764
rect 376536 129752 376542 129804
rect 378962 129752 378968 129804
rect 379020 129792 379026 129804
rect 379974 129792 379980 129804
rect 379020 129764 379980 129792
rect 379020 129752 379026 129764
rect 379974 129752 379980 129764
rect 380032 129752 380038 129804
rect 50522 129684 50528 129736
rect 50580 129724 50586 129736
rect 54478 129724 54484 129736
rect 50580 129696 54484 129724
rect 50580 129684 50586 129696
rect 54478 129684 54484 129696
rect 54536 129684 54542 129736
rect 54570 129684 54576 129736
rect 54628 129724 54634 129736
rect 55858 129724 55864 129736
rect 54628 129696 55864 129724
rect 54628 129684 54634 129696
rect 55858 129684 55864 129696
rect 55916 129684 55922 129736
rect 213454 129684 213460 129736
rect 213512 129724 213518 129736
rect 215938 129724 215944 129736
rect 213512 129696 215944 129724
rect 213512 129684 213518 129696
rect 215938 129684 215944 129696
rect 215996 129684 216002 129736
rect 300762 129684 300768 129736
rect 300820 129724 300826 129736
rect 356606 129724 356612 129736
rect 300820 129696 356612 129724
rect 300820 129684 300826 129696
rect 356606 129684 356612 129696
rect 356664 129684 356670 129736
rect 373074 129684 373080 129736
rect 373132 129724 373138 129736
rect 376110 129724 376116 129736
rect 373132 129696 376116 129724
rect 373132 129684 373138 129696
rect 376110 129684 376116 129696
rect 376168 129724 376174 129736
rect 376570 129724 376576 129736
rect 376168 129696 376576 129724
rect 376168 129684 376174 129696
rect 376570 129684 376576 129696
rect 376628 129684 376634 129736
rect 466454 129684 466460 129736
rect 466512 129724 466518 129736
rect 516594 129724 516600 129736
rect 466512 129696 516600 129724
rect 466512 129684 466518 129696
rect 516594 129684 516600 129696
rect 516652 129684 516658 129736
rect 212902 129616 212908 129668
rect 212960 129656 212966 129668
rect 215846 129656 215852 129668
rect 212960 129628 215852 129656
rect 212960 129616 212966 129628
rect 215846 129616 215852 129628
rect 215904 129616 215910 129668
rect 302234 129004 302240 129056
rect 302292 129044 302298 129056
rect 356790 129044 356796 129056
rect 302292 129016 356796 129044
rect 302292 129004 302298 129016
rect 356790 129004 356796 129016
rect 356848 129044 356854 129056
rect 357526 129044 357532 129056
rect 356848 129016 357532 129044
rect 356848 129004 356854 129016
rect 357526 129004 357532 129016
rect 357584 129004 357590 129056
rect 375742 128664 375748 128716
rect 375800 128704 375806 128716
rect 376570 128704 376576 128716
rect 375800 128676 376576 128704
rect 375800 128664 375806 128676
rect 376570 128664 376576 128676
rect 376628 128664 376634 128716
rect 215846 127576 215852 127628
rect 215904 127616 215910 127628
rect 215904 127588 215984 127616
rect 215904 127576 215910 127588
rect 215956 127424 215984 127588
rect 215938 127372 215944 127424
rect 215996 127372 216002 127424
rect 2958 120028 2964 120080
rect 3016 120068 3022 120080
rect 11698 120068 11704 120080
rect 3016 120040 11704 120068
rect 3016 120028 3022 120040
rect 11698 120028 11704 120040
rect 11756 120028 11762 120080
rect 57790 81404 57796 81456
rect 57848 81444 57854 81456
rect 59354 81444 59360 81456
rect 57848 81416 59360 81444
rect 57848 81404 57854 81416
rect 59354 81404 59360 81416
rect 59412 81404 59418 81456
rect 366450 55156 366456 55208
rect 366508 55196 366514 55208
rect 376938 55196 376944 55208
rect 366508 55168 376944 55196
rect 366508 55156 366514 55168
rect 376938 55156 376944 55168
rect 376996 55156 377002 55208
rect 214558 53116 214564 53168
rect 214616 53156 214622 53168
rect 215202 53156 215208 53168
rect 214616 53128 215208 53156
rect 214616 53116 214622 53128
rect 215202 53116 215208 53128
rect 215260 53156 215266 53168
rect 216674 53156 216680 53168
rect 215260 53128 216680 53156
rect 215260 53116 215266 53128
rect 216674 53116 216680 53128
rect 216732 53116 216738 53168
rect 358722 53048 358728 53100
rect 358780 53088 358786 53100
rect 376938 53088 376944 53100
rect 358780 53060 376944 53088
rect 358780 53048 358786 53060
rect 376938 53048 376944 53060
rect 376996 53048 377002 53100
rect 358078 52436 358084 52488
rect 358136 52476 358142 52488
rect 358722 52476 358728 52488
rect 358136 52448 358728 52476
rect 358136 52436 358142 52448
rect 358722 52436 358728 52448
rect 358780 52436 358786 52488
rect 378686 44684 378692 44736
rect 378744 44724 378750 44736
rect 397086 44724 397092 44736
rect 378744 44696 397092 44724
rect 378744 44684 378750 44696
rect 397086 44684 397092 44696
rect 397144 44684 397150 44736
rect 378594 44616 378600 44668
rect 378652 44656 378658 44668
rect 396074 44656 396080 44668
rect 378652 44628 396080 44656
rect 378652 44616 378658 44628
rect 396074 44616 396080 44628
rect 396132 44616 396138 44668
rect 218606 44548 218612 44600
rect 218664 44588 218670 44600
rect 235994 44588 236000 44600
rect 218664 44560 236000 44588
rect 218664 44548 218670 44560
rect 235994 44548 236000 44560
rect 236052 44548 236058 44600
rect 374638 44548 374644 44600
rect 374696 44588 374702 44600
rect 403066 44588 403072 44600
rect 374696 44560 403072 44588
rect 374696 44548 374702 44560
rect 403066 44548 403072 44560
rect 403124 44548 403130 44600
rect 54202 44480 54208 44532
rect 54260 44520 54266 44532
rect 77110 44520 77116 44532
rect 54260 44492 77116 44520
rect 54260 44480 54266 44492
rect 77110 44480 77116 44492
rect 77168 44480 77174 44532
rect 215754 44480 215760 44532
rect 215812 44520 215818 44532
rect 237098 44520 237104 44532
rect 215812 44492 237104 44520
rect 215812 44480 215818 44492
rect 237098 44480 237104 44492
rect 237156 44480 237162 44532
rect 379882 44480 379888 44532
rect 379940 44520 379946 44532
rect 414566 44520 414572 44532
rect 379940 44492 414572 44520
rect 379940 44480 379946 44492
rect 414566 44480 414572 44492
rect 414624 44480 414630 44532
rect 55950 44412 55956 44464
rect 56008 44452 56014 44464
rect 83090 44452 83096 44464
rect 56008 44424 83096 44452
rect 56008 44412 56014 44424
rect 83090 44412 83096 44424
rect 83148 44412 83154 44464
rect 214466 44412 214472 44464
rect 214524 44452 214530 44464
rect 243078 44452 243084 44464
rect 214524 44424 243084 44452
rect 214524 44412 214530 44424
rect 243078 44412 243084 44424
rect 243136 44412 243142 44464
rect 377214 44412 377220 44464
rect 377272 44452 377278 44464
rect 416958 44452 416964 44464
rect 377272 44424 416964 44452
rect 377272 44412 377278 44424
rect 416958 44412 416964 44424
rect 417016 44412 417022 44464
rect 58986 44344 58992 44396
rect 59044 44384 59050 44396
rect 101766 44384 101772 44396
rect 59044 44356 101772 44384
rect 59044 44344 59050 44356
rect 101766 44344 101772 44356
rect 101824 44344 101830 44396
rect 217226 44344 217232 44396
rect 217284 44384 217290 44396
rect 255866 44384 255872 44396
rect 217284 44356 255872 44384
rect 217284 44344 217290 44356
rect 255866 44344 255872 44356
rect 255924 44344 255930 44396
rect 376202 44344 376208 44396
rect 376260 44384 376266 44396
rect 419442 44384 419448 44396
rect 376260 44356 419448 44384
rect 376260 44344 376266 44356
rect 419442 44344 419448 44356
rect 419500 44344 419506 44396
rect 54846 44276 54852 44328
rect 54904 44316 54910 44328
rect 100754 44316 100760 44328
rect 54904 44288 100760 44316
rect 54904 44276 54910 44288
rect 100754 44276 100760 44288
rect 100812 44276 100818 44328
rect 218514 44276 218520 44328
rect 218572 44316 218578 44328
rect 256970 44316 256976 44328
rect 218572 44288 256976 44316
rect 218572 44276 218578 44288
rect 256970 44276 256976 44288
rect 257028 44276 257034 44328
rect 374914 44276 374920 44328
rect 374972 44316 374978 44328
rect 418154 44316 418160 44328
rect 374972 44288 418160 44316
rect 374972 44276 374978 44288
rect 418154 44276 418160 44288
rect 418212 44276 418218 44328
rect 54386 44208 54392 44260
rect 54444 44248 54450 44260
rect 143534 44248 143540 44260
rect 54444 44220 143540 44248
rect 54444 44208 54450 44220
rect 143534 44208 143540 44220
rect 143592 44208 143598 44260
rect 217134 44208 217140 44260
rect 217192 44248 217198 44260
rect 258074 44248 258080 44260
rect 217192 44220 258080 44248
rect 217192 44208 217198 44220
rect 258074 44208 258080 44220
rect 258132 44208 258138 44260
rect 379698 44208 379704 44260
rect 379756 44248 379762 44260
rect 423950 44248 423956 44260
rect 379756 44220 423956 44248
rect 379756 44208 379762 44220
rect 423950 44208 423956 44220
rect 424008 44208 424014 44260
rect 51442 44140 51448 44192
rect 51500 44180 51506 44192
rect 145926 44180 145932 44192
rect 51500 44152 145932 44180
rect 51500 44140 51506 44152
rect 145926 44140 145932 44152
rect 145984 44140 145990 44192
rect 216122 44140 216128 44192
rect 216180 44180 216186 44192
rect 262858 44180 262864 44192
rect 216180 44152 262864 44180
rect 216180 44140 216186 44152
rect 262858 44140 262864 44152
rect 262916 44140 262922 44192
rect 363598 44140 363604 44192
rect 363656 44180 363662 44192
rect 410702 44180 410708 44192
rect 363656 44152 410708 44180
rect 363656 44140 363662 44152
rect 410702 44140 410708 44152
rect 410760 44140 410766 44192
rect 57882 44072 57888 44124
rect 57940 44112 57946 44124
rect 215202 44112 215208 44124
rect 57940 44084 215208 44112
rect 57940 44072 57946 44084
rect 215202 44072 215208 44084
rect 215260 44112 215266 44124
rect 358078 44112 358084 44124
rect 215260 44084 358084 44112
rect 215260 44072 215266 44084
rect 358078 44072 358084 44084
rect 358136 44072 358142 44124
rect 376386 44072 376392 44124
rect 376444 44112 376450 44124
rect 406470 44112 406476 44124
rect 376444 44084 406476 44112
rect 376444 44072 376450 44084
rect 406470 44072 406476 44084
rect 406528 44072 406534 44124
rect 3418 44004 3424 44056
rect 3476 44044 3482 44056
rect 7558 44044 7564 44056
rect 3476 44016 7564 44044
rect 3476 44004 3482 44016
rect 7558 44004 7564 44016
rect 7616 44004 7622 44056
rect 54478 44004 54484 44056
rect 54536 44044 54542 44056
rect 84194 44044 84200 44056
rect 54536 44016 84200 44044
rect 54536 44004 54542 44016
rect 84194 44004 84200 44016
rect 84252 44004 84258 44056
rect 215846 44004 215852 44056
rect 215904 44044 215910 44056
rect 244274 44044 244280 44056
rect 215904 44016 244280 44044
rect 215904 44004 215910 44016
rect 244274 44004 244280 44016
rect 244332 44004 244338 44056
rect 374730 44004 374736 44056
rect 374788 44044 374794 44056
rect 405458 44044 405464 44056
rect 374788 44016 405464 44044
rect 374788 44004 374794 44016
rect 405458 44004 405464 44016
rect 405516 44004 405522 44056
rect 59814 43936 59820 43988
rect 59872 43976 59878 43988
rect 94498 43976 94504 43988
rect 59872 43948 94504 43976
rect 59872 43936 59878 43948
rect 94498 43936 94504 43948
rect 94556 43936 94562 43988
rect 218882 43936 218888 43988
rect 218940 43976 218946 43988
rect 259454 43976 259460 43988
rect 218940 43948 259460 43976
rect 218940 43936 218946 43948
rect 259454 43936 259460 43948
rect 259512 43936 259518 43988
rect 379238 43936 379244 43988
rect 379296 43976 379302 43988
rect 420638 43976 420644 43988
rect 379296 43948 420644 43976
rect 379296 43936 379302 43948
rect 420638 43936 420644 43948
rect 420696 43936 420702 43988
rect 57054 43868 57060 43920
rect 57112 43908 57118 43920
rect 96982 43908 96988 43920
rect 57112 43880 96988 43908
rect 57112 43868 57118 43880
rect 96982 43868 96988 43880
rect 97040 43868 97046 43920
rect 219618 43868 219624 43920
rect 219676 43908 219682 43920
rect 263870 43908 263876 43920
rect 219676 43880 263876 43908
rect 219676 43868 219682 43880
rect 263870 43868 263876 43880
rect 263928 43868 263934 43920
rect 376294 43868 376300 43920
rect 376352 43908 376358 43920
rect 421742 43908 421748 43920
rect 376352 43880 421748 43908
rect 376352 43868 376358 43880
rect 421742 43868 421748 43880
rect 421800 43868 421806 43920
rect 54938 43800 54944 43852
rect 54996 43840 55002 43852
rect 98086 43840 98092 43852
rect 54996 43812 98092 43840
rect 54996 43800 55002 43812
rect 98086 43800 98092 43812
rect 98144 43800 98150 43852
rect 216214 43800 216220 43852
rect 216272 43840 216278 43852
rect 261754 43840 261760 43852
rect 216272 43812 261760 43840
rect 216272 43800 216278 43812
rect 261754 43800 261760 43812
rect 261812 43800 261818 43852
rect 379790 43800 379796 43852
rect 379848 43840 379854 43852
rect 425238 43840 425244 43852
rect 379848 43812 425244 43840
rect 379848 43800 379854 43812
rect 425238 43800 425244 43812
rect 425296 43800 425302 43852
rect 56042 43732 56048 43784
rect 56100 43772 56106 43784
rect 102778 43772 102784 43784
rect 56100 43744 102784 43772
rect 56100 43732 56106 43744
rect 102778 43732 102784 43744
rect 102836 43732 102842 43784
rect 214190 43732 214196 43784
rect 214248 43772 214254 43784
rect 260650 43772 260656 43784
rect 214248 43744 260656 43772
rect 214248 43732 214254 43744
rect 260650 43732 260656 43744
rect 260708 43732 260714 43784
rect 279234 43732 279240 43784
rect 279292 43772 279298 43784
rect 356974 43772 356980 43784
rect 279292 43744 356980 43772
rect 279292 43732 279298 43744
rect 356974 43732 356980 43744
rect 357032 43732 357038 43784
rect 375834 43732 375840 43784
rect 375892 43772 375898 43784
rect 422846 43772 422852 43784
rect 375892 43744 422852 43772
rect 375892 43732 375898 43744
rect 422846 43732 422852 43744
rect 422904 43732 422910 43784
rect 56318 43664 56324 43716
rect 56376 43704 56382 43716
rect 103882 43704 103888 43716
rect 56376 43676 103888 43704
rect 56376 43664 56382 43676
rect 103882 43664 103888 43676
rect 103940 43664 103946 43716
rect 212442 43664 212448 43716
rect 212500 43704 212506 43716
rect 308490 43704 308496 43716
rect 212500 43676 308496 43704
rect 212500 43664 212506 43676
rect 308490 43664 308496 43676
rect 308548 43664 308554 43716
rect 356698 43664 356704 43716
rect 356756 43704 356762 43716
rect 425974 43704 425980 43716
rect 356756 43676 425980 43704
rect 356756 43664 356762 43676
rect 425974 43664 425980 43676
rect 426032 43664 426038 43716
rect 53282 43596 53288 43648
rect 53340 43636 53346 43648
rect 113266 43636 113272 43648
rect 53340 43608 113272 43636
rect 53340 43596 53346 43608
rect 113266 43596 113272 43608
rect 113324 43596 113330 43648
rect 213730 43596 213736 43648
rect 213788 43636 213794 43648
rect 315850 43636 315856 43648
rect 213788 43608 315856 43636
rect 213788 43596 213794 43608
rect 315850 43596 315856 43608
rect 315908 43596 315914 43648
rect 366358 43596 366364 43648
rect 366416 43636 366422 43648
rect 458450 43636 458456 43648
rect 366416 43608 458456 43636
rect 366416 43596 366422 43608
rect 458450 43596 458456 43608
rect 458508 43596 458514 43648
rect 42518 43528 42524 43580
rect 42576 43568 42582 43580
rect 115934 43568 115940 43580
rect 42576 43540 115940 43568
rect 42576 43528 42582 43540
rect 115934 43528 115940 43540
rect 115992 43528 115998 43580
rect 219250 43528 219256 43580
rect 219308 43568 219314 43580
rect 421006 43568 421012 43580
rect 219308 43540 421012 43568
rect 219308 43528 219314 43540
rect 421006 43528 421012 43540
rect 421064 43528 421070 43580
rect 56226 43460 56232 43512
rect 56284 43500 56290 43512
rect 158438 43500 158444 43512
rect 56284 43472 158444 43500
rect 56284 43460 56290 43472
rect 158438 43460 158444 43472
rect 158496 43460 158502 43512
rect 198642 43460 198648 43512
rect 198700 43500 198706 43512
rect 300854 43500 300860 43512
rect 198700 43472 300860 43500
rect 198700 43460 198706 43472
rect 300854 43460 300860 43472
rect 300912 43460 300918 43512
rect 358170 43460 358176 43512
rect 358228 43500 358234 43512
rect 455874 43500 455880 43512
rect 358228 43472 455880 43500
rect 358228 43460 358234 43472
rect 455874 43460 455880 43472
rect 455932 43460 455938 43512
rect 49602 43392 49608 43444
rect 49660 43432 49666 43444
rect 160830 43432 160836 43444
rect 49660 43404 160836 43432
rect 49660 43392 49666 43404
rect 160830 43392 160836 43404
rect 160888 43392 160894 43444
rect 218974 43392 218980 43444
rect 219032 43432 219038 43444
rect 428182 43432 428188 43444
rect 219032 43404 428188 43432
rect 219032 43392 219038 43404
rect 428182 43392 428188 43404
rect 428240 43392 428246 43444
rect 439222 43392 439228 43444
rect 439280 43432 439286 43444
rect 516594 43432 516600 43444
rect 439280 43404 516600 43432
rect 439280 43392 439286 43404
rect 516594 43392 516600 43404
rect 516652 43392 516658 43444
rect 378870 43324 378876 43376
rect 378928 43364 378934 43376
rect 407574 43364 407580 43376
rect 378928 43336 407580 43364
rect 378928 43324 378934 43336
rect 407574 43324 407580 43336
rect 407632 43324 407638 43376
rect 375926 43256 375932 43308
rect 375984 43296 375990 43308
rect 404170 43296 404176 43308
rect 375984 43268 404176 43296
rect 375984 43256 375990 43268
rect 404170 43256 404176 43268
rect 404228 43256 404234 43308
rect 57238 42780 57244 42832
rect 57296 42820 57302 42832
rect 57882 42820 57888 42832
rect 57296 42792 57888 42820
rect 57296 42780 57302 42792
rect 57882 42780 57888 42792
rect 57940 42780 57946 42832
rect 50982 42712 50988 42764
rect 51040 42752 51046 42764
rect 155954 42752 155960 42764
rect 51040 42724 155960 42752
rect 51040 42712 51046 42724
rect 155954 42712 155960 42724
rect 156012 42712 156018 42764
rect 183462 42712 183468 42764
rect 183520 42752 183526 42764
rect 197446 42752 197452 42764
rect 183520 42724 197452 42752
rect 183520 42712 183526 42724
rect 197446 42712 197452 42724
rect 197504 42712 197510 42764
rect 209590 42712 209596 42764
rect 209648 42752 209654 42764
rect 320910 42752 320916 42764
rect 209648 42724 320916 42752
rect 209648 42712 209654 42724
rect 320910 42712 320916 42724
rect 320968 42712 320974 42764
rect 343174 42712 343180 42764
rect 343232 42752 343238 42764
rect 357618 42752 357624 42764
rect 343232 42724 357624 42752
rect 343232 42712 343238 42724
rect 357618 42712 357624 42724
rect 357676 42712 357682 42764
rect 378502 42712 378508 42764
rect 378560 42752 378566 42764
rect 485958 42752 485964 42764
rect 378560 42724 485964 42752
rect 378560 42712 378566 42724
rect 485958 42712 485964 42724
rect 486016 42712 486022 42764
rect 503254 42712 503260 42764
rect 503312 42752 503318 42764
rect 517606 42752 517612 42764
rect 503312 42724 517612 42752
rect 503312 42712 503318 42724
rect 517606 42712 517612 42724
rect 517664 42712 517670 42764
rect 52270 42644 52276 42696
rect 52328 42684 52334 42696
rect 135898 42684 135904 42696
rect 52328 42656 135904 42684
rect 52328 42644 52334 42656
rect 135898 42644 135904 42656
rect 135956 42644 135962 42696
rect 183186 42644 183192 42696
rect 183244 42684 183250 42696
rect 197354 42684 197360 42696
rect 183244 42656 197360 42684
rect 183244 42644 183250 42656
rect 197354 42644 197360 42656
rect 197412 42644 197418 42696
rect 218238 42644 218244 42696
rect 218296 42684 218302 42696
rect 325878 42684 325884 42696
rect 218296 42656 325884 42684
rect 218296 42644 218302 42656
rect 325878 42644 325884 42656
rect 325936 42644 325942 42696
rect 343450 42644 343456 42696
rect 343508 42684 343514 42696
rect 357434 42684 357440 42696
rect 343508 42656 357440 42684
rect 343508 42644 343514 42656
rect 357434 42644 357440 42656
rect 357492 42644 357498 42696
rect 365070 42644 365076 42696
rect 365128 42684 365134 42696
rect 453390 42684 453396 42696
rect 365128 42656 453396 42684
rect 365128 42644 365134 42656
rect 453390 42644 453396 42656
rect 453448 42644 453454 42696
rect 503530 42644 503536 42696
rect 503588 42684 503594 42696
rect 517514 42684 517520 42696
rect 503588 42656 517520 42684
rect 503588 42644 503594 42656
rect 517514 42644 517520 42656
rect 517572 42644 517578 42696
rect 53742 42576 53748 42628
rect 53800 42616 53806 42628
rect 133414 42616 133420 42628
rect 53800 42588 133420 42616
rect 53800 42576 53806 42588
rect 133414 42576 133420 42588
rect 133472 42576 133478 42628
rect 216582 42576 216588 42628
rect 216640 42616 216646 42628
rect 318334 42616 318340 42628
rect 216640 42588 318340 42616
rect 216640 42576 216646 42588
rect 318334 42576 318340 42588
rect 318392 42576 318398 42628
rect 360930 42576 360936 42628
rect 360988 42616 360994 42628
rect 448238 42616 448244 42628
rect 360988 42588 448244 42616
rect 360988 42576 360994 42588
rect 448238 42576 448244 42588
rect 448296 42576 448302 42628
rect 56502 42508 56508 42560
rect 56560 42548 56566 42560
rect 128354 42548 128360 42560
rect 56560 42520 128360 42548
rect 56560 42508 56566 42520
rect 128354 42508 128360 42520
rect 128412 42508 128418 42560
rect 211062 42508 211068 42560
rect 211120 42548 211126 42560
rect 310974 42548 310980 42560
rect 211120 42520 310980 42548
rect 211120 42508 211126 42520
rect 310974 42508 310980 42520
rect 311032 42508 311038 42560
rect 364978 42508 364984 42560
rect 365036 42548 365042 42560
rect 445846 42548 445852 42560
rect 365036 42520 445852 42548
rect 365036 42508 365042 42520
rect 445846 42508 445852 42520
rect 445904 42508 445910 42560
rect 55122 42440 55128 42492
rect 55180 42480 55186 42492
rect 118234 42480 118240 42492
rect 55180 42452 118240 42480
rect 55180 42440 55186 42452
rect 118234 42440 118240 42452
rect 118292 42440 118298 42492
rect 213822 42440 213828 42492
rect 213880 42480 213886 42492
rect 313366 42480 313372 42492
rect 213880 42452 313372 42480
rect 213880 42440 213886 42452
rect 313366 42440 313372 42452
rect 313424 42440 313430 42492
rect 367738 42440 367744 42492
rect 367796 42480 367802 42492
rect 443454 42480 443460 42492
rect 367796 42452 443460 42480
rect 367796 42440 367802 42452
rect 443454 42440 443460 42452
rect 443512 42440 443518 42492
rect 52362 42372 52368 42424
rect 52420 42412 52426 42424
rect 113174 42412 113180 42424
rect 52420 42384 113180 42412
rect 52420 42372 52426 42384
rect 113174 42372 113180 42384
rect 113232 42372 113238 42424
rect 215110 42372 215116 42424
rect 215168 42412 215174 42424
rect 298462 42412 298468 42424
rect 215168 42384 298468 42412
rect 215168 42372 215174 42384
rect 298462 42372 298468 42384
rect 298520 42372 298526 42424
rect 361022 42372 361028 42424
rect 361080 42412 361086 42424
rect 435910 42412 435916 42424
rect 361080 42384 435916 42412
rect 361080 42372 361086 42384
rect 435910 42372 435916 42384
rect 435968 42372 435974 42424
rect 43990 42304 43996 42356
rect 44048 42344 44054 42356
rect 96246 42344 96252 42356
rect 44048 42316 96252 42344
rect 44048 42304 44054 42316
rect 96246 42304 96252 42316
rect 96304 42304 96310 42356
rect 209682 42304 209688 42356
rect 209740 42344 209746 42356
rect 293310 42344 293316 42356
rect 209740 42316 293316 42344
rect 209740 42304 209746 42316
rect 293310 42304 293316 42316
rect 293368 42304 293374 42356
rect 370498 42304 370504 42356
rect 370556 42344 370562 42356
rect 440878 42344 440884 42356
rect 370556 42316 440884 42344
rect 370556 42304 370562 42316
rect 440878 42304 440884 42316
rect 440936 42304 440942 42356
rect 59906 42236 59912 42288
rect 59964 42276 59970 42288
rect 108574 42276 108580 42288
rect 59964 42248 108580 42276
rect 59964 42236 59970 42248
rect 108574 42236 108580 42248
rect 108632 42236 108638 42288
rect 218422 42236 218428 42288
rect 218480 42276 218486 42288
rect 302510 42276 302516 42288
rect 218480 42248 302516 42276
rect 218480 42236 218486 42248
rect 302510 42236 302516 42248
rect 302568 42236 302574 42288
rect 371878 42236 371884 42288
rect 371936 42276 371942 42288
rect 438486 42276 438492 42288
rect 371936 42248 438492 42276
rect 371936 42236 371942 42248
rect 438486 42236 438492 42248
rect 438544 42236 438550 42288
rect 56134 42168 56140 42220
rect 56192 42208 56198 42220
rect 95878 42208 95884 42220
rect 56192 42180 95884 42208
rect 56192 42168 56198 42180
rect 95878 42168 95884 42180
rect 95936 42168 95942 42220
rect 211798 42168 211804 42220
rect 211856 42208 211862 42220
rect 276106 42208 276112 42220
rect 211856 42180 276112 42208
rect 211856 42168 211862 42180
rect 276106 42168 276112 42180
rect 276164 42168 276170 42220
rect 278314 42168 278320 42220
rect 278372 42208 278378 42220
rect 356790 42208 356796 42220
rect 278372 42180 356796 42208
rect 278372 42168 278378 42180
rect 356790 42168 356796 42180
rect 356848 42168 356854 42220
rect 378778 42168 378784 42220
rect 378836 42208 378842 42220
rect 430942 42208 430948 42220
rect 378836 42180 430948 42208
rect 378836 42168 378842 42180
rect 430942 42168 430948 42180
rect 431000 42168 431006 42220
rect 50154 42100 50160 42152
rect 50212 42140 50218 42152
rect 88334 42140 88340 42152
rect 50212 42112 88340 42140
rect 50212 42100 50218 42112
rect 88334 42100 88340 42112
rect 88392 42100 88398 42152
rect 218698 42100 218704 42152
rect 218756 42140 218762 42152
rect 268194 42140 268200 42152
rect 218756 42112 268200 42140
rect 218756 42100 218762 42112
rect 268194 42100 268200 42112
rect 268252 42100 268258 42152
rect 363690 42100 363696 42152
rect 363748 42140 363754 42152
rect 413646 42140 413652 42152
rect 363748 42112 413652 42140
rect 363748 42100 363754 42112
rect 413646 42100 413652 42112
rect 413704 42100 413710 42152
rect 54662 42032 54668 42084
rect 54720 42072 54726 42084
rect 76006 42072 76012 42084
rect 54720 42044 76012 42072
rect 54720 42032 54726 42044
rect 76006 42032 76012 42044
rect 76064 42032 76070 42084
rect 211890 42032 211896 42084
rect 211948 42072 211954 42084
rect 260926 42072 260932 42084
rect 211948 42044 260932 42072
rect 211948 42032 211954 42044
rect 260926 42032 260932 42044
rect 260984 42032 260990 42084
rect 379606 42032 379612 42084
rect 379664 42072 379670 42084
rect 427630 42072 427636 42084
rect 379664 42044 427636 42072
rect 379664 42032 379670 42044
rect 427630 42032 427636 42044
rect 427688 42032 427694 42084
rect 378962 41964 378968 42016
rect 379020 42004 379026 42016
rect 415486 42004 415492 42016
rect 379020 41976 415492 42004
rect 379020 41964 379026 41976
rect 415486 41964 415492 41976
rect 415544 41964 415550 42016
rect 52086 41352 52092 41404
rect 52144 41392 52150 41404
rect 115750 41392 115756 41404
rect 52144 41364 115756 41392
rect 52144 41352 52150 41364
rect 115750 41352 115756 41364
rect 115808 41352 115814 41404
rect 219986 41352 219992 41404
rect 220044 41392 220050 41404
rect 408310 41392 408316 41404
rect 220044 41364 408316 41392
rect 220044 41352 220050 41364
rect 408310 41352 408316 41364
rect 408368 41352 408374 41404
rect 57790 41284 57796 41336
rect 57848 41324 57854 41336
rect 119062 41324 119068 41336
rect 57848 41296 119068 41324
rect 57848 41284 57854 41296
rect 119062 41284 119068 41296
rect 119120 41284 119126 41336
rect 216490 41284 216496 41336
rect 216548 41324 216554 41336
rect 276934 41324 276940 41336
rect 216548 41296 276940 41324
rect 216548 41284 216554 41296
rect 276934 41284 276940 41296
rect 276992 41284 276998 41336
rect 376110 41284 376116 41336
rect 376168 41324 376174 41336
rect 429654 41324 429660 41336
rect 376168 41296 429660 41324
rect 376168 41284 376174 41296
rect 429654 41284 429660 41296
rect 429712 41284 429718 41336
rect 53558 41216 53564 41268
rect 53616 41256 53622 41268
rect 114186 41256 114192 41268
rect 53616 41228 114192 41256
rect 53616 41216 53622 41228
rect 114186 41216 114192 41228
rect 114244 41216 114250 41268
rect 214374 41216 214380 41268
rect 214432 41256 214438 41268
rect 273254 41256 273260 41268
rect 214432 41228 273260 41256
rect 214432 41216 214438 41228
rect 273254 41216 273260 41228
rect 273312 41216 273318 41268
rect 379422 41216 379428 41268
rect 379480 41256 379486 41268
rect 426434 41256 426440 41268
rect 379480 41228 426440 41256
rect 379480 41216 379486 41228
rect 426434 41216 426440 41228
rect 426492 41216 426498 41268
rect 42610 41148 42616 41200
rect 42668 41188 42674 41200
rect 93670 41188 93676 41200
rect 42668 41160 93676 41188
rect 42668 41148 42674 41160
rect 93670 41148 93676 41160
rect 93728 41148 93734 41200
rect 214926 41148 214932 41200
rect 214984 41188 214990 41200
rect 271230 41188 271236 41200
rect 214984 41160 271236 41188
rect 214984 41148 214990 41160
rect 271230 41148 271236 41160
rect 271288 41148 271294 41200
rect 379146 41148 379152 41200
rect 379204 41188 379210 41200
rect 413278 41188 413284 41200
rect 379204 41160 413284 41188
rect 379204 41148 379210 41160
rect 413278 41148 413284 41160
rect 413336 41148 413342 41200
rect 58618 41080 58624 41132
rect 58676 41120 58682 41132
rect 107010 41120 107016 41132
rect 58676 41092 107016 41120
rect 58676 41080 58682 41092
rect 107010 41080 107016 41092
rect 107068 41080 107074 41132
rect 212258 41080 212264 41132
rect 212316 41120 212322 41132
rect 268470 41120 268476 41132
rect 212316 41092 268476 41120
rect 212316 41080 212322 41092
rect 268470 41080 268476 41092
rect 268528 41080 268534 41132
rect 377674 41080 377680 41132
rect 377732 41120 377738 41132
rect 409966 41120 409972 41132
rect 377732 41092 409972 41120
rect 377732 41080 377738 41092
rect 409966 41080 409972 41092
rect 410024 41080 410030 41132
rect 59998 41012 60004 41064
rect 60056 41052 60062 41064
rect 106366 41052 106372 41064
rect 60056 41024 106372 41052
rect 60056 41012 60062 41024
rect 106366 41012 106372 41024
rect 106424 41012 106430 41064
rect 219342 41012 219348 41064
rect 219400 41052 219406 41064
rect 265158 41052 265164 41064
rect 219400 41024 265164 41052
rect 219400 41012 219406 41024
rect 265158 41012 265164 41024
rect 265216 41012 265222 41064
rect 373902 41012 373908 41064
rect 373960 41052 373966 41064
rect 401686 41052 401692 41064
rect 373960 41024 401692 41052
rect 373960 41012 373966 41024
rect 401686 41012 401692 41024
rect 401744 41012 401750 41064
rect 51718 40944 51724 40996
rect 51776 40984 51782 40996
rect 85390 40984 85396 40996
rect 51776 40956 85396 40984
rect 51776 40944 51782 40956
rect 85390 40944 85396 40956
rect 85448 40944 85454 40996
rect 218790 40944 218796 40996
rect 218848 40984 218854 40996
rect 253382 40984 253388 40996
rect 218848 40956 253388 40984
rect 218848 40944 218854 40956
rect 253382 40944 253388 40956
rect 253440 40944 253446 40996
rect 374822 40944 374828 40996
rect 374880 40984 374886 40996
rect 398190 40984 398196 40996
rect 374880 40956 398196 40984
rect 374880 40944 374886 40956
rect 398190 40944 398196 40956
rect 398248 40944 398254 40996
rect 53374 40876 53380 40928
rect 53432 40916 53438 40928
rect 86494 40916 86500 40928
rect 53432 40888 86500 40916
rect 53432 40876 53438 40888
rect 86494 40876 86500 40888
rect 86552 40876 86558 40928
rect 219066 40876 219072 40928
rect 219124 40916 219130 40928
rect 251174 40916 251180 40928
rect 219124 40888 251180 40916
rect 219124 40876 219130 40888
rect 251174 40876 251180 40888
rect 251232 40876 251238 40928
rect 59078 40808 59084 40860
rect 59136 40848 59142 40860
rect 92382 40848 92388 40860
rect 59136 40820 92388 40848
rect 59136 40808 59142 40820
rect 92382 40808 92388 40820
rect 92440 40808 92446 40860
rect 216030 40808 216036 40860
rect 216088 40848 216094 40860
rect 246390 40848 246396 40860
rect 216088 40820 246396 40848
rect 216088 40808 216094 40820
rect 246390 40808 246396 40820
rect 246448 40808 246454 40860
rect 55858 40740 55864 40792
rect 55916 40780 55922 40792
rect 87598 40780 87604 40792
rect 55916 40752 87604 40780
rect 55916 40740 55922 40752
rect 87598 40740 87604 40752
rect 87656 40740 87662 40792
rect 214650 40740 214656 40792
rect 214708 40780 214714 40792
rect 245286 40780 245292 40792
rect 214708 40752 245292 40780
rect 214708 40740 214714 40752
rect 245286 40740 245292 40752
rect 245344 40740 245350 40792
rect 51626 40672 51632 40724
rect 51684 40712 51690 40724
rect 78214 40712 78220 40724
rect 51684 40684 78220 40712
rect 51684 40672 51690 40684
rect 78214 40672 78220 40684
rect 78272 40672 78278 40724
rect 213362 40672 213368 40724
rect 213420 40712 213426 40724
rect 239122 40712 239128 40724
rect 213420 40684 239128 40712
rect 213420 40672 213426 40684
rect 239122 40672 239128 40684
rect 239180 40672 239186 40724
rect 53466 40604 53472 40656
rect 53524 40644 53530 40656
rect 80422 40644 80428 40656
rect 53524 40616 80428 40644
rect 53524 40604 53530 40616
rect 80422 40604 80428 40616
rect 80480 40604 80486 40656
rect 215018 40604 215024 40656
rect 215076 40644 215082 40656
rect 241606 40644 241612 40656
rect 215076 40616 241612 40644
rect 215076 40604 215082 40616
rect 241606 40604 241612 40616
rect 241664 40604 241670 40656
rect 54754 39992 54760 40044
rect 54812 40032 54818 40044
rect 116302 40032 116308 40044
rect 54812 40004 116308 40032
rect 54812 39992 54818 40004
rect 116302 39992 116308 40004
rect 116360 39992 116366 40044
rect 213638 39992 213644 40044
rect 213696 40032 213702 40044
rect 240502 40032 240508 40044
rect 213696 40004 240508 40032
rect 213696 39992 213702 40004
rect 240502 39992 240508 40004
rect 240560 39992 240566 40044
rect 375190 39992 375196 40044
rect 375248 40032 375254 40044
rect 399386 40032 399392 40044
rect 375248 40004 399392 40032
rect 375248 39992 375254 40004
rect 399386 39992 399392 40004
rect 399444 39992 399450 40044
rect 51994 39924 52000 39976
rect 52052 39964 52058 39976
rect 111886 39964 111892 39976
rect 52052 39936 111892 39964
rect 52052 39924 52058 39936
rect 111886 39924 111892 39936
rect 111944 39924 111950 39976
rect 214834 39924 214840 39976
rect 214892 39964 214898 39976
rect 238110 39964 238116 39976
rect 214892 39936 238116 39964
rect 214892 39924 214898 39936
rect 238110 39924 238116 39936
rect 238168 39924 238174 39976
rect 376662 39924 376668 39976
rect 376720 39964 376726 39976
rect 436370 39964 436376 39976
rect 376720 39936 436376 39964
rect 376720 39924 376726 39936
rect 436370 39924 436376 39936
rect 436428 39924 436434 39976
rect 52178 39856 52184 39908
rect 52236 39896 52242 39908
rect 111150 39896 111156 39908
rect 52236 39868 111156 39896
rect 52236 39856 52242 39868
rect 111150 39856 111156 39868
rect 111208 39856 111214 39908
rect 216398 39856 216404 39908
rect 216456 39896 216462 39908
rect 272150 39896 272156 39908
rect 216456 39868 272156 39896
rect 216456 39856 216462 39868
rect 272150 39856 272156 39868
rect 272208 39856 272214 39908
rect 374454 39856 374460 39908
rect 374512 39896 374518 39908
rect 434622 39896 434628 39908
rect 374512 39868 434628 39896
rect 374512 39856 374518 39868
rect 434622 39856 434628 39868
rect 434680 39856 434686 39908
rect 55030 39788 55036 39840
rect 55088 39828 55094 39840
rect 109310 39828 109316 39840
rect 55088 39800 109316 39828
rect 55088 39788 55094 39800
rect 109310 39788 109316 39800
rect 109368 39788 109374 39840
rect 215938 39788 215944 39840
rect 215996 39828 216002 39840
rect 269758 39828 269764 39840
rect 215996 39800 269764 39828
rect 215996 39788 216002 39800
rect 269758 39788 269764 39800
rect 269816 39788 269822 39840
rect 373810 39788 373816 39840
rect 373868 39828 373874 39840
rect 432138 39828 432144 39840
rect 373868 39800 432144 39828
rect 373868 39788 373874 39800
rect 432138 39788 432144 39800
rect 432196 39788 432202 39840
rect 44082 39720 44088 39772
rect 44140 39760 44146 39772
rect 90726 39760 90732 39772
rect 44140 39732 90732 39760
rect 44140 39720 44146 39732
rect 90726 39720 90732 39732
rect 90784 39720 90790 39772
rect 219802 39720 219808 39772
rect 219860 39760 219866 39772
rect 266630 39760 266636 39772
rect 219860 39732 266636 39760
rect 219860 39720 219866 39732
rect 266630 39720 266636 39732
rect 266688 39720 266694 39772
rect 375282 39720 375288 39772
rect 375340 39760 375346 39772
rect 431126 39760 431132 39772
rect 375340 39732 431132 39760
rect 375340 39720 375346 39732
rect 431126 39720 431132 39732
rect 431184 39720 431190 39772
rect 56962 39652 56968 39704
rect 57020 39692 57026 39704
rect 91278 39692 91284 39704
rect 57020 39664 91284 39692
rect 57020 39652 57026 39664
rect 91278 39652 91284 39664
rect 91336 39652 91342 39704
rect 219894 39652 219900 39704
rect 219952 39692 219958 39704
rect 266354 39692 266360 39704
rect 219952 39664 266360 39692
rect 219952 39652 219958 39664
rect 266354 39652 266360 39664
rect 266412 39652 266418 39704
rect 377582 39652 377588 39704
rect 377640 39692 377646 39704
rect 411898 39692 411904 39704
rect 377640 39664 411904 39692
rect 377640 39652 377646 39664
rect 411898 39652 411904 39664
rect 411956 39652 411962 39704
rect 59170 39584 59176 39636
rect 59228 39624 59234 39636
rect 93302 39624 93308 39636
rect 59228 39596 93308 39624
rect 59228 39584 59234 39596
rect 93302 39584 93308 39596
rect 93360 39584 93366 39636
rect 219710 39584 219716 39636
rect 219768 39624 219774 39636
rect 254118 39624 254124 39636
rect 219768 39596 254124 39624
rect 219768 39584 219774 39596
rect 254118 39584 254124 39596
rect 254176 39584 254182 39636
rect 379330 39584 379336 39636
rect 379388 39624 379394 39636
rect 411254 39624 411260 39636
rect 379388 39596 411260 39624
rect 379388 39584 379394 39596
rect 411254 39584 411260 39596
rect 411312 39584 411318 39636
rect 56410 39516 56416 39568
rect 56468 39556 56474 39568
rect 88610 39556 88616 39568
rect 56468 39528 88616 39556
rect 56468 39516 56474 39528
rect 88610 39516 88616 39528
rect 88668 39516 88674 39568
rect 217594 39516 217600 39568
rect 217652 39556 217658 39568
rect 251726 39556 251732 39568
rect 217652 39528 251732 39556
rect 217652 39516 217658 39528
rect 251726 39516 251732 39528
rect 251784 39516 251790 39568
rect 376570 39516 376576 39568
rect 376628 39556 376634 39568
rect 408678 39556 408684 39568
rect 376628 39528 408684 39556
rect 376628 39516 376634 39528
rect 408678 39516 408684 39528
rect 408736 39516 408742 39568
rect 59262 39448 59268 39500
rect 59320 39488 59326 39500
rect 89990 39488 89996 39500
rect 59320 39460 89996 39488
rect 59320 39448 59326 39460
rect 89990 39448 89996 39460
rect 90048 39448 90054 39500
rect 216306 39448 216312 39500
rect 216364 39488 216370 39500
rect 248598 39488 248604 39500
rect 216364 39460 248604 39488
rect 216364 39448 216370 39460
rect 248598 39448 248604 39460
rect 248656 39448 248662 39500
rect 372430 39448 372436 39500
rect 372488 39488 372494 39500
rect 400306 39488 400312 39500
rect 372488 39460 400312 39488
rect 372488 39448 372494 39460
rect 400306 39448 400312 39460
rect 400364 39448 400370 39500
rect 53650 39380 53656 39432
rect 53708 39420 53714 39432
rect 81802 39420 81808 39432
rect 53708 39392 81808 39420
rect 53708 39380 53714 39392
rect 81802 39380 81808 39392
rect 81860 39380 81866 39432
rect 219158 39380 219164 39432
rect 219216 39420 219222 39432
rect 247678 39420 247684 39432
rect 219216 39392 247684 39420
rect 219216 39380 219222 39392
rect 247678 39380 247684 39392
rect 247736 39380 247742 39432
rect 375006 39380 375012 39432
rect 375064 39420 375070 39432
rect 435174 39420 435180 39432
rect 375064 39392 435180 39420
rect 375064 39380 375070 39392
rect 435174 39380 435180 39392
rect 435232 39380 435238 39432
rect 51902 39312 51908 39364
rect 51960 39352 51966 39364
rect 78766 39352 78772 39364
rect 51960 39324 78772 39352
rect 51960 39312 51966 39324
rect 78766 39312 78772 39324
rect 78824 39312 78830 39364
rect 213546 39312 213552 39364
rect 213604 39352 213610 39364
rect 274726 39352 274732 39364
rect 213604 39324 274732 39352
rect 213604 39312 213610 39324
rect 274726 39312 274732 39324
rect 274784 39312 274790 39364
rect 212350 39244 212356 39296
rect 212408 39284 212414 39296
rect 273530 39284 273536 39296
rect 212408 39256 273536 39284
rect 212408 39244 212414 39256
rect 273530 39244 273536 39256
rect 273588 39244 273594 39296
rect 2774 31696 2780 31748
rect 2832 31736 2838 31748
rect 580442 31736 580448 31748
rect 2832 31708 580448 31736
rect 2832 31696 2838 31708
rect 580442 31696 580448 31708
rect 580500 31696 580506 31748
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2774 3516 2780 3528
rect 1728 3488 2780 3516
rect 1728 3476 1734 3488
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 57238 3448 57244 3460
rect 624 3420 57244 3448
rect 624 3408 630 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
<< via1 >>
rect 38384 700952 38436 701004
rect 99840 700952 99892 701004
rect 161296 700952 161348 701004
rect 222752 700952 222804 701004
rect 284208 700952 284260 701004
rect 345756 700952 345808 701004
rect 407212 700952 407264 701004
rect 468668 700952 468720 701004
rect 530124 700952 530176 701004
rect 531228 700952 531280 701004
rect 253480 700340 253532 700392
rect 305644 700340 305696 700392
rect 69112 700272 69164 700324
rect 304264 700272 304316 700324
rect 531228 700272 531280 700324
rect 580264 700272 580316 700324
rect 37924 699660 37976 699712
rect 38384 699660 38436 699712
rect 436744 699660 436796 699712
rect 437940 699660 437992 699712
rect 315028 698912 315080 698964
rect 400220 698912 400272 698964
rect 59268 697552 59320 697604
rect 545488 697552 545540 697604
rect 3424 684496 3476 684548
rect 316684 684496 316736 684548
rect 2780 660288 2832 660340
rect 37924 660288 37976 660340
rect 137560 658248 137612 658300
rect 579896 658248 579948 658300
rect 318800 651992 318852 652044
rect 498200 651992 498252 652044
rect 129740 650632 129792 650684
rect 429292 650632 429344 650684
rect 291200 650020 291252 650072
rect 457444 650020 457496 650072
rect 191840 649272 191892 649324
rect 430580 649272 430632 649324
rect 280988 648728 281040 648780
rect 430672 648728 430724 648780
rect 289820 648660 289872 648712
rect 489920 648660 489972 648712
rect 217784 648592 217836 648644
rect 580264 648592 580316 648644
rect 318248 648116 318300 648168
rect 427820 648116 427872 648168
rect 312544 648048 312596 648100
rect 332600 648048 332652 648100
rect 298744 647980 298796 648032
rect 378324 647980 378376 648032
rect 319720 647912 319772 647964
rect 355140 647912 355192 647964
rect 313924 647844 313976 647896
rect 359556 647844 359608 647896
rect 375380 647844 375432 647896
rect 423864 647844 423916 647896
rect 316868 647776 316920 647828
rect 364340 647776 364392 647828
rect 319812 647708 319864 647760
rect 373172 647708 373224 647760
rect 315304 647640 315356 647692
rect 368572 647640 368624 647692
rect 284944 647572 284996 647624
rect 350540 647572 350592 647624
rect 314016 647504 314068 647556
rect 382740 647504 382792 647556
rect 318156 647436 318208 647488
rect 387340 647436 387392 647488
rect 316776 647368 316828 647420
rect 396356 647368 396408 647420
rect 318064 647300 318116 647352
rect 337108 647300 337160 647352
rect 319628 647232 319680 647284
rect 323492 647232 323544 647284
rect 280712 646620 280764 646672
rect 341524 646620 341576 646672
rect 296720 646552 296772 646604
rect 429936 646552 429988 646604
rect 298100 646484 298152 646536
rect 432604 646484 432656 646536
rect 291292 646416 291344 646468
rect 428464 646416 428516 646468
rect 288532 646348 288584 646400
rect 429844 646348 429896 646400
rect 319444 646280 319496 646332
rect 466736 646280 466788 646332
rect 282184 646212 282236 646264
rect 430764 646212 430816 646264
rect 293960 646144 294012 646196
rect 497648 646144 497700 646196
rect 296812 646076 296864 646128
rect 512000 646076 512052 646128
rect 288440 646008 288492 646060
rect 510620 646008 510672 646060
rect 40684 645940 40736 645992
rect 409880 645940 409932 645992
rect 218704 645872 218756 645924
rect 414388 645872 414440 645924
rect 302884 644444 302936 644496
rect 317604 644444 317656 644496
rect 136548 640840 136600 640892
rect 149060 640840 149112 640892
rect 134892 640772 134944 640824
rect 140320 640772 140372 640824
rect 213920 640772 213972 640824
rect 225788 640772 225840 640824
rect 100576 640704 100628 640756
rect 124496 640704 124548 640756
rect 139860 640704 139912 640756
rect 157432 640704 157484 640756
rect 212540 640704 212592 640756
rect 272156 640704 272208 640756
rect 115388 640636 115440 640688
rect 124588 640636 124640 640688
rect 137836 640636 137888 640688
rect 160652 640636 160704 640688
rect 217876 640636 217928 640688
rect 243176 640636 243228 640688
rect 56508 640568 56560 640620
rect 77392 640568 77444 640620
rect 112168 640568 112220 640620
rect 124680 640568 124732 640620
rect 134984 640568 135036 640620
rect 140228 640568 140280 640620
rect 140320 640568 140372 640620
rect 166448 640568 166500 640620
rect 218888 640568 218940 640620
rect 252192 640568 252244 640620
rect 54944 640500 54996 640552
rect 80612 640500 80664 640552
rect 109592 640500 109644 640552
rect 122840 640500 122892 640552
rect 139216 640500 139268 640552
rect 174820 640500 174872 640552
rect 189632 640500 189684 640552
rect 205640 640500 205692 640552
rect 218796 640500 218848 640552
rect 263784 640500 263836 640552
rect 54852 640432 54904 640484
rect 88984 640432 89036 640484
rect 106372 640432 106424 640484
rect 121460 640432 121512 640484
rect 137652 640432 137704 640484
rect 140136 640432 140188 640484
rect 140228 640432 140280 640484
rect 180616 640432 180668 640484
rect 214012 640432 214064 640484
rect 269580 640432 269632 640484
rect 55128 640364 55180 640416
rect 92204 640364 92256 640416
rect 103796 640364 103848 640416
rect 120816 640364 120868 640416
rect 124220 640364 124272 640416
rect 172244 640364 172296 640416
rect 192208 640364 192260 640416
rect 204352 640364 204404 640416
rect 219348 640364 219400 640416
rect 275376 640364 275428 640416
rect 55036 640296 55088 640348
rect 94780 640296 94832 640348
rect 133880 640296 133932 640348
rect 140044 640296 140096 640348
rect 140136 640296 140188 640348
rect 186412 640296 186464 640348
rect 195428 640296 195480 640348
rect 200856 640296 200908 640348
rect 217324 640296 217376 640348
rect 231584 640296 231636 640348
rect 287704 640296 287756 640348
rect 317696 640296 317748 640348
rect 215300 639208 215352 639260
rect 234804 639208 234856 639260
rect 219624 639140 219676 639192
rect 246396 639140 246448 639192
rect 210424 639072 210476 639124
rect 237380 639072 237432 639124
rect 133144 639004 133196 639056
rect 151636 639004 151688 639056
rect 206284 639004 206336 639056
rect 254768 639004 254820 639056
rect 69020 638936 69072 638988
rect 124312 638936 124364 638988
rect 135260 638936 135312 638988
rect 183836 638936 183888 638988
rect 204260 638936 204312 638988
rect 277952 638936 278004 638988
rect 223764 638188 223816 638240
rect 215944 638120 215996 638172
rect 217968 638052 218020 638104
rect 228732 638052 228784 638104
rect 126244 637984 126296 638036
rect 177856 637984 177908 638036
rect 204904 637984 204956 638036
rect 223764 637984 223816 638036
rect 135168 637916 135220 637968
rect 145564 637916 145616 637968
rect 213184 637916 213236 637968
rect 222844 637916 222896 637968
rect 266268 637984 266320 638036
rect 260196 637916 260248 637968
rect 57796 637848 57848 637900
rect 71228 637848 71280 637900
rect 136456 637848 136508 637900
rect 154580 637848 154632 637900
rect 208400 637848 208452 637900
rect 240324 637848 240376 637900
rect 56324 637780 56376 637832
rect 65524 637780 65576 637832
rect 135076 637780 135128 637832
rect 162860 637780 162912 637832
rect 206376 637780 206428 637832
rect 248696 637780 248748 637832
rect 59360 637712 59412 637764
rect 97908 637712 97960 637764
rect 56416 637644 56468 637696
rect 62948 637644 63000 637696
rect 86776 637644 86828 637696
rect 124404 637712 124456 637764
rect 138664 637712 138716 637764
rect 168748 637712 168800 637764
rect 210516 637712 210568 637764
rect 257620 637712 257672 637764
rect 59176 637576 59228 637628
rect 74632 637576 74684 637628
rect 83464 637576 83516 637628
rect 121644 637644 121696 637696
rect 138756 637644 138808 637696
rect 142988 637644 143040 637696
rect 198280 637644 198332 637696
rect 201500 637644 201552 637696
rect 216036 637644 216088 637696
rect 219716 637644 219768 637696
rect 118240 637576 118292 637628
rect 120908 637576 120960 637628
rect 137928 637576 137980 637628
rect 218704 637576 218756 637628
rect 280712 637440 280764 637492
rect 280712 637236 280764 637288
rect 429936 636896 429988 636948
rect 474740 636896 474792 636948
rect 432604 636828 432656 636880
rect 505468 636828 505520 636880
rect 482928 636216 482980 636268
rect 511356 636216 511408 636268
rect 206468 634788 206520 634840
rect 216680 634788 216732 634840
rect 289084 634788 289136 634840
rect 317972 634788 318024 634840
rect 428464 634720 428516 634772
rect 456800 634720 456852 634772
rect 208492 632068 208544 632120
rect 216680 632068 216732 632120
rect 307024 630640 307076 630692
rect 317420 630640 317472 630692
rect 211804 626560 211856 626612
rect 216680 626560 216732 626612
rect 429844 626492 429896 626544
rect 456800 626492 456852 626544
rect 311164 625132 311216 625184
rect 317972 625132 318024 625184
rect 132500 622412 132552 622464
rect 136640 622412 136692 622464
rect 204996 622412 205048 622464
rect 216680 622412 216732 622464
rect 287796 620984 287848 621036
rect 317972 620984 318024 621036
rect 135352 618196 135404 618248
rect 137284 618196 137336 618248
rect 295984 615476 296036 615528
rect 317420 615476 317472 615528
rect 286324 611328 286376 611380
rect 317972 611328 318024 611380
rect 134524 604460 134576 604512
rect 137376 604460 137428 604512
rect 213276 604460 213328 604512
rect 216680 604460 216732 604512
rect 124128 603100 124180 603152
rect 134616 603100 134668 603152
rect 203892 603100 203944 603152
rect 216772 603100 216824 603152
rect 283656 603100 283708 603152
rect 300216 603100 300268 603152
rect 211160 601672 211212 601724
rect 216680 601672 216732 601724
rect 296076 601672 296128 601724
rect 317972 601672 318024 601724
rect 57428 600244 57480 600296
rect 58624 600244 58676 600296
rect 214564 597524 214616 597576
rect 217048 597524 217100 597576
rect 286416 597524 286468 597576
rect 317972 597524 318024 597576
rect 217692 595960 217744 596012
rect 218704 595960 218756 596012
rect 125600 592016 125652 592068
rect 136640 592016 136692 592068
rect 210608 592016 210660 592068
rect 216680 592016 216732 592068
rect 300124 592016 300176 592068
rect 317972 592016 318024 592068
rect 130384 589296 130436 589348
rect 136640 589296 136692 589348
rect 209044 589296 209096 589348
rect 216680 589296 216732 589348
rect 210700 586508 210752 586560
rect 216680 586508 216732 586560
rect 289176 586508 289228 586560
rect 317420 586508 317472 586560
rect 300216 584128 300268 584180
rect 302240 584128 302292 584180
rect 281632 583312 281684 583364
rect 282276 583312 282328 583364
rect 207020 577464 207072 577516
rect 217416 577464 217468 577516
rect 57888 576172 57940 576224
rect 137284 576172 137336 576224
rect 217692 576172 217744 576224
rect 219900 576172 219952 576224
rect 57244 575492 57296 575544
rect 60372 575492 60424 575544
rect 137376 575492 137428 575544
rect 140136 575492 140188 575544
rect 200948 575492 201000 575544
rect 203340 575492 203392 575544
rect 3516 575424 3568 575476
rect 286416 575424 286468 575476
rect 134616 575356 134668 575408
rect 216772 575356 216824 575408
rect 302240 575356 302292 575408
rect 58440 575220 58492 575272
rect 62396 575220 62448 575272
rect 139216 575220 139268 575272
rect 142160 575220 142212 575272
rect 139860 575152 139912 575204
rect 140780 575152 140832 575204
rect 164332 575152 164384 575204
rect 200856 575152 200908 575204
rect 106280 575084 106332 575136
rect 124588 575084 124640 575136
rect 137652 575084 137704 575136
rect 145472 575084 145524 575136
rect 183468 575084 183520 575136
rect 218888 575084 218940 575136
rect 100392 575016 100444 575068
rect 121552 575016 121604 575068
rect 156236 575016 156288 575068
rect 205640 575016 205692 575068
rect 98184 574948 98236 575000
rect 122840 574948 122892 575000
rect 138848 574948 138900 575000
rect 149152 574948 149204 575000
rect 154580 574948 154632 575000
rect 204352 574948 204404 575000
rect 219348 574948 219400 575000
rect 223580 574948 223632 575000
rect 273260 574948 273312 575000
rect 318248 574948 318300 575000
rect 54852 574880 54904 574932
rect 78680 574880 78732 574932
rect 97448 574880 97500 574932
rect 124680 574880 124732 574932
rect 129740 574880 129792 574932
rect 202972 574880 203024 574932
rect 217876 574880 217928 574932
rect 222200 574880 222252 574932
rect 229284 574880 229336 574932
rect 281264 574880 281316 574932
rect 57612 574812 57664 574864
rect 83188 574812 83240 574864
rect 93860 574812 93912 574864
rect 124496 574812 124548 574864
rect 134984 574812 135036 574864
rect 151912 574812 151964 574864
rect 197084 574812 197136 574864
rect 282000 574812 282052 574864
rect 63500 574744 63552 574796
rect 123576 574744 123628 574796
rect 134892 574744 134944 574796
rect 161940 574744 161992 574796
rect 179420 574744 179472 574796
rect 281632 574744 281684 574796
rect 58808 574268 58860 574320
rect 60924 574268 60976 574320
rect 139032 574200 139084 574252
rect 141240 574200 141292 574252
rect 302240 574064 302292 574116
rect 302976 574064 303028 574116
rect 59452 573860 59504 573912
rect 63224 573860 63276 573912
rect 112536 573656 112588 573708
rect 123024 573656 123076 573708
rect 88156 573588 88208 573640
rect 120908 573588 120960 573640
rect 129004 573588 129056 573640
rect 203156 573588 203208 573640
rect 57152 573520 57204 573572
rect 81716 573520 81768 573572
rect 86960 573520 87012 573572
rect 121460 573520 121512 573572
rect 126152 573520 126204 573572
rect 201960 573520 202012 573572
rect 219256 573520 219308 573572
rect 224316 573520 224368 573572
rect 240784 573520 240836 573572
rect 315304 573520 315356 573572
rect 59268 573452 59320 573504
rect 68836 573452 68888 573504
rect 78864 573452 78916 573504
rect 122288 573452 122340 573504
rect 186320 573452 186372 573504
rect 282920 573452 282972 573504
rect 67640 573384 67692 573436
rect 121828 573384 121880 573436
rect 139124 573384 139176 573436
rect 150624 573384 150676 573436
rect 182272 573384 182324 573436
rect 281540 573384 281592 573436
rect 64512 573316 64564 573368
rect 122932 573316 122984 573368
rect 137008 573316 137060 573368
rect 160560 573316 160612 573368
rect 180800 573316 180852 573368
rect 283380 573316 283432 573368
rect 268016 572704 268068 572756
rect 317972 572704 318024 572756
rect 150992 572500 151044 572552
rect 160744 572500 160796 572552
rect 198004 572500 198056 572552
rect 200580 572500 200632 572552
rect 267004 572500 267056 572552
rect 268936 572500 268988 572552
rect 148416 572432 148468 572484
rect 159364 572432 159416 572484
rect 143540 572364 143592 572416
rect 156788 572364 156840 572416
rect 160008 572364 160060 572416
rect 164884 572364 164936 572416
rect 82544 572296 82596 572348
rect 88984 572296 89036 572348
rect 147680 572296 147732 572348
rect 162584 572296 162636 572348
rect 74540 572228 74592 572280
rect 97356 572228 97408 572280
rect 99932 572228 99984 572280
rect 115480 572228 115532 572280
rect 154856 572228 154908 572280
rect 171600 572228 171652 572280
rect 232228 572228 232280 572280
rect 259920 572228 259972 572280
rect 62580 572160 62632 572212
rect 71044 572160 71096 572212
rect 85764 572160 85816 572212
rect 108304 572160 108356 572212
rect 129832 572160 129884 572212
rect 154212 572160 154264 572212
rect 158720 572160 158772 572212
rect 183192 572160 183244 572212
rect 188344 572160 188396 572212
rect 203432 572160 203484 572212
rect 222292 572160 222344 572212
rect 254124 572160 254176 572212
rect 269672 572160 269724 572212
rect 286324 572160 286376 572212
rect 68376 572092 68428 572144
rect 105544 572092 105596 572144
rect 119712 572092 119764 572144
rect 145196 572092 145248 572144
rect 147772 572092 147824 572144
rect 185768 572092 185820 572144
rect 190460 572092 190512 572144
rect 257344 572092 257396 572144
rect 263692 572092 263744 572144
rect 312544 572092 312596 572144
rect 70952 572024 71004 572076
rect 108396 572024 108448 572076
rect 110420 572024 110472 572076
rect 120724 572024 120776 572076
rect 134156 572024 134208 572076
rect 197360 572024 197412 572076
rect 227904 572024 227956 572076
rect 245752 572024 245804 572076
rect 247040 572024 247092 572076
rect 319812 572024 319864 572076
rect 58900 571956 58952 572008
rect 74632 571956 74684 572008
rect 76840 571956 76892 572008
rect 117320 571956 117372 572008
rect 132684 571956 132736 572008
rect 177396 571956 177448 572008
rect 192760 571956 192812 572008
rect 277308 571956 277360 572008
rect 113272 571616 113324 571668
rect 121092 571616 121144 571668
rect 94136 571412 94188 571464
rect 101404 571412 101456 571464
rect 262864 571412 262916 571464
rect 265716 571412 265768 571464
rect 60004 571344 60056 571396
rect 61384 571344 61436 571396
rect 72424 571344 72476 571396
rect 74172 571344 74224 571396
rect 76748 571344 76800 571396
rect 83464 571344 83516 571396
rect 91560 571344 91612 571396
rect 93124 571344 93176 571396
rect 100760 571344 100812 571396
rect 103152 571344 103204 571396
rect 106924 571344 106976 571396
rect 108948 571344 109000 571396
rect 116584 571344 116636 571396
rect 120540 571344 120592 571396
rect 165804 571344 165856 571396
rect 167828 571344 167880 571396
rect 171784 571344 171836 571396
rect 174176 571344 174228 571396
rect 184204 571344 184256 571396
rect 188988 571344 189040 571396
rect 219992 571344 220044 571396
rect 221464 571344 221516 571396
rect 222568 571344 222620 571396
rect 224960 571344 225012 571396
rect 225052 571344 225104 571396
rect 228364 571344 228416 571396
rect 260104 571344 260156 571396
rect 263140 571344 263192 571396
rect 269764 571344 269816 571396
rect 271512 571344 271564 571396
rect 278044 571344 278096 571396
rect 280528 571344 280580 571396
rect 193220 570868 193272 570920
rect 218796 570868 218848 570920
rect 94596 570800 94648 570852
rect 123300 570800 123352 570852
rect 168472 570800 168524 570852
rect 200672 570800 200724 570852
rect 57336 570732 57388 570784
rect 89812 570732 89864 570784
rect 122840 570732 122892 570784
rect 202144 570732 202196 570784
rect 215852 570732 215904 570784
rect 281172 570732 281224 570784
rect 65984 570664 66036 570716
rect 121920 570664 121972 570716
rect 137928 570664 137980 570716
rect 169116 570664 169168 570716
rect 180616 570664 180668 570716
rect 282276 570664 282328 570716
rect 7564 570596 7616 570648
rect 317512 570596 317564 570648
rect 266636 569440 266688 569492
rect 298744 569440 298796 569492
rect 59084 569372 59136 569424
rect 92572 569372 92624 569424
rect 138296 569372 138348 569424
rect 200764 569372 200816 569424
rect 250076 569372 250128 569424
rect 295984 569372 296036 569424
rect 79968 569304 80020 569356
rect 114744 569304 114796 569356
rect 195244 569304 195296 569356
rect 283012 569304 283064 569356
rect 69020 569236 69072 569288
rect 123484 569236 123536 569288
rect 138480 569236 138532 569288
rect 159088 569236 159140 569288
rect 181352 569236 181404 569288
rect 281908 569236 281960 569288
rect 3424 569168 3476 569220
rect 319812 569168 319864 569220
rect 193496 568012 193548 568064
rect 206468 568012 206520 568064
rect 259460 568012 259512 568064
rect 302884 568012 302936 568064
rect 170588 567944 170640 567996
rect 201776 567944 201828 567996
rect 255320 567944 255372 567996
rect 309784 567944 309836 567996
rect 57060 567876 57112 567928
rect 101496 567876 101548 567928
rect 187056 567876 187108 567928
rect 283288 567876 283340 567928
rect 70952 567808 71004 567860
rect 123208 567808 123260 567860
rect 137100 567808 137152 567860
rect 166264 567808 166316 567860
rect 183560 567808 183612 567860
rect 281724 567808 281776 567860
rect 11704 567196 11756 567248
rect 317972 567196 318024 567248
rect 266544 566720 266596 566772
rect 284944 566720 284996 566772
rect 84568 566652 84620 566704
rect 122104 566652 122156 566704
rect 157984 566652 158036 566704
rect 203064 566652 203116 566704
rect 226432 566652 226484 566704
rect 280804 566652 280856 566704
rect 188068 566584 188120 566636
rect 233240 566584 233292 566636
rect 257988 566584 258040 566636
rect 314016 566584 314068 566636
rect 58992 566516 59044 566568
rect 108212 566516 108264 566568
rect 122564 566516 122616 566568
rect 201592 566516 201644 566568
rect 213920 566516 213972 566568
rect 215024 566516 215076 566568
rect 245108 566516 245160 566568
rect 313924 566516 313976 566568
rect 65248 566448 65300 566500
rect 123392 566448 123444 566500
rect 138572 566448 138624 566500
rect 160652 566448 160704 566500
rect 194968 566448 195020 566500
rect 283564 566448 283616 566500
rect 220728 565360 220780 565412
rect 247132 565360 247184 565412
rect 190644 565292 190696 565344
rect 204996 565292 205048 565344
rect 228640 565292 228692 565344
rect 282092 565292 282144 565344
rect 88340 565224 88392 565276
rect 104624 565224 104676 565276
rect 177028 565224 177080 565276
rect 213276 565224 213328 565276
rect 246488 565224 246540 565276
rect 311164 565224 311216 565276
rect 71044 565156 71096 565208
rect 109684 565156 109736 565208
rect 142620 565156 142672 565208
rect 202052 565156 202104 565208
rect 206376 565156 206428 565208
rect 241520 565156 241572 565208
rect 242900 565156 242952 565208
rect 318156 565156 318208 565208
rect 57704 565088 57756 565140
rect 76840 565088 76892 565140
rect 80336 565088 80388 565140
rect 122012 565088 122064 565140
rect 122104 565088 122156 565140
rect 190552 565088 190604 565140
rect 196348 565088 196400 565140
rect 283104 565088 283156 565140
rect 135260 564884 135312 564936
rect 136180 564884 136232 564936
rect 304264 564340 304316 564392
rect 317972 564340 318024 564392
rect 197820 564000 197872 564052
rect 210700 564000 210752 564052
rect 177764 563932 177816 563984
rect 225144 563932 225196 563984
rect 89628 563864 89680 563916
rect 104900 563864 104952 563916
rect 144092 563864 144144 563916
rect 201684 563864 201736 563916
rect 260196 563864 260248 563916
rect 289176 563864 289228 563916
rect 80980 563796 81032 563848
rect 121000 563796 121052 563848
rect 189172 563796 189224 563848
rect 267004 563796 267056 563848
rect 59544 563728 59596 563780
rect 101036 563728 101088 563780
rect 142252 563728 142304 563780
rect 167736 563728 167788 563780
rect 200672 563728 200724 563780
rect 281816 563728 281868 563780
rect 66720 563660 66772 563712
rect 121184 563660 121236 563712
rect 121552 563660 121604 563712
rect 201132 563660 201184 563712
rect 234344 563660 234396 563712
rect 319720 563660 319772 563712
rect 158720 563388 158772 563440
rect 159824 563388 159876 563440
rect 189908 562572 189960 562624
rect 217324 562572 217376 562624
rect 205732 562504 205784 562556
rect 262864 562504 262916 562556
rect 86040 562436 86092 562488
rect 122196 562436 122248 562488
rect 138480 562436 138532 562488
rect 203248 562436 203300 562488
rect 212172 562436 212224 562488
rect 280896 562436 280948 562488
rect 58532 562368 58584 562420
rect 63132 562300 63184 562352
rect 69020 562232 69072 562284
rect 70308 562232 70360 562284
rect 74540 562232 74592 562284
rect 75276 562232 75328 562284
rect 78680 562232 78732 562284
rect 79600 562232 79652 562284
rect 89812 562300 89864 562352
rect 91008 562300 91060 562352
rect 100760 562368 100812 562420
rect 101772 562368 101824 562420
rect 127624 562368 127676 562420
rect 194600 562368 194652 562420
rect 199200 562368 199252 562420
rect 211804 562368 211856 562420
rect 218152 562368 218204 562420
rect 219256 562368 219308 562420
rect 222200 562368 222252 562420
rect 222844 562368 222896 562420
rect 224960 562368 225012 562420
rect 225788 562368 225840 562420
rect 255320 562368 255372 562420
rect 256516 562368 256568 562420
rect 102508 562300 102560 562352
rect 106280 562300 106332 562352
rect 107568 562300 107620 562352
rect 124220 562300 124272 562352
rect 125416 562300 125468 562352
rect 125600 562300 125652 562352
rect 126888 562300 126940 562352
rect 140780 562300 140832 562352
rect 141884 562300 141936 562352
rect 137468 562232 137520 562284
rect 173164 562300 173216 562352
rect 180800 562300 180852 562352
rect 181996 562300 182048 562352
rect 185584 562300 185636 562352
rect 143540 562232 143592 562284
rect 144736 562232 144788 562284
rect 147680 562232 147732 562284
rect 148324 562232 148376 562284
rect 154580 562232 154632 562284
rect 155500 562232 155552 562284
rect 164332 562232 164384 562284
rect 165528 562232 165580 562284
rect 208400 562232 208452 562284
rect 209228 562232 209280 562284
rect 110512 562164 110564 562216
rect 142160 562164 142212 562216
rect 143356 562164 143408 562216
rect 250812 562232 250864 562284
rect 319628 562368 319680 562420
rect 273260 562300 273312 562352
rect 274456 562300 274508 562352
rect 275192 562300 275244 562352
rect 318064 562300 318116 562352
rect 274640 562232 274692 562284
rect 283748 561824 283800 561876
rect 287796 561824 287848 561876
rect 192116 561212 192168 561264
rect 216036 561212 216088 561264
rect 178500 561144 178552 561196
rect 209044 561144 209096 561196
rect 217876 561144 217928 561196
rect 260104 561144 260156 561196
rect 61384 561076 61436 561128
rect 105360 561076 105412 561128
rect 140504 561076 140556 561128
rect 198004 561076 198056 561128
rect 209136 561076 209188 561128
rect 236000 561076 236052 561128
rect 251548 561076 251600 561128
rect 316868 561076 316920 561128
rect 69572 561008 69624 561060
rect 114652 561008 114704 561060
rect 139492 561008 139544 561060
rect 163412 561008 163464 561060
rect 198556 561008 198608 561060
rect 278044 561008 278096 561060
rect 279516 561008 279568 561060
rect 289084 561008 289136 561060
rect 71688 560940 71740 560992
rect 121736 560940 121788 560992
rect 124036 560940 124088 560992
rect 201868 560940 201920 560992
rect 207112 560940 207164 560992
rect 214564 560940 214616 560992
rect 235080 560940 235132 560992
rect 319536 560940 319588 560992
rect 190460 560804 190512 560856
rect 191380 560804 191432 560856
rect 237932 559852 237984 559904
rect 315488 559852 315540 559904
rect 269488 559784 269540 559836
rect 300124 559784 300176 559836
rect 57520 559716 57572 559768
rect 88248 559716 88300 559768
rect 184940 559716 184992 559768
rect 210608 559716 210660 559768
rect 253664 559716 253716 559768
rect 316776 559716 316828 559768
rect 73160 559648 73212 559700
rect 106924 559648 106976 559700
rect 136916 559648 136968 559700
rect 202236 559648 202288 559700
rect 210700 559648 210752 559700
rect 283196 559648 283248 559700
rect 82452 559580 82504 559632
rect 116584 559580 116636 559632
rect 124680 559580 124732 559632
rect 201224 559580 201276 559632
rect 202144 559580 202196 559632
rect 283472 559580 283524 559632
rect 58716 559512 58768 559564
rect 111064 559512 111116 559564
rect 120448 559512 120500 559564
rect 130384 559512 130436 559564
rect 179144 559512 179196 559564
rect 269764 559512 269816 559564
rect 282368 559512 282420 559564
rect 296076 559512 296128 559564
rect 293776 559444 293828 559496
rect 312728 559444 312780 559496
rect 286692 559376 286744 559428
rect 309784 559376 309836 559428
rect 288072 559308 288124 559360
rect 312544 559308 312596 559360
rect 285220 559240 285272 559292
rect 312820 559240 312872 559292
rect 284944 559172 284996 559224
rect 315304 559172 315356 559224
rect 284484 559104 284536 559156
rect 315580 559104 315632 559156
rect 284208 559036 284260 559088
rect 315396 559036 315448 559088
rect 193220 558968 193272 559020
rect 194232 558968 194284 559020
rect 242256 558968 242308 559020
rect 318248 558968 318300 559020
rect 293132 558900 293184 558952
rect 312912 558900 312964 558952
rect 138940 558288 138992 558340
rect 149796 558288 149848 558340
rect 152648 558288 152700 558340
rect 202880 558288 202932 558340
rect 244372 558288 244424 558340
rect 318064 558288 318116 558340
rect 131212 558220 131264 558272
rect 184204 558220 184256 558272
rect 219164 558220 219216 558272
rect 227168 558220 227220 558272
rect 271604 558220 271656 558272
rect 287704 558220 287756 558272
rect 57428 558152 57480 558204
rect 99196 558152 99248 558204
rect 99288 558152 99340 558204
rect 123116 558152 123168 558204
rect 128268 558152 128320 558204
rect 201040 558152 201092 558204
rect 212816 557948 212868 558000
rect 251180 558152 251232 558204
rect 265900 558152 265952 558204
rect 301504 558152 301556 558204
rect 273076 558084 273128 558136
rect 311164 558084 311216 558136
rect 264428 558016 264480 558068
rect 304356 558016 304408 558068
rect 260840 557948 260892 558000
rect 304264 557948 304316 558000
rect 273720 557880 273772 557932
rect 318156 557880 318208 557932
rect 272340 557812 272392 557864
rect 316684 557812 316736 557864
rect 254400 557744 254452 557796
rect 319628 557744 319680 557796
rect 252284 557676 252336 557728
rect 317972 557676 318024 557728
rect 247224 557608 247276 557660
rect 319536 557608 319588 557660
rect 287336 557540 287388 557592
rect 312636 557540 312688 557592
rect 61660 557472 61712 557524
rect 64880 557472 64932 557524
rect 83464 557472 83516 557524
rect 86776 557472 86828 557524
rect 131856 557472 131908 557524
rect 133144 557472 133196 557524
rect 187792 557472 187844 557524
rect 195244 557472 195296 557524
rect 511356 557472 511408 557524
rect 580172 557472 580224 557524
rect 55128 557404 55180 557456
rect 67364 557404 67416 557456
rect 68376 557404 68428 557456
rect 77392 557404 77444 557456
rect 101404 557404 101456 557456
rect 106096 557404 106148 557456
rect 108396 557404 108448 557456
rect 114652 557404 114704 557456
rect 277308 557404 277360 557456
rect 301688 557404 301740 557456
rect 56508 557336 56560 557388
rect 83924 557336 83976 557388
rect 138756 557336 138808 557388
rect 146944 557336 146996 557388
rect 164884 557336 164936 557388
rect 173440 557336 173492 557388
rect 278044 557336 278096 557388
rect 318616 557336 318668 557388
rect 55036 557268 55088 557320
rect 85304 557268 85356 557320
rect 137836 557268 137888 557320
rect 151268 557268 151320 557320
rect 159364 557268 159416 557320
rect 167000 557268 167052 557320
rect 257252 557268 257304 557320
rect 303068 557268 303120 557320
rect 56416 557200 56468 557252
rect 88892 557200 88944 557252
rect 60372 557132 60424 557184
rect 95332 557200 95384 557252
rect 139860 557200 139912 557252
rect 153384 557200 153436 557252
rect 164148 557200 164200 557252
rect 171784 557200 171836 557252
rect 252928 557200 252980 557252
rect 319352 557200 319404 557252
rect 114008 557132 114060 557184
rect 124312 557132 124364 557184
rect 135168 557132 135220 557184
rect 156972 557132 157024 557184
rect 160744 557132 160796 557184
rect 172704 557132 172756 557184
rect 255872 557132 255924 557184
rect 301780 557132 301832 557184
rect 54944 557064 54996 557116
rect 93032 557064 93084 557116
rect 93124 557064 93176 557116
rect 96804 557064 96856 557116
rect 99196 557064 99248 557116
rect 116860 557064 116912 557116
rect 118240 557064 118292 557116
rect 126244 557064 126296 557116
rect 135076 557064 135128 557116
rect 164884 557064 164936 557116
rect 58624 556996 58676 557048
rect 68376 556996 68428 557048
rect 68468 556996 68520 557048
rect 99656 556996 99708 557048
rect 106832 556996 106884 557048
rect 121644 556996 121696 557048
rect 136548 556996 136600 557048
rect 171968 557064 172020 557116
rect 176292 557064 176344 557116
rect 210516 557064 210568 557116
rect 261576 557064 261628 557116
rect 282184 557064 282236 557116
rect 171324 556996 171376 557048
rect 188344 556996 188396 557048
rect 199936 556996 199988 557048
rect 210424 556996 210476 557048
rect 217968 556996 218020 557048
rect 218612 556996 218664 557048
rect 245844 556996 245896 557048
rect 281080 556996 281132 557048
rect 63224 556928 63276 556980
rect 76012 556928 76064 556980
rect 76840 556928 76892 556980
rect 117596 556928 117648 556980
rect 118976 556928 119028 556980
rect 134524 556928 134576 556980
rect 137744 556928 137796 556980
rect 175556 556928 175608 556980
rect 195612 556928 195664 556980
rect 206468 556928 206520 556980
rect 218060 556928 218112 556980
rect 230020 556928 230072 556980
rect 231492 556928 231544 556980
rect 238760 556928 238812 556980
rect 239404 556928 239456 556980
rect 280988 556928 281040 556980
rect 56324 556860 56376 556912
rect 98920 556860 98972 556912
rect 103980 556860 104032 556912
rect 124404 556860 124456 556912
rect 136456 556860 136508 556912
rect 157708 556860 157760 556912
rect 158352 556860 158404 556912
rect 200948 556860 201000 556912
rect 220084 556860 220136 556912
rect 232872 556860 232924 556912
rect 238668 556860 238720 556912
rect 284944 556860 284996 556912
rect 57796 556792 57848 556844
rect 73804 556792 73856 556844
rect 78128 556792 78180 556844
rect 120816 556792 120868 556844
rect 146208 556792 146260 556844
rect 201500 556792 201552 556844
rect 204996 556792 205048 556844
rect 213184 556792 213236 556844
rect 218704 556792 218756 556844
rect 233608 556792 233660 556844
rect 237196 556792 237248 556844
rect 284208 556792 284260 556844
rect 299572 556792 299624 556844
rect 319444 556792 319496 556844
rect 59176 556724 59228 556776
rect 68468 556724 68520 556776
rect 105544 556724 105596 556776
rect 108948 556724 109000 556776
rect 275928 556724 275980 556776
rect 300400 556724 300452 556776
rect 270868 556656 270920 556708
rect 300216 556656 300268 556708
rect 285956 556588 286008 556640
rect 319720 556588 319772 556640
rect 280160 556520 280212 556572
rect 316868 556520 316920 556572
rect 88984 556452 89036 556504
rect 90364 556452 90416 556504
rect 262312 556452 262364 556504
rect 300308 556452 300360 556504
rect 173164 556384 173216 556436
rect 174912 556384 174964 556436
rect 240048 556384 240100 556436
rect 266360 556384 266412 556436
rect 281632 556384 281684 556436
rect 300124 556384 300176 556436
rect 101496 556316 101548 556368
rect 103244 556316 103296 556368
rect 108304 556316 108356 556368
rect 111800 556316 111852 556368
rect 202788 556316 202840 556368
rect 209136 556316 209188 556368
rect 283104 556316 283156 556368
rect 301596 556316 301648 556368
rect 88248 556248 88300 556300
rect 91744 556248 91796 556300
rect 137652 556248 137704 556300
rect 138664 556248 138716 556300
rect 162676 556248 162728 556300
rect 168380 556248 168432 556300
rect 174176 556248 174228 556300
rect 179512 556248 179564 556300
rect 201408 556248 201460 556300
rect 206284 556248 206336 556300
rect 209964 556248 210016 556300
rect 215944 556248 215996 556300
rect 293960 556248 294012 556300
rect 295248 556248 295300 556300
rect 296720 556248 296772 556300
rect 297364 556248 297416 556300
rect 298100 556248 298152 556300
rect 316776 556248 316828 556300
rect 96068 556180 96120 556232
rect 99288 556180 99340 556232
rect 115480 556180 115532 556232
rect 116124 556180 116176 556232
rect 121092 556180 121144 556232
rect 122104 556180 122156 556232
rect 154120 556180 154172 556232
rect 157984 556180 158036 556232
rect 167828 556180 167880 556232
rect 169852 556180 169904 556232
rect 203524 556180 203576 556232
rect 204904 556180 204956 556232
rect 276572 556180 276624 556232
rect 301872 556180 301924 556232
rect 295984 555704 296036 555756
rect 313096 555704 313148 555756
rect 294512 555636 294564 555688
rect 315672 555636 315724 555688
rect 278780 555568 278832 555620
rect 300768 555568 300820 555620
rect 268752 555500 268804 555552
rect 302884 555500 302936 555552
rect 266360 555432 266412 555484
rect 318708 555432 318760 555484
rect 263048 555364 263100 555416
rect 301964 555364 302016 555416
rect 265164 555296 265216 555348
rect 313004 555296 313056 555348
rect 243636 555228 243688 555280
rect 305736 555228 305788 555280
rect 236476 555160 236528 555212
rect 301412 555160 301464 555212
rect 249448 555092 249500 555144
rect 318432 555092 318484 555144
rect 235908 555024 235960 555076
rect 319444 555024 319496 555076
rect 300768 554684 300820 554736
rect 317972 554684 318024 554736
rect 301412 550536 301464 550588
rect 317420 550536 317472 550588
rect 305736 545028 305788 545080
rect 317972 545028 318024 545080
rect 430948 543192 431000 543244
rect 431408 543192 431460 543244
rect 430764 543056 430816 543108
rect 430948 543056 431000 543108
rect 319260 542988 319312 543040
rect 319444 542988 319496 543040
rect 319168 536256 319220 536308
rect 319536 536256 319588 536308
rect 312912 535372 312964 535424
rect 512184 535372 512236 535424
rect 313096 535304 313148 535356
rect 505100 535304 505152 535356
rect 312820 535236 312872 535288
rect 466460 535236 466512 535288
rect 300492 535168 300544 535220
rect 430672 535168 430724 535220
rect 300676 535100 300728 535152
rect 430764 535100 430816 535152
rect 303068 535032 303120 535084
rect 431316 535032 431368 535084
rect 315580 534964 315632 535016
rect 429476 534964 429528 535016
rect 316868 534896 316920 534948
rect 430580 534896 430632 534948
rect 318616 534828 318668 534880
rect 431224 534828 431276 534880
rect 319352 534760 319404 534812
rect 431132 534760 431184 534812
rect 318248 534692 318300 534744
rect 428464 534692 428516 534744
rect 300400 534148 300452 534200
rect 351276 534148 351328 534200
rect 305644 534080 305696 534132
rect 369308 534080 369360 534132
rect 309784 534012 309836 534064
rect 512092 534012 512144 534064
rect 318340 533944 318392 533996
rect 489920 533944 489972 533996
rect 319536 533876 319588 533928
rect 483020 533876 483072 533928
rect 302976 533808 303028 533860
rect 457628 533808 457680 533860
rect 312728 533740 312780 533792
rect 459560 533740 459612 533792
rect 315672 533672 315724 533724
rect 457536 533672 457588 533724
rect 316776 533604 316828 533656
rect 457444 533604 457496 533656
rect 300124 533536 300176 533588
rect 431040 533536 431092 533588
rect 300216 533468 300268 533520
rect 430856 533468 430908 533520
rect 301688 533400 301740 533452
rect 431408 533400 431460 533452
rect 301596 533332 301648 533384
rect 430948 533332 431000 533384
rect 301872 533264 301924 533316
rect 414940 533264 414992 533316
rect 301780 533196 301832 533248
rect 405924 533196 405976 533248
rect 300308 533128 300360 533180
rect 328644 533128 328696 533180
rect 304264 532652 304316 532704
rect 342260 532652 342312 532704
rect 313004 532584 313056 532636
rect 319628 532584 319680 532636
rect 319444 532516 319496 532568
rect 346676 532584 346728 532636
rect 319260 532448 319312 532500
rect 333244 532516 333296 532568
rect 319904 532448 319956 532500
rect 410524 532448 410576 532500
rect 302884 532380 302936 532432
rect 387892 532380 387944 532432
rect 301504 532312 301556 532364
rect 383660 532312 383712 532364
rect 318156 532244 318208 532296
rect 396908 532244 396960 532296
rect 304356 532176 304408 532228
rect 374460 532176 374512 532228
rect 311164 532108 311216 532160
rect 364708 532108 364760 532160
rect 319168 532040 319220 532092
rect 360292 532040 360344 532092
rect 318524 531972 318576 532024
rect 356244 531972 356296 532024
rect 316684 531904 316736 531956
rect 319904 531904 319956 531956
rect 319996 531904 320048 531956
rect 419540 531904 419592 531956
rect 318432 531836 318484 531888
rect 423956 531836 424008 531888
rect 301964 531768 302016 531820
rect 401600 531768 401652 531820
rect 318064 531700 318116 531752
rect 319996 531700 320048 531752
rect 312636 531224 312688 531276
rect 474740 531224 474792 531276
rect 315488 531156 315540 531208
rect 428372 531156 428424 531208
rect 303252 530544 303304 530596
rect 518164 530544 518216 530596
rect 312544 529864 312596 529916
rect 512000 529864 512052 529916
rect 315304 529796 315356 529848
rect 429384 529796 429436 529848
rect 315396 529728 315448 529780
rect 428556 529728 428608 529780
rect 302332 529184 302384 529236
rect 578884 529184 578936 529236
rect 42708 525036 42760 525088
rect 57704 525036 57756 525088
rect 302884 502324 302936 502376
rect 540244 502324 540296 502376
rect 82912 494912 82964 494964
rect 83188 494912 83240 494964
rect 128360 494912 128412 494964
rect 128544 494912 128596 494964
rect 136640 494912 136692 494964
rect 136916 494912 136968 494964
rect 176752 494912 176804 494964
rect 177028 494912 177080 494964
rect 229100 494912 229152 494964
rect 229468 494912 229520 494964
rect 259552 494912 259604 494964
rect 259828 494912 259880 494964
rect 197560 494776 197612 494828
rect 198280 494776 198332 494828
rect 207220 494776 207272 494828
rect 207388 494776 207440 494828
rect 242916 494776 242968 494828
rect 243084 494776 243136 494828
rect 244372 494776 244424 494828
rect 244556 494776 244608 494828
rect 273276 494776 273328 494828
rect 273444 494776 273496 494828
rect 284316 494776 284368 494828
rect 284484 494776 284536 494828
rect 498200 493960 498252 494012
rect 580172 493960 580224 494012
rect 56324 493348 56376 493400
rect 90548 493348 90600 493400
rect 51816 493280 51868 493332
rect 99380 493280 99432 493332
rect 109776 493280 109828 493332
rect 207112 493280 207164 493332
rect 161572 492736 161624 492788
rect 161940 492736 161992 492788
rect 167000 492736 167052 492788
rect 167736 492736 167788 492788
rect 219532 492736 219584 492788
rect 221004 492736 221056 492788
rect 221188 492736 221240 492788
rect 69112 492668 69164 492720
rect 69940 492668 69992 492720
rect 74632 492668 74684 492720
rect 75276 492668 75328 492720
rect 75920 492668 75972 492720
rect 76564 492668 76616 492720
rect 78680 492668 78732 492720
rect 79692 492668 79744 492720
rect 161480 492668 161532 492720
rect 161756 492668 161808 492720
rect 162860 492668 162912 492720
rect 163320 492668 163372 492720
rect 164240 492668 164292 492720
rect 165068 492668 165120 492720
rect 167092 492668 167144 492720
rect 167276 492668 167328 492720
rect 168472 492668 168524 492720
rect 169116 492668 169168 492720
rect 169852 492668 169904 492720
rect 170404 492668 170456 492720
rect 171232 492668 171284 492720
rect 172060 492668 172112 492720
rect 172612 492668 172664 492720
rect 173532 492668 173584 492720
rect 173992 492668 174044 492720
rect 174820 492668 174872 492720
rect 175280 492668 175332 492720
rect 176108 492668 176160 492720
rect 176660 492668 176712 492720
rect 177396 492668 177448 492720
rect 178040 492668 178092 492720
rect 178684 492668 178736 492720
rect 179420 492668 179472 492720
rect 180064 492668 180116 492720
rect 180892 492668 180944 492720
rect 181444 492668 181496 492720
rect 182180 492668 182232 492720
rect 182732 492668 182784 492720
rect 184940 492668 184992 492720
rect 185860 492668 185912 492720
rect 59268 492600 59320 492652
rect 60096 492532 60148 492584
rect 61936 492532 61988 492584
rect 62120 492532 62172 492584
rect 62948 492532 63000 492584
rect 63040 492532 63092 492584
rect 88800 492532 88852 492584
rect 139400 492600 139452 492652
rect 139860 492600 139912 492652
rect 150440 492600 150492 492652
rect 91100 492532 91152 492584
rect 92572 492532 92624 492584
rect 93308 492532 93360 492584
rect 129924 492532 129976 492584
rect 130108 492532 130160 492584
rect 50896 492464 50948 492516
rect 84384 492464 84436 492516
rect 92480 492464 92532 492516
rect 92940 492464 92992 492516
rect 102232 492464 102284 492516
rect 103060 492464 103112 492516
rect 106372 492464 106424 492516
rect 106924 492464 106976 492516
rect 107660 492464 107712 492516
rect 107844 492464 107896 492516
rect 118700 492464 118752 492516
rect 119252 492464 119304 492516
rect 120080 492464 120132 492516
rect 120540 492464 120592 492516
rect 122932 492464 122984 492516
rect 123300 492464 123352 492516
rect 124312 492464 124364 492516
rect 124956 492464 125008 492516
rect 125692 492464 125744 492516
rect 125876 492464 125928 492516
rect 126980 492464 127032 492516
rect 127164 492464 127216 492516
rect 129740 492464 129792 492516
rect 130660 492464 130712 492516
rect 131120 492464 131172 492516
rect 131580 492464 131632 492516
rect 133972 492464 134024 492516
rect 134708 492464 134760 492516
rect 135352 492464 135404 492516
rect 135996 492464 136048 492516
rect 138020 492464 138072 492516
rect 138664 492464 138716 492516
rect 139400 492464 139452 492516
rect 140044 492464 140096 492516
rect 140964 492464 141016 492516
rect 141700 492464 141752 492516
rect 143540 492464 143592 492516
rect 143908 492464 143960 492516
rect 146300 492464 146352 492516
rect 147036 492464 147088 492516
rect 150440 492464 150492 492516
rect 151544 492464 151596 492516
rect 50528 492396 50580 492448
rect 62028 492328 62080 492380
rect 62764 492328 62816 492380
rect 64880 492328 64932 492380
rect 65524 492328 65576 492380
rect 56416 492260 56468 492312
rect 63040 492260 63092 492312
rect 67732 492396 67784 492448
rect 68192 492396 68244 492448
rect 68284 492396 68336 492448
rect 67640 492328 67692 492380
rect 67916 492328 67968 492380
rect 68376 492328 68428 492380
rect 71780 492396 71832 492448
rect 72148 492396 72200 492448
rect 72516 492396 72568 492448
rect 106280 492396 106332 492448
rect 122840 492396 122892 492448
rect 123668 492396 123720 492448
rect 125600 492396 125652 492448
rect 126336 492396 126388 492448
rect 131212 492396 131264 492448
rect 132132 492396 132184 492448
rect 68928 492260 68980 492312
rect 104624 492328 104676 492380
rect 156696 492600 156748 492652
rect 212816 492600 212868 492652
rect 248604 492668 248656 492720
rect 255320 492600 255372 492652
rect 256332 492600 256384 492652
rect 155316 492532 155368 492584
rect 211160 492532 211212 492584
rect 219532 492532 219584 492584
rect 240048 492532 240100 492584
rect 157340 492464 157392 492516
rect 158076 492464 158128 492516
rect 160100 492464 160152 492516
rect 160652 492464 160704 492516
rect 153108 492396 153160 492448
rect 160836 492396 160888 492448
rect 200856 492328 200908 492380
rect 104900 492260 104952 492312
rect 151452 492260 151504 492312
rect 191104 492260 191156 492312
rect 201592 492464 201644 492516
rect 202052 492464 202104 492516
rect 202972 492464 203024 492516
rect 203892 492464 203944 492516
rect 208492 492464 208544 492516
rect 208676 492464 208728 492516
rect 209872 492464 209924 492516
rect 210516 492464 210568 492516
rect 212724 492464 212776 492516
rect 213460 492464 213512 492516
rect 215300 492464 215352 492516
rect 216220 492464 216272 492516
rect 218060 492464 218112 492516
rect 218796 492464 218848 492516
rect 223580 492464 223632 492516
rect 223764 492464 223816 492516
rect 255412 492532 255464 492584
rect 255780 492532 255832 492584
rect 258172 492668 258224 492720
rect 258908 492668 258960 492720
rect 262404 492668 262456 492720
rect 262588 492668 262640 492720
rect 283012 492668 283064 492720
rect 283564 492668 283616 492720
rect 291200 492668 291252 492720
rect 291936 492668 291988 492720
rect 295340 492668 295392 492720
rect 295892 492668 295944 492720
rect 256700 492600 256752 492652
rect 257068 492600 257120 492652
rect 258080 492600 258132 492652
rect 258540 492600 258592 492652
rect 259460 492600 259512 492652
rect 260196 492600 260248 492652
rect 260840 492600 260892 492652
rect 261484 492600 261536 492652
rect 262220 492600 262272 492652
rect 262864 492600 262916 492652
rect 264980 492600 265032 492652
rect 265900 492600 265952 492652
rect 267832 492600 267884 492652
rect 268660 492600 268712 492652
rect 269120 492600 269172 492652
rect 269948 492600 270000 492652
rect 270592 492600 270644 492652
rect 271236 492600 271288 492652
rect 271972 492600 272024 492652
rect 272524 492600 272576 492652
rect 282920 492600 282972 492652
rect 283196 492600 283248 492652
rect 284300 492600 284352 492652
rect 284852 492600 284904 492652
rect 285680 492600 285732 492652
rect 286692 492600 286744 492652
rect 288440 492600 288492 492652
rect 289268 492600 289320 492652
rect 291292 492600 291344 492652
rect 291476 492600 291528 492652
rect 295524 492600 295576 492652
rect 296260 492600 296312 492652
rect 296720 492600 296772 492652
rect 297732 492600 297784 492652
rect 298192 492600 298244 492652
rect 299020 492600 299072 492652
rect 356796 492532 356848 492584
rect 358360 492464 358412 492516
rect 208400 492396 208452 492448
rect 209136 492396 209188 492448
rect 220912 492396 220964 492448
rect 221464 492396 221516 492448
rect 239680 492396 239732 492448
rect 358268 492396 358320 492448
rect 205732 492328 205784 492380
rect 206376 492328 206428 492380
rect 209228 492328 209280 492380
rect 219992 492328 220044 492380
rect 222660 492328 222712 492380
rect 240784 492328 240836 492380
rect 362316 492328 362368 492380
rect 201776 492260 201828 492312
rect 240600 492260 240652 492312
rect 366548 492260 366600 492312
rect 57244 492192 57296 492244
rect 102416 492192 102468 492244
rect 121460 492192 121512 492244
rect 121920 492192 121972 492244
rect 155224 492192 155276 492244
rect 200672 492192 200724 492244
rect 53380 492124 53432 492176
rect 100208 492124 100260 492176
rect 152280 492124 152332 492176
rect 160836 492124 160888 492176
rect 160928 492124 160980 492176
rect 190184 492124 190236 492176
rect 49148 492056 49200 492108
rect 97540 492056 97592 492108
rect 110144 492056 110196 492108
rect 162124 492056 162176 492108
rect 164148 492056 164200 492108
rect 194968 492124 195020 492176
rect 196992 492124 197044 492176
rect 218336 492124 218388 492176
rect 226156 492192 226208 492244
rect 231400 492192 231452 492244
rect 358176 492192 358228 492244
rect 226064 492124 226116 492176
rect 356704 492124 356756 492176
rect 202144 492056 202196 492108
rect 202788 492056 202840 492108
rect 212080 492056 212132 492108
rect 231768 492056 231820 492108
rect 366364 492056 366416 492108
rect 62856 491988 62908 492040
rect 129648 491988 129700 492040
rect 139860 491988 139912 492040
rect 190092 491988 190144 492040
rect 190184 491988 190236 492040
rect 197636 491988 197688 492040
rect 200304 491988 200356 492040
rect 217416 491988 217468 492040
rect 225604 491988 225656 492040
rect 362224 491988 362276 492040
rect 43904 491920 43956 491972
rect 95332 491920 95384 491972
rect 110328 491920 110380 491972
rect 192484 491920 192536 491972
rect 194508 491920 194560 491972
rect 212448 491920 212500 491972
rect 223488 491920 223540 491972
rect 363604 491920 363656 491972
rect 55036 491852 55088 491904
rect 81716 491852 81768 491904
rect 157984 491852 158036 491904
rect 197360 491852 197412 491904
rect 253940 491852 253992 491904
rect 254216 491852 254268 491904
rect 256792 491852 256844 491904
rect 257620 491852 257672 491904
rect 53748 491784 53800 491836
rect 74540 491784 74592 491836
rect 153936 491784 153988 491836
rect 160928 491784 160980 491836
rect 169760 491784 169812 491836
rect 170036 491784 170088 491836
rect 52368 491716 52420 491768
rect 71964 491716 72016 491768
rect 166908 491716 166960 491768
rect 198096 491784 198148 491836
rect 292580 491784 292632 491836
rect 292764 491784 292816 491836
rect 183468 491716 183520 491768
rect 198188 491716 198240 491768
rect 253940 491716 253992 491768
rect 254860 491716 254912 491768
rect 56508 491648 56560 491700
rect 73804 491648 73856 491700
rect 191104 491648 191156 491700
rect 197728 491648 197780 491700
rect 207204 491648 207256 491700
rect 207756 491648 207808 491700
rect 190092 491580 190144 491632
rect 193864 491580 193916 491632
rect 204168 491376 204220 491428
rect 211620 491376 211672 491428
rect 199016 491308 199068 491360
rect 202420 491308 202472 491360
rect 142160 491240 142212 491292
rect 142620 491240 142672 491292
rect 267096 490764 267148 490816
rect 359464 490764 359516 490816
rect 70400 490696 70452 490748
rect 70860 490696 70912 490748
rect 260932 490696 260984 490748
rect 368112 490696 368164 490748
rect 246488 490628 246540 490680
rect 376116 490628 376168 490680
rect 58992 490560 59044 490612
rect 96252 490560 96304 490612
rect 191840 490560 191892 490612
rect 192392 490560 192444 490612
rect 222568 490560 222620 490612
rect 376024 490560 376076 490612
rect 85764 490424 85816 490476
rect 85948 490424 86000 490476
rect 87052 490424 87104 490476
rect 87604 490424 87656 490476
rect 237472 490424 237524 490476
rect 237748 490424 237800 490476
rect 274824 490424 274876 490476
rect 275192 490424 275244 490476
rect 276020 490424 276072 490476
rect 276940 490424 276992 490476
rect 80060 490356 80112 490408
rect 80980 490356 81032 490408
rect 81532 490356 81584 490408
rect 82268 490356 82320 490408
rect 82820 490356 82872 490408
rect 83556 490356 83608 490408
rect 84292 490356 84344 490408
rect 84936 490356 84988 490408
rect 85580 490356 85632 490408
rect 86316 490356 86368 490408
rect 86960 490356 87012 490408
rect 87236 490356 87288 490408
rect 111892 490356 111944 490408
rect 112628 490356 112680 490408
rect 186320 490356 186372 490408
rect 187148 490356 187200 490408
rect 192116 490356 192168 490408
rect 192852 490356 192904 490408
rect 193220 490356 193272 490408
rect 193772 490356 193824 490408
rect 194600 490356 194652 490408
rect 195428 490356 195480 490408
rect 231860 490356 231912 490408
rect 232412 490356 232464 490408
rect 233240 490356 233292 490408
rect 234252 490356 234304 490408
rect 237380 490356 237432 490408
rect 238208 490356 238260 490408
rect 242900 490356 242952 490408
rect 243452 490356 243504 490408
rect 244372 490356 244424 490408
rect 245292 490356 245344 490408
rect 245660 490356 245712 490408
rect 246580 490356 246632 490408
rect 249800 490356 249852 490408
rect 250536 490356 250588 490408
rect 273260 490356 273312 490408
rect 273812 490356 273864 490408
rect 274640 490356 274692 490408
rect 275652 490356 275704 490408
rect 276112 490356 276164 490408
rect 276572 490356 276624 490408
rect 277492 490356 277544 490408
rect 278228 490356 278280 490408
rect 280160 490356 280212 490408
rect 280988 490356 281040 490408
rect 60740 490288 60792 490340
rect 61108 490288 61160 490340
rect 187700 490152 187752 490204
rect 188436 490152 188488 490204
rect 244648 490152 244700 490204
rect 244556 489948 244608 490000
rect 50344 489812 50396 489864
rect 98092 489812 98144 489864
rect 59820 489744 59872 489796
rect 118700 489744 118752 489796
rect 48228 489676 48280 489728
rect 111248 489676 111300 489728
rect 48044 489608 48096 489660
rect 112076 489608 112128 489660
rect 46572 489540 46624 489592
rect 111708 489540 111760 489592
rect 46296 489472 46348 489524
rect 110788 489472 110840 489524
rect 138204 489472 138256 489524
rect 200304 489472 200356 489524
rect 51724 489404 51776 489456
rect 116032 489404 116084 489456
rect 136732 489404 136784 489456
rect 198924 489404 198976 489456
rect 48964 489336 49016 489388
rect 115204 489336 115256 489388
rect 138112 489336 138164 489388
rect 200396 489336 200448 489388
rect 281816 489336 281868 489388
rect 359556 489336 359608 489388
rect 57152 489268 57204 489320
rect 132500 489268 132552 489320
rect 135444 489268 135496 489320
rect 203248 489268 203300 489320
rect 247316 489268 247368 489320
rect 370596 489268 370648 489320
rect 48688 489200 48740 489252
rect 129740 489200 129792 489252
rect 136824 489200 136876 489252
rect 205824 489200 205876 489252
rect 236736 489200 236788 489252
rect 366456 489200 366508 489252
rect 61936 489132 61988 489184
rect 180064 489132 180116 489184
rect 204352 489132 204404 489184
rect 217324 489132 217376 489184
rect 239312 489132 239364 489184
rect 376208 489132 376260 489184
rect 50436 489064 50488 489116
rect 98000 489064 98052 489116
rect 54668 488996 54720 489048
rect 96712 488996 96764 489048
rect 55772 488928 55824 488980
rect 96804 488928 96856 488980
rect 283104 487840 283156 487892
rect 359832 487840 359884 487892
rect 57704 487772 57756 487824
rect 114284 487772 114336 487824
rect 158904 487772 158956 487824
rect 218796 487772 218848 487824
rect 227628 487772 227680 487824
rect 227812 487772 227864 487824
rect 244464 487772 244516 487824
rect 244740 487772 244792 487824
rect 260932 487772 260984 487824
rect 366732 487772 366784 487824
rect 226432 487296 226484 487348
rect 226708 487296 226760 487348
rect 53196 487092 53248 487144
rect 116952 487092 117004 487144
rect 53288 487024 53340 487076
rect 116492 487024 116544 487076
rect 58624 486956 58676 487008
rect 121552 486956 121604 487008
rect 59728 486888 59780 486940
rect 130016 486888 130068 486940
rect 46664 486820 46716 486872
rect 117412 486820 117464 486872
rect 229192 486820 229244 486872
rect 229836 486820 229888 486872
rect 46388 486752 46440 486804
rect 117872 486752 117924 486804
rect 189080 486752 189132 486804
rect 189724 486752 189776 486804
rect 226340 486752 226392 486804
rect 227260 486752 227312 486804
rect 46480 486684 46532 486736
rect 118240 486684 118292 486736
rect 54392 486616 54444 486668
rect 129924 486616 129976 486668
rect 50804 486548 50856 486600
rect 131304 486548 131356 486600
rect 47952 486480 48004 486532
rect 128544 486480 128596 486532
rect 242072 486480 242124 486532
rect 370688 486480 370740 486532
rect 47860 486412 47912 486464
rect 129832 486412 129884 486464
rect 223672 486412 223724 486464
rect 363696 486412 363748 486464
rect 58900 486344 58952 486396
rect 118792 486344 118844 486396
rect 58808 486276 58860 486328
rect 118884 486276 118936 486328
rect 57888 486208 57940 486260
rect 113916 486208 113968 486260
rect 256884 485188 256936 485240
rect 369308 485188 369360 485240
rect 243084 485120 243136 485172
rect 371976 485120 372028 485172
rect 165712 485052 165764 485104
rect 209044 485052 209096 485104
rect 229284 485052 229336 485104
rect 364984 485052 365036 485104
rect 57060 484304 57112 484356
rect 128452 484304 128504 484356
rect 58716 484236 58768 484288
rect 134064 484236 134116 484288
rect 48780 484168 48832 484220
rect 124220 484168 124272 484220
rect 59636 484100 59688 484152
rect 135352 484100 135404 484152
rect 45468 484032 45520 484084
rect 124312 484032 124364 484084
rect 43628 483964 43680 484016
rect 122932 483964 122984 484016
rect 42248 483896 42300 483948
rect 124404 483896 124456 483948
rect 48872 483828 48924 483880
rect 132684 483828 132736 483880
rect 46112 483760 46164 483812
rect 132592 483760 132644 483812
rect 43352 483692 43404 483744
rect 131212 483692 131264 483744
rect 292764 483692 292816 483744
rect 379980 483692 380032 483744
rect 46020 483624 46072 483676
rect 143632 483624 143684 483676
rect 167184 483624 167236 483676
rect 215944 483624 215996 483676
rect 237564 483624 237616 483676
rect 378876 483624 378928 483676
rect 58532 483556 58584 483608
rect 128360 483556 128412 483608
rect 59360 483488 59412 483540
rect 86224 483488 86276 483540
rect 262404 482400 262456 482452
rect 373448 482400 373500 482452
rect 205640 482332 205692 482384
rect 217600 482332 217652 482384
rect 236000 482332 236052 482384
rect 367836 482332 367888 482384
rect 57612 482264 57664 482316
rect 114560 482264 114612 482316
rect 168564 482264 168616 482316
rect 210424 482264 210476 482316
rect 229100 482264 229152 482316
rect 360936 482264 360988 482316
rect 295616 481108 295668 481160
rect 376760 481108 376812 481160
rect 242992 481040 243044 481092
rect 363788 481040 363840 481092
rect 149060 480972 149112 481024
rect 211804 480972 211856 481024
rect 254216 480972 254268 481024
rect 379060 480972 379112 481024
rect 60832 480904 60884 480956
rect 199200 480904 199252 480956
rect 230480 480904 230532 480956
rect 365076 480904 365128 480956
rect 296904 480156 296956 480208
rect 358636 480156 358688 480208
rect 295432 480088 295484 480140
rect 362684 480088 362736 480140
rect 295340 480020 295392 480072
rect 364156 480020 364208 480072
rect 295524 479952 295576 480004
rect 366916 479952 366968 480004
rect 294144 479884 294196 479936
rect 365628 479884 365680 479936
rect 296812 479816 296864 479868
rect 369584 479816 369636 479868
rect 298284 479748 298336 479800
rect 379520 479748 379572 479800
rect 287244 479680 287296 479732
rect 373724 479680 373776 479732
rect 284484 479612 284536 479664
rect 377404 479612 377456 479664
rect 178224 479544 178276 479596
rect 210608 479544 210660 479596
rect 252744 479544 252796 479596
rect 374828 479544 374880 479596
rect 161756 479476 161808 479528
rect 216036 479476 216088 479528
rect 244556 479476 244608 479528
rect 369124 479476 369176 479528
rect 256792 478252 256844 478304
rect 361304 478252 361356 478304
rect 252652 478184 252704 478236
rect 369400 478184 369452 478236
rect 146392 478116 146444 478168
rect 211896 478116 211948 478168
rect 244464 478116 244516 478168
rect 374644 478116 374696 478168
rect 292672 477436 292724 477488
rect 357164 477436 357216 477488
rect 294052 477368 294104 477420
rect 368388 477368 368440 477420
rect 293960 477300 294012 477352
rect 371148 477300 371200 477352
rect 291384 477232 291436 477284
rect 374460 477232 374512 477284
rect 291292 477164 291344 477216
rect 376484 477164 376536 477216
rect 285956 477096 286008 477148
rect 371792 477096 371844 477148
rect 281632 477028 281684 477080
rect 368296 477028 368348 477080
rect 290004 476960 290056 477012
rect 377220 476960 377272 477012
rect 256700 476892 256752 476944
rect 365352 476892 365404 476944
rect 244372 476824 244424 476876
rect 373264 476824 373316 476876
rect 158812 476756 158864 476808
rect 203616 476756 203668 476808
rect 226524 476756 226576 476808
rect 378784 476756 378836 476808
rect 262312 475464 262364 475516
rect 379244 475464 379296 475516
rect 252560 475396 252612 475448
rect 374920 475396 374972 475448
rect 62764 475328 62816 475380
rect 199384 475328 199436 475380
rect 227904 475328 227956 475380
rect 367744 475328 367796 475380
rect 289912 474580 289964 474632
rect 373172 474580 373224 474632
rect 267832 474512 267884 474564
rect 359648 474512 359700 474564
rect 270684 474444 270736 474496
rect 362776 474444 362828 474496
rect 267924 474376 267976 474428
rect 361396 474376 361448 474428
rect 270592 474308 270644 474360
rect 364892 474308 364944 474360
rect 269304 474240 269356 474292
rect 369676 474240 369728 474292
rect 269212 474172 269264 474224
rect 372436 474172 372488 474224
rect 259644 474104 259696 474156
rect 372252 474104 372304 474156
rect 244280 474036 244332 474088
rect 358452 474036 358504 474088
rect 161664 473968 161716 474020
rect 213184 473968 213236 474020
rect 237472 473968 237524 474020
rect 372068 473968 372120 474020
rect 185032 472744 185084 472796
rect 210700 472744 210752 472796
rect 258264 472744 258316 472796
rect 373540 472744 373592 472796
rect 178132 472676 178184 472728
rect 205088 472676 205140 472728
rect 245752 472676 245804 472728
rect 361120 472676 361172 472728
rect 3608 472608 3660 472660
rect 307024 472608 307076 472660
rect 3516 471928 3568 471980
rect 429200 471928 429252 471980
rect 273444 471860 273496 471912
rect 359740 471860 359792 471912
rect 276204 471792 276256 471844
rect 364248 471792 364300 471844
rect 277584 471724 277636 471776
rect 369032 471724 369084 471776
rect 274916 471656 274968 471708
rect 367652 471656 367704 471708
rect 284392 471588 284444 471640
rect 377680 471588 377732 471640
rect 267740 471520 267792 471572
rect 361488 471520 361540 471572
rect 272064 471452 272116 471504
rect 367008 471452 367060 471504
rect 273352 471384 273404 471436
rect 377496 471384 377548 471436
rect 176844 471316 176896 471368
rect 206560 471316 206612 471368
rect 259552 471316 259604 471368
rect 370872 471316 370924 471368
rect 164424 471248 164476 471300
rect 211988 471248 212040 471300
rect 251364 471248 251416 471300
rect 363972 471248 364024 471300
rect 284300 470024 284352 470076
rect 377772 470024 377824 470076
rect 251272 469956 251324 470008
rect 362408 469956 362460 470008
rect 176752 469888 176804 469940
rect 212172 469888 212224 469940
rect 241612 469888 241664 469940
rect 365168 469888 365220 469940
rect 4804 469820 4856 469872
rect 391940 469820 391992 469872
rect 48136 469140 48188 469192
rect 72424 469140 72476 469192
rect 285864 469140 285916 469192
rect 370412 469140 370464 469192
rect 42616 469072 42668 469124
rect 67824 469072 67876 469124
rect 266452 469072 266504 469124
rect 360752 469072 360804 469124
rect 42524 469004 42576 469056
rect 70584 469004 70636 469056
rect 276112 469004 276164 469056
rect 375104 469004 375156 469056
rect 42432 468936 42484 468988
rect 94044 468936 94096 468988
rect 259460 468936 259512 468988
rect 362500 468936 362552 468988
rect 46204 468868 46256 468920
rect 104992 468868 105044 468920
rect 254032 468868 254084 468920
rect 362592 468868 362644 468920
rect 43536 468800 43588 468852
rect 103612 468800 103664 468852
rect 255320 468800 255372 468852
rect 365444 468800 365496 468852
rect 42156 468732 42208 468784
rect 102232 468732 102284 468784
rect 254124 468732 254176 468784
rect 368204 468732 368256 468784
rect 45376 468664 45428 468716
rect 106372 468664 106424 468716
rect 255504 468664 255556 468716
rect 373632 468664 373684 468716
rect 45284 468596 45336 468648
rect 106464 468596 106516 468648
rect 255412 468596 255464 468648
rect 376300 468596 376352 468648
rect 43444 468528 43496 468580
rect 105084 468528 105136 468580
rect 174084 468528 174136 468580
rect 214656 468528 214708 468580
rect 247132 468528 247184 468580
rect 378968 468528 379020 468580
rect 18604 468460 18656 468512
rect 378140 468460 378192 468512
rect 44088 468392 44140 468444
rect 66352 468392 66404 468444
rect 288624 468392 288676 468444
rect 367560 468392 367612 468444
rect 175464 467236 175516 467288
rect 200856 467236 200908 467288
rect 175372 467168 175424 467220
rect 202236 467168 202288 467220
rect 57520 467100 57572 467152
rect 111892 467100 111944 467152
rect 162952 467100 163004 467152
rect 209136 467100 209188 467152
rect 209228 467100 209280 467152
rect 217784 467100 217836 467152
rect 227812 467100 227864 467152
rect 371884 467100 371936 467152
rect 45192 466352 45244 466404
rect 68284 466352 68336 466404
rect 190644 466352 190696 466404
rect 212908 466352 212960 466404
rect 280344 466352 280396 466404
rect 357256 466352 357308 466404
rect 45100 466284 45152 466336
rect 68376 466284 68428 466336
rect 176660 466284 176712 466336
rect 209320 466284 209372 466336
rect 298192 466284 298244 466336
rect 376576 466284 376628 466336
rect 52092 466216 52144 466268
rect 82820 466216 82872 466268
rect 173992 466216 174044 466268
rect 207848 466216 207900 466268
rect 289820 466216 289872 466268
rect 373080 466216 373132 466268
rect 50712 466148 50764 466200
rect 83004 466148 83056 466200
rect 140780 466148 140832 466200
rect 197820 466148 197872 466200
rect 271972 466148 272024 466200
rect 358728 466148 358780 466200
rect 49516 466080 49568 466132
rect 82912 466080 82964 466132
rect 139400 466080 139452 466132
rect 197084 466080 197136 466132
rect 263784 466080 263836 466132
rect 356888 466080 356940 466132
rect 57796 466012 57848 466064
rect 102324 466012 102376 466064
rect 140872 466012 140924 466064
rect 200488 466012 200540 466064
rect 263692 466012 263744 466064
rect 366824 466012 366876 466064
rect 54576 465944 54628 465996
rect 100944 465944 100996 465996
rect 140964 465944 141016 465996
rect 201776 465944 201828 465996
rect 265256 465944 265308 465996
rect 372344 465944 372396 465996
rect 53104 465876 53156 465928
rect 100852 465876 100904 465928
rect 141056 465876 141108 465928
rect 203340 465876 203392 465928
rect 265164 465876 265216 465928
rect 375012 465876 375064 465928
rect 57428 465808 57480 465860
rect 113364 465808 113416 465860
rect 139492 465808 139544 465860
rect 204536 465808 204588 465860
rect 260840 465808 260892 465860
rect 376392 465808 376444 465860
rect 50252 465740 50304 465792
rect 98184 465740 98236 465792
rect 107844 465740 107896 465792
rect 204352 465740 204404 465792
rect 226340 465740 226392 465792
rect 361028 465740 361080 465792
rect 51632 465672 51684 465724
rect 99472 465672 99524 465724
rect 109040 465672 109092 465724
rect 205640 465672 205692 465724
rect 227720 465672 227772 465724
rect 370504 465672 370556 465724
rect 44732 465604 44784 465656
rect 65064 465604 65116 465656
rect 187884 465604 187936 465656
rect 206652 465604 206704 465656
rect 44824 465536 44876 465588
rect 64972 465536 65024 465588
rect 182364 465536 182416 465588
rect 200948 465536 201000 465588
rect 44916 465468 44968 465520
rect 64880 465468 64932 465520
rect 192116 465468 192168 465520
rect 205364 465468 205416 465520
rect 287152 464448 287204 464500
rect 370320 464448 370372 464500
rect 164240 464380 164292 464432
rect 216128 464380 216180 464432
rect 274824 464380 274876 464432
rect 364800 464380 364852 464432
rect 160192 464312 160244 464364
rect 214564 464312 214616 464364
rect 285772 464312 285824 464364
rect 377588 464312 377640 464364
rect 59912 463632 59964 463684
rect 91192 463632 91244 463684
rect 190552 463632 190604 463684
rect 214380 463632 214432 463684
rect 54944 463564 54996 463616
rect 86960 463564 87012 463616
rect 190460 463564 190512 463616
rect 217508 463564 217560 463616
rect 277492 463564 277544 463616
rect 357348 463564 357400 463616
rect 49608 463496 49660 463548
rect 81624 463496 81676 463548
rect 184940 463496 184992 463548
rect 213276 463496 213328 463548
rect 288532 463496 288584 463548
rect 368940 463496 368992 463548
rect 55956 463428 56008 463480
rect 88616 463428 88668 463480
rect 183744 463428 183796 463480
rect 212264 463428 212316 463480
rect 277400 463428 277452 463480
rect 366272 463428 366324 463480
rect 52000 463360 52052 463412
rect 85672 463360 85724 463412
rect 175280 463360 175332 463412
rect 207940 463360 207992 463412
rect 276020 463360 276072 463412
rect 371700 463360 371752 463412
rect 56232 463292 56284 463344
rect 89812 463292 89864 463344
rect 180984 463292 181036 463344
rect 216220 463292 216272 463344
rect 269120 463292 269172 463344
rect 366180 463292 366232 463344
rect 54852 463224 54904 463276
rect 88524 463224 88576 463276
rect 160100 463224 160152 463276
rect 200764 463224 200816 463276
rect 263600 463224 263652 463276
rect 363880 463224 363932 463276
rect 54760 463156 54812 463208
rect 88432 463156 88484 463208
rect 168472 463156 168524 463208
rect 210516 463156 210568 463208
rect 262220 463156 262272 463208
rect 365536 463156 365588 463208
rect 53012 463088 53064 463140
rect 87144 463088 87196 463140
rect 142344 463088 142396 463140
rect 199108 463088 199160 463140
rect 241520 463088 241572 463140
rect 358544 463088 358596 463140
rect 59084 463020 59136 463072
rect 95424 463020 95476 463072
rect 142252 463020 142304 463072
rect 207480 463020 207532 463072
rect 251180 463020 251232 463072
rect 370780 463020 370832 463072
rect 52828 462952 52880 463004
rect 100760 462952 100812 463004
rect 107752 462952 107804 463004
rect 197636 462952 197688 463004
rect 240140 462952 240192 463004
rect 361212 462952 361264 463004
rect 56048 462884 56100 462936
rect 87052 462884 87104 462936
rect 180892 462884 180944 462936
rect 203708 462884 203760 462936
rect 55864 462816 55916 462868
rect 85580 462816 85632 462868
rect 187792 462816 187844 462868
rect 205180 462816 205232 462868
rect 44640 462748 44692 462800
rect 63684 462748 63736 462800
rect 193312 462748 193364 462800
rect 206836 462748 206888 462800
rect 207020 462340 207072 462392
rect 207296 462340 207348 462392
rect 217692 462340 217744 462392
rect 86224 462272 86276 462324
rect 178316 462272 178368 462324
rect 180064 462272 180116 462324
rect 199568 462272 199620 462324
rect 203156 462272 203208 462324
rect 206284 462272 206336 462324
rect 192484 462204 192536 462256
rect 210056 462204 210108 462256
rect 186412 462136 186464 462188
rect 205272 462136 205324 462188
rect 191932 462068 191984 462120
rect 215852 462068 215904 462120
rect 283012 462068 283064 462120
rect 360844 462068 360896 462120
rect 192024 462000 192076 462052
rect 218428 462000 218480 462052
rect 278780 462000 278832 462052
rect 357900 462000 357952 462052
rect 182272 461932 182324 461984
rect 209412 461932 209464 461984
rect 287060 461932 287112 461984
rect 372528 461932 372580 461984
rect 182180 461864 182232 461916
rect 211436 461864 211488 461916
rect 285680 461864 285732 461916
rect 374000 461864 374052 461916
rect 511264 461864 511316 461916
rect 517520 461864 517572 461916
rect 171232 461796 171284 461848
rect 212080 461796 212132 461848
rect 271880 461796 271932 461848
rect 363512 461796 363564 461848
rect 57336 461728 57388 461780
rect 111984 461728 112036 461780
rect 165620 461728 165672 461780
rect 218888 461728 218940 461780
rect 280252 461728 280304 461780
rect 375748 461728 375800 461780
rect 62212 461660 62264 461712
rect 199476 461660 199528 461712
rect 199568 461660 199620 461712
rect 339684 461660 339736 461712
rect 47584 461592 47636 461644
rect 207020 461592 207072 461644
rect 274732 461592 274784 461644
rect 371056 461592 371108 461644
rect 339684 461048 339736 461100
rect 360108 461048 360160 461100
rect 499856 461048 499908 461100
rect 500868 461048 500920 461100
rect 178316 460980 178368 461032
rect 200580 460980 200632 461032
rect 338304 460980 338356 461032
rect 357072 460980 357124 461032
rect 498476 460980 498528 461032
rect 517796 460980 517848 461032
rect 190920 460912 190972 460964
rect 207020 460912 207072 460964
rect 351000 460912 351052 460964
rect 361580 460912 361632 460964
rect 500868 460912 500920 460964
rect 517612 460912 517664 460964
rect 49240 460844 49292 460896
rect 78864 460844 78916 460896
rect 183560 460844 183612 460896
rect 202328 460844 202380 460896
rect 299480 460844 299532 460896
rect 379428 460844 379480 460896
rect 50988 460776 51040 460828
rect 78680 460776 78732 460828
rect 193864 460776 193916 460828
rect 213000 460776 213052 460828
rect 266360 460776 266412 460828
rect 358084 460776 358136 460828
rect 53472 460708 53524 460760
rect 77300 460708 77352 460760
rect 189264 460708 189316 460760
rect 210240 460708 210292 460760
rect 281540 460708 281592 460760
rect 379336 460708 379388 460760
rect 52276 460640 52328 460692
rect 75920 460640 75972 460692
rect 172612 460640 172664 460692
rect 207756 460640 207808 460692
rect 258080 460640 258132 460692
rect 364064 460640 364116 460692
rect 55496 460572 55548 460624
rect 78772 460572 78824 460624
rect 179512 460572 179564 460624
rect 214748 460572 214800 460624
rect 248420 460572 248472 460624
rect 366640 460572 366692 460624
rect 55128 460504 55180 460556
rect 71872 460504 71924 460556
rect 179420 460504 179472 460556
rect 214840 460504 214892 460556
rect 249800 460504 249852 460556
rect 368020 460504 368072 460556
rect 52368 460436 52420 460488
rect 70400 460436 70452 460488
rect 162124 460436 162176 460488
rect 197728 460436 197780 460488
rect 249984 460436 250036 460488
rect 369216 460436 369268 460488
rect 43996 460368 44048 460420
rect 67640 460368 67692 460420
rect 167092 460368 167144 460420
rect 204996 460368 205048 460420
rect 242900 460368 242952 460420
rect 365260 460368 365312 460420
rect 51908 460300 51960 460352
rect 92572 460300 92624 460352
rect 168380 460300 168432 460352
rect 206376 460300 206428 460352
rect 249892 460300 249944 460352
rect 373356 460300 373408 460352
rect 45008 460232 45060 460284
rect 103704 460232 103756 460284
rect 125600 460232 125652 460284
rect 196900 460232 196952 460284
rect 248512 460232 248564 460284
rect 372160 460232 372212 460284
rect 47676 460164 47728 460216
rect 63500 460164 63552 460216
rect 63592 460164 63644 460216
rect 199016 460164 199068 460216
rect 237380 460164 237432 460216
rect 374736 460164 374788 460216
rect 50160 460096 50212 460148
rect 66260 460096 66312 460148
rect 187700 460096 187752 460148
rect 203800 460096 203852 460148
rect 280160 460096 280212 460148
rect 357992 460096 358044 460148
rect 47768 460028 47820 460080
rect 62120 460028 62172 460080
rect 193220 460028 193272 460080
rect 208860 460028 208912 460080
rect 194692 459960 194744 460012
rect 203524 459960 203576 460012
rect 214288 459620 214340 459672
rect 220912 459620 220964 459672
rect 216312 459552 216364 459604
rect 220820 459552 220872 459604
rect 191840 459484 191892 459536
rect 208032 459484 208084 459536
rect 194600 459416 194652 459468
rect 211528 459416 211580 459468
rect 291200 459416 291252 459468
rect 360660 459416 360712 459468
rect 189172 459348 189224 459400
rect 209504 459348 209556 459400
rect 282920 459348 282972 459400
rect 359924 459348 359976 459400
rect 180800 459280 180852 459332
rect 210792 459280 210844 459332
rect 288440 459280 288492 459332
rect 374552 459280 374604 459332
rect 59176 459212 59228 459264
rect 92480 459212 92532 459264
rect 173900 459212 173952 459264
rect 206744 459212 206796 459264
rect 274640 459212 274692 459264
rect 362868 459212 362920 459264
rect 51540 459144 51592 459196
rect 99564 459144 99616 459196
rect 178040 459144 178092 459196
rect 218980 459144 219032 459196
rect 270500 459144 270552 459196
rect 363420 459144 363472 459196
rect 52736 459076 52788 459128
rect 120080 459076 120132 459128
rect 142160 459076 142212 459128
rect 198004 459076 198056 459128
rect 273260 459076 273312 459128
rect 372988 459076 373040 459128
rect 54300 459008 54352 459060
rect 131120 459008 131172 459060
rect 136640 459008 136692 459060
rect 199292 459008 199344 459060
rect 264980 459008 265032 459060
rect 369492 459008 369544 459060
rect 56232 458940 56284 458992
rect 133972 458940 134024 458992
rect 135260 458940 135312 458992
rect 197912 458940 197964 458992
rect 253940 458940 253992 458992
rect 370964 458940 371016 458992
rect 52276 458872 52328 458924
rect 133880 458872 133932 458924
rect 138020 458872 138072 458924
rect 201868 458872 201920 458924
rect 247040 458872 247092 458924
rect 367928 458872 367980 458924
rect 60740 458804 60792 458856
rect 199568 458804 199620 458856
rect 245660 458804 245712 458856
rect 379152 458804 379204 458856
rect 189080 458736 189132 458788
rect 201040 458736 201092 458788
rect 199016 458328 199068 458380
rect 47492 458260 47544 458312
rect 358820 458260 358872 458312
rect 516600 458260 516652 458312
rect 207388 458192 207440 458244
rect 208124 458192 208176 458244
rect 53012 457784 53064 457836
rect 53472 457784 53524 457836
rect 49240 456084 49292 456136
rect 49608 456084 49660 456136
rect 518164 441532 518216 441584
rect 579896 441532 579948 441584
rect 3148 422220 3200 422272
rect 18604 422220 18656 422272
rect 54484 416644 54536 416696
rect 57244 416644 57296 416696
rect 56232 415352 56284 415404
rect 56600 415352 56652 415404
rect 47584 412564 47636 412616
rect 57244 412564 57296 412616
rect 47492 411204 47544 411256
rect 57244 411204 57296 411256
rect 50804 411068 50856 411120
rect 55680 411068 55732 411120
rect 208124 410524 208176 410576
rect 216772 410524 216824 410576
rect 205732 409096 205784 409148
rect 216772 409096 216824 409148
rect 56232 408552 56284 408604
rect 56600 408552 56652 408604
rect 57060 408552 57112 408604
rect 57980 408552 58032 408604
rect 47584 408484 47636 408536
rect 57244 408484 57296 408536
rect 58532 407736 58584 407788
rect 59360 407736 59412 407788
rect 57060 407464 57112 407516
rect 59636 407464 59688 407516
rect 47492 407124 47544 407176
rect 57244 407124 57296 407176
rect 360844 406376 360896 406428
rect 377404 406376 377456 406428
rect 47400 405696 47452 405748
rect 57244 405696 57296 405748
rect 204444 404948 204496 405000
rect 216864 404948 216916 405000
rect 359924 404948 359976 405000
rect 377680 404948 377732 405000
rect 50804 404336 50856 404388
rect 57244 404336 57296 404388
rect 359832 403588 359884 403640
rect 377772 403588 377824 403640
rect 50988 402976 51040 403028
rect 57244 402976 57296 403028
rect 360108 389308 360160 389360
rect 361672 389308 361724 389360
rect 46020 384956 46072 385008
rect 57244 384956 57296 385008
rect 206284 384956 206336 385008
rect 216680 384956 216732 385008
rect 359556 384956 359608 385008
rect 376944 384956 376996 385008
rect 47952 383596 48004 383648
rect 56876 383596 56928 383648
rect 207020 383596 207072 383648
rect 216680 383596 216732 383648
rect 361580 383596 361632 383648
rect 376944 383596 376996 383648
rect 57152 383528 57204 383580
rect 57612 383528 57664 383580
rect 209504 383528 209556 383580
rect 217048 383528 217100 383580
rect 359464 383528 359516 383580
rect 376852 383528 376904 383580
rect 56968 382304 57020 382356
rect 57244 382304 57296 382356
rect 206284 382236 206336 382288
rect 207020 382236 207072 382288
rect 360844 382236 360896 382288
rect 361580 382236 361632 382288
rect 42708 382168 42760 382220
rect 57244 382168 57296 382220
rect 57520 382168 57572 382220
rect 47952 380876 48004 380928
rect 48780 380876 48832 380928
rect 212908 380672 212960 380724
rect 212908 380468 212960 380520
rect 57152 377748 57204 377800
rect 57612 377748 57664 377800
rect 216772 375300 216824 375352
rect 217784 375300 217836 375352
rect 47584 375028 47636 375080
rect 216772 375028 216824 375080
rect 47492 374960 47544 375012
rect 217232 374960 217284 375012
rect 58808 374892 58860 374944
rect 60740 374892 60792 374944
rect 58900 374824 58952 374876
rect 62120 374824 62172 374876
rect 208952 374824 209004 374876
rect 218244 374824 218296 374876
rect 140964 374756 141016 374808
rect 201868 374756 201920 374808
rect 203064 374756 203116 374808
rect 281448 374756 281500 374808
rect 359740 374756 359792 374808
rect 440332 374756 440384 374808
rect 201500 374688 201552 374740
rect 311808 374688 311860 374740
rect 358636 374688 358688 374740
rect 372896 374688 372948 374740
rect 201684 374620 201736 374672
rect 314568 374620 314620 374672
rect 372436 374620 372488 374672
rect 418252 374620 418304 374672
rect 165988 374552 166040 374604
rect 199108 374552 199160 374604
rect 360752 374552 360804 374604
rect 407764 374552 407816 374604
rect 163412 374484 163464 374536
rect 198004 374484 198056 374536
rect 361488 374484 361540 374536
rect 410708 374484 410760 374536
rect 158536 374416 158588 374468
rect 201776 374416 201828 374468
rect 213552 374416 213604 374468
rect 244280 374416 244332 374468
rect 372896 374416 372948 374468
rect 373816 374416 373868 374468
rect 433340 374416 433392 374468
rect 160928 374348 160980 374400
rect 207480 374348 207532 374400
rect 241244 374348 241296 374400
rect 248696 374348 248748 374400
rect 377496 374348 377548 374400
rect 443092 374348 443144 374400
rect 153476 374280 153528 374332
rect 200488 374280 200540 374332
rect 241152 374280 241204 374332
rect 250076 374280 250128 374332
rect 367008 374280 367060 374332
rect 434812 374280 434864 374332
rect 148968 374212 149020 374264
rect 197084 374212 197136 374264
rect 215484 374212 215536 374264
rect 263692 374212 263744 374264
rect 363512 374212 363564 374264
rect 433616 374212 433668 374264
rect 146208 374144 146260 374196
rect 204536 374144 204588 374196
rect 218244 374144 218296 374196
rect 271144 374144 271196 374196
rect 372988 374144 373040 374196
rect 445944 374144 445996 374196
rect 143540 374076 143592 374128
rect 213092 374076 213144 374128
rect 219624 374076 219676 374128
rect 222016 374076 222068 374128
rect 270316 374076 270368 374128
rect 275836 374076 275888 374128
rect 371056 374076 371108 374128
rect 448244 374076 448296 374128
rect 56968 374008 57020 374060
rect 105452 374008 105504 374060
rect 201592 374008 201644 374060
rect 320916 374008 320968 374060
rect 373908 374008 373960 374060
rect 47400 373940 47452 373992
rect 217600 373940 217652 373992
rect 404820 373940 404872 373992
rect 58716 373872 58768 373924
rect 116124 373872 116176 373924
rect 139216 373872 139268 373924
rect 200304 373872 200356 373924
rect 369676 373872 369728 373924
rect 421012 373872 421064 373924
rect 43352 373804 43404 373856
rect 103520 373804 103572 373856
rect 136456 373804 136508 373856
rect 200396 373804 200448 373856
rect 366180 373804 366232 373856
rect 423036 373804 423088 373856
rect 52276 373736 52328 373788
rect 113548 373736 113600 373788
rect 131028 373736 131080 373788
rect 199292 373736 199344 373788
rect 219440 373736 219492 373788
rect 219624 373736 219676 373788
rect 368388 373736 368440 373788
rect 376852 373736 376904 373788
rect 379428 373736 379480 373788
rect 439412 373736 439464 373788
rect 56232 373668 56284 373720
rect 118332 373668 118384 373720
rect 128912 373668 128964 373720
rect 198924 373668 198976 373720
rect 215300 373668 215352 373720
rect 215576 373668 215628 373720
rect 219256 373668 219308 373720
rect 363420 373668 363472 373720
rect 425428 373668 425480 373720
rect 57060 373600 57112 373652
rect 125692 373600 125744 373652
rect 133696 373600 133748 373652
rect 205824 373600 205876 373652
rect 367652 373600 367704 373652
rect 450268 373600 450320 373652
rect 48872 373532 48924 373584
rect 110420 373532 110472 373584
rect 121368 373532 121420 373584
rect 197912 373532 197964 373584
rect 215300 373532 215352 373584
rect 216496 373532 216548 373584
rect 236460 373532 236512 373584
rect 375104 373532 375156 373584
rect 460940 373532 460992 373584
rect 46112 373464 46164 373516
rect 107844 373464 107896 373516
rect 124128 373464 124180 373516
rect 203248 373464 203300 373516
rect 209780 373464 209832 373516
rect 211068 373464 211120 373516
rect 214932 373464 214984 373516
rect 224224 373464 224276 373516
rect 364800 373464 364852 373516
rect 452844 373464 452896 373516
rect 55680 373396 55732 373448
rect 98276 373396 98328 373448
rect 98368 373396 98420 373448
rect 212724 373396 212776 373448
rect 215024 373396 215076 373448
rect 242900 373396 242952 373448
rect 371700 373396 371752 373448
rect 462780 373396 462832 373448
rect 48688 373328 48740 373380
rect 96068 373328 96120 373380
rect 96160 373328 96212 373380
rect 212632 373328 212684 373380
rect 47860 373260 47912 373312
rect 90180 373260 90232 373312
rect 95056 373260 95108 373312
rect 212540 373260 212592 373312
rect 362868 373328 362920 373380
rect 455420 373328 455472 373380
rect 219348 373260 219400 373312
rect 269212 373260 269264 373312
rect 364248 373260 364300 373312
rect 458180 373260 458232 373312
rect 54300 373192 54352 373244
rect 100852 373192 100904 373244
rect 151728 373192 151780 373244
rect 197820 373192 197872 373244
rect 219164 373192 219216 373244
rect 253940 373192 253992 373244
rect 365628 373192 365680 373244
rect 380900 373192 380952 373244
rect 54392 373124 54444 373176
rect 88340 373124 88392 373176
rect 156512 373124 156564 373176
rect 203340 373124 203392 373176
rect 212632 373124 212684 373176
rect 217968 373124 218020 373176
rect 255412 373124 255464 373176
rect 59728 373056 59780 373108
rect 93676 373056 93728 373108
rect 212724 373056 212776 373108
rect 219072 373056 219124 373108
rect 258080 373056 258132 373108
rect 212816 372988 212868 373040
rect 213644 372988 213696 373040
rect 256700 372988 256752 373040
rect 214012 372920 214064 372972
rect 259644 372920 259696 372972
rect 216956 372852 217008 372904
rect 217600 372852 217652 372904
rect 100024 372784 100076 372836
rect 213920 372784 213972 372836
rect 215208 372784 215260 372836
rect 259460 372852 259512 372904
rect 204260 372716 204312 372768
rect 215300 372716 215352 372768
rect 207204 372648 207256 372700
rect 215024 372648 215076 372700
rect 215392 372648 215444 372700
rect 216404 372648 216456 372700
rect 220728 372784 220780 372836
rect 219256 372716 219308 372768
rect 264980 372784 265032 372836
rect 220912 372716 220964 372768
rect 266360 372716 266412 372768
rect 214104 372580 214156 372632
rect 261300 372648 261352 372700
rect 380900 372648 380952 372700
rect 426440 372648 426492 372700
rect 220728 372580 220780 372632
rect 262220 372580 262272 372632
rect 275836 372580 275888 372632
rect 356612 372580 356664 372632
rect 369768 372580 369820 372632
rect 84752 372512 84804 372564
rect 208492 372512 208544 372564
rect 210976 372512 211028 372564
rect 212724 372512 212776 372564
rect 219440 372512 219492 372564
rect 273260 372512 273312 372564
rect 281448 372512 281500 372564
rect 326068 372512 326120 372564
rect 370320 372512 370372 372564
rect 375104 372512 375156 372564
rect 86776 372444 86828 372496
rect 208400 372444 208452 372496
rect 210332 372444 210384 372496
rect 218060 372444 218112 372496
rect 271880 372444 271932 372496
rect 376852 372580 376904 372632
rect 378048 372580 378100 372632
rect 425060 372580 425112 372632
rect 439412 372580 439464 372632
rect 516692 372648 516744 372700
rect 511908 372580 511960 372632
rect 517520 372580 517572 372632
rect 376576 372512 376628 372564
rect 438216 372512 438268 372564
rect 376760 372444 376812 372496
rect 427820 372444 427872 372496
rect 91560 372376 91612 372428
rect 92388 372308 92440 372360
rect 204168 372308 204220 372360
rect 93400 372240 93452 372292
rect 202788 372240 202840 372292
rect 52920 372172 52972 372224
rect 54392 372172 54444 372224
rect 79508 372172 79560 372224
rect 213368 372376 213420 372428
rect 368940 372308 368992 372360
rect 379612 372308 379664 372360
rect 210976 372240 211028 372292
rect 244280 372240 244332 372292
rect 211344 372172 211396 372224
rect 219900 372172 219952 372224
rect 220544 372172 220596 372224
rect 215300 372104 215352 372156
rect 220452 372104 220504 372156
rect 251180 372172 251232 372224
rect 373080 372104 373132 372156
rect 379520 372104 379572 372156
rect 202788 372036 202840 372088
rect 220820 372036 220872 372088
rect 221924 372036 221976 372088
rect 367560 372036 367612 372088
rect 376760 372036 376812 372088
rect 112996 371968 113048 372020
rect 210332 371968 210384 372020
rect 220636 371968 220688 372020
rect 241244 371968 241296 372020
rect 379336 371968 379388 372020
rect 396080 371968 396132 372020
rect 204168 371900 204220 371952
rect 219532 371900 219584 371952
rect 220452 371900 220504 371952
rect 182732 371764 182784 371816
rect 202972 371764 203024 371816
rect 204168 371764 204220 371816
rect 114468 371696 114520 371748
rect 212724 371696 212776 371748
rect 88064 371628 88116 371680
rect 211068 371628 211120 371680
rect 90916 371560 90968 371612
rect 209872 371560 209924 371612
rect 219808 371832 219860 371884
rect 241152 371900 241204 371952
rect 371056 371900 371108 371952
rect 398840 371900 398892 371952
rect 224224 371832 224276 371884
rect 247132 371832 247184 371884
rect 372528 371832 372580 371884
rect 405740 371832 405792 371884
rect 215300 371764 215352 371816
rect 216312 371764 216364 371816
rect 239128 371764 239180 371816
rect 240048 371764 240100 371816
rect 213368 371696 213420 371748
rect 245660 371696 245712 371748
rect 220544 371628 220596 371680
rect 251180 371628 251232 371680
rect 274640 371628 274692 371680
rect 302240 371628 302292 371680
rect 280068 371560 280120 371612
rect 359280 371560 359332 371612
rect 89352 371492 89404 371544
rect 209964 371492 210016 371544
rect 219716 371492 219768 371544
rect 220636 371492 220688 371544
rect 221924 371492 221976 371544
rect 252560 371492 252612 371544
rect 276020 371492 276072 371544
rect 356980 371492 357032 371544
rect 44640 371424 44692 371476
rect 47492 371424 47544 371476
rect 78312 371424 78364 371476
rect 369676 371764 369728 371816
rect 397460 371764 397512 371816
rect 379612 371696 379664 371748
rect 379796 371696 379848 371748
rect 409880 371696 409932 371748
rect 374552 371628 374604 371680
rect 380072 371628 380124 371680
rect 411260 371628 411312 371680
rect 375104 371560 375156 371612
rect 407120 371560 407172 371612
rect 379520 371492 379572 371544
rect 379888 371492 379940 371544
rect 412640 371492 412692 371544
rect 44732 371356 44784 371408
rect 47584 371356 47636 371408
rect 80060 371356 80112 371408
rect 210884 371356 210936 371408
rect 238116 371356 238168 371408
rect 373172 371424 373224 371476
rect 373724 371424 373776 371476
rect 376760 371424 376812 371476
rect 378048 371424 378100 371476
rect 411260 371424 411312 371476
rect 240048 371356 240100 371408
rect 371056 371356 371108 371408
rect 379980 371356 380032 371408
rect 380992 371356 381044 371408
rect 422300 371356 422352 371408
rect 438216 371356 438268 371408
rect 516600 371356 516652 371408
rect 44824 371288 44876 371340
rect 46112 371288 46164 371340
rect 79508 371288 79560 371340
rect 204168 371288 204220 371340
rect 343180 371288 343232 371340
rect 360292 371288 360344 371340
rect 503168 371288 503220 371340
rect 517888 371288 517940 371340
rect 44916 371220 44968 371272
rect 47860 371220 47912 371272
rect 81440 371220 81492 371272
rect 84568 371220 84620 371272
rect 106188 371220 106240 371272
rect 3516 371152 3568 371204
rect 40684 371152 40736 371204
rect 47676 371152 47728 371204
rect 183284 371152 183336 371204
rect 201592 371220 201644 371272
rect 343456 371220 343508 371272
rect 357440 371220 357492 371272
rect 502340 371220 502392 371272
rect 198832 371152 198884 371204
rect 305000 371152 305052 371204
rect 357900 371152 357952 371204
rect 473360 371152 473412 371204
rect 47768 371084 47820 371136
rect 182732 371084 182784 371136
rect 197544 371084 197596 371136
rect 298100 371084 298152 371136
rect 357348 371084 357400 371136
rect 470600 371084 470652 371136
rect 104624 371016 104676 371068
rect 215484 371016 215536 371068
rect 217416 371016 217468 371068
rect 307760 371016 307812 371068
rect 366272 371016 366324 371068
rect 465080 371016 465132 371068
rect 196716 370948 196768 371000
rect 287244 370948 287296 371000
rect 369032 370948 369084 371000
rect 467840 370948 467892 371000
rect 202420 370880 202472 370932
rect 300860 370880 300912 370932
rect 358728 370880 358780 370932
rect 437480 370880 437532 370932
rect 197452 370812 197504 370864
rect 295340 370812 295392 370864
rect 359648 370812 359700 370864
rect 415400 370812 415452 370864
rect 198280 370744 198332 370796
rect 292580 370744 292632 370796
rect 361396 370744 361448 370796
rect 412824 370744 412876 370796
rect 196808 370676 196860 370728
rect 289820 370676 289872 370728
rect 368296 370676 368348 370728
rect 374552 370676 374604 370728
rect 377128 370676 377180 370728
rect 416780 370676 416832 370728
rect 196624 370608 196676 370660
rect 285680 370608 285732 370660
rect 373080 370608 373132 370660
rect 379612 370608 379664 370660
rect 414020 370608 414072 370660
rect 196992 370540 197044 370592
rect 277400 370540 277452 370592
rect 374552 370540 374604 370592
rect 396080 370540 396132 370592
rect 52920 370472 52972 370524
rect 58624 370472 58676 370524
rect 198740 370472 198792 370524
rect 274640 370472 274692 370524
rect 374460 370472 374512 370524
rect 377128 370472 377180 370524
rect 206836 370404 206888 370456
rect 270500 370404 270552 370456
rect 106188 370336 106240 370388
rect 212448 370336 212500 370388
rect 276020 370336 276072 370388
rect 370412 370336 370464 370388
rect 376668 370336 376720 370388
rect 402980 370472 403032 370524
rect 208032 370268 208084 370320
rect 264980 370268 265032 370320
rect 371792 370268 371844 370320
rect 377496 370268 377548 370320
rect 403256 370336 403308 370388
rect 208584 370200 208636 370252
rect 213552 370200 213604 370252
rect 215484 369860 215536 369912
rect 217232 369860 217284 369912
rect 202880 369792 202932 369844
rect 322940 369792 322992 369844
rect 357992 369792 358044 369844
rect 485780 369792 485832 369844
rect 200672 369724 200724 369776
rect 313280 369724 313332 369776
rect 357256 369724 357308 369776
rect 483020 369724 483072 369776
rect 200212 369656 200264 369708
rect 310520 369656 310572 369708
rect 375748 369656 375800 369708
rect 480260 369656 480312 369708
rect 203524 369588 203576 369640
rect 280160 369588 280212 369640
rect 364892 369588 364944 369640
rect 430580 369588 430632 369640
rect 76840 369520 76892 369572
rect 203064 369520 203116 369572
rect 211528 369520 211580 369572
rect 282920 369520 282972 369572
rect 362776 369520 362828 369572
rect 427820 369520 427872 369572
rect 205364 369452 205416 369504
rect 267740 369452 267792 369504
rect 376484 369452 376536 369504
rect 418160 369452 418212 369504
rect 77208 369384 77260 369436
rect 204260 369384 204312 369436
rect 212908 369384 212960 369436
rect 258172 369384 258224 369436
rect 373724 369384 373776 369436
rect 373908 369384 373960 369436
rect 377220 369384 377272 369436
rect 378692 369384 378744 369436
rect 415676 369384 415728 369436
rect 108856 369316 108908 369368
rect 208124 369316 208176 369368
rect 208860 369316 208912 369368
rect 273260 369316 273312 369368
rect 357164 369316 357216 369368
rect 379336 369316 379388 369368
rect 419540 369316 419592 369368
rect 111616 369248 111668 369300
rect 208952 369248 209004 369300
rect 218428 369248 218480 369300
rect 263600 369248 263652 369300
rect 201040 369180 201092 369232
rect 249800 369180 249852 369232
rect 360660 369180 360712 369232
rect 373080 369180 373132 369232
rect 418252 369248 418304 369300
rect 375840 369180 375892 369232
rect 376484 369180 376536 369232
rect 102048 369112 102100 369164
rect 214104 369112 214156 369164
rect 214472 369112 214524 369164
rect 215852 369112 215904 369164
rect 260840 369112 260892 369164
rect 371148 369112 371200 369164
rect 375932 369112 375984 369164
rect 423680 369180 423732 369232
rect 83832 369044 83884 369096
rect 207204 369044 207256 369096
rect 214380 369044 214432 369096
rect 255320 369044 255372 369096
rect 369584 369044 369636 369096
rect 371792 369044 371844 369096
rect 431960 369112 432012 369164
rect 210240 368976 210292 369028
rect 247040 368976 247092 369028
rect 101680 368908 101732 368960
rect 214012 368908 214064 368960
rect 215300 368908 215352 368960
rect 217508 368908 217560 368960
rect 252652 368908 252704 368960
rect 102784 368840 102836 368892
rect 216404 368840 216456 368892
rect 105636 368772 105688 368824
rect 215576 368772 215628 368824
rect 376576 368432 376628 368484
rect 379704 368432 379756 368484
rect 436100 368432 436152 368484
rect 379796 368228 379848 368280
rect 380072 368228 380124 368280
rect 359004 367956 359056 368008
rect 359556 367956 359608 368008
rect 373172 367956 373224 368008
rect 376484 367956 376536 368008
rect 408500 367956 408552 368008
rect 362684 367888 362736 367940
rect 379428 367888 379480 367940
rect 426440 367888 426492 367940
rect 364156 367820 364208 367872
rect 374460 367820 374512 367872
rect 429200 367820 429252 367872
rect 199384 367752 199436 367804
rect 359004 367752 359056 367804
rect 366916 367752 366968 367804
rect 371148 367752 371200 367804
rect 430672 367752 430724 367804
rect 359924 366324 359976 366376
rect 519360 366324 519412 366376
rect 199844 363604 199896 363656
rect 358912 363604 358964 363656
rect 359832 360816 359884 360868
rect 519084 360816 519136 360868
rect 519636 360816 519688 360868
rect 358912 359524 358964 359576
rect 359648 359524 359700 359576
rect 519176 359524 519228 359576
rect 519360 359524 519412 359576
rect 199568 359456 199620 359508
rect 199752 359456 199804 359508
rect 359096 359456 359148 359508
rect 359924 359456 359976 359508
rect 359188 358708 359240 358760
rect 359464 358708 359516 358760
rect 359464 358028 359516 358080
rect 519268 358028 519320 358080
rect 359556 356736 359608 356788
rect 518992 356736 519044 356788
rect 519544 356736 519596 356788
rect 199660 356668 199712 356720
rect 359004 356668 359056 356720
rect 359832 356668 359884 356720
rect 179328 351908 179380 351960
rect 201500 351908 201552 351960
rect 203064 351908 203116 351960
rect 206284 351908 206336 351960
rect 338488 351296 338540 351348
rect 357072 351296 357124 351348
rect 340512 351228 340564 351280
rect 361580 351296 361632 351348
rect 500592 351296 500644 351348
rect 517704 351296 517756 351348
rect 360200 351228 360252 351280
rect 360844 351228 360896 351280
rect 499028 351228 499080 351280
rect 517796 351228 517848 351280
rect 191288 351160 191340 351212
rect 202880 351160 202932 351212
rect 203064 351160 203116 351212
rect 351644 351160 351696 351212
rect 179696 350548 179748 350600
rect 196624 350548 196676 350600
rect 510896 350548 510948 350600
rect 511908 350548 511960 350600
rect 517520 350548 517572 350600
rect 219348 350480 219400 350532
rect 220820 350480 220872 350532
rect 277308 349800 277360 349852
rect 357532 349800 357584 349852
rect 502248 349800 502300 349852
rect 517612 349800 517664 349852
rect 378600 349528 378652 349580
rect 380900 349528 380952 349580
rect 216772 349188 216824 349240
rect 220912 349188 220964 349240
rect 58624 349052 58676 349104
rect 60740 349052 60792 349104
rect 58900 348644 58952 348696
rect 62120 348644 62172 348696
rect 57152 346876 57204 346928
rect 59360 346876 59412 346928
rect 540244 339396 540296 339448
rect 580172 339396 580224 339448
rect 52920 320084 52972 320136
rect 54300 320084 54352 320136
rect 48044 292476 48096 292528
rect 57060 292476 57112 292528
rect 57336 292476 57388 292528
rect 57152 292204 57204 292256
rect 59728 292204 59780 292256
rect 56876 291864 56928 291916
rect 57980 291864 58032 291916
rect 376944 276224 376996 276276
rect 376944 276020 376996 276072
rect 46296 275952 46348 276004
rect 57612 275952 57664 276004
rect 203800 275952 203852 276004
rect 216680 275952 216732 276004
rect 358084 275952 358136 276004
rect 376852 275952 376904 276004
rect 202880 274592 202932 274644
rect 216680 274592 216732 274644
rect 360200 274592 360252 274644
rect 376760 274592 376812 274644
rect 198004 273912 198056 273964
rect 202880 273912 202932 273964
rect 358084 273232 358136 273284
rect 360200 273232 360252 273284
rect 206744 273164 206796 273216
rect 216680 273164 216732 273216
rect 363972 273164 364024 273216
rect 376760 273164 376812 273216
rect 376852 272484 376904 272536
rect 377036 272484 377088 272536
rect 54300 271124 54352 271176
rect 57980 271124 58032 271176
rect 214380 265344 214432 265396
rect 215024 265344 215076 265396
rect 214656 265208 214708 265260
rect 215024 265208 215076 265260
rect 48872 264936 48924 264988
rect 58624 264936 58676 264988
rect 51540 264868 51592 264920
rect 110972 264868 111024 264920
rect 219164 264868 219216 264920
rect 221188 264868 221240 264920
rect 373632 264868 373684 264920
rect 425980 264868 426032 264920
rect 42156 264800 42208 264852
rect 125968 264800 126020 264852
rect 218612 264800 218664 264852
rect 221096 264800 221148 264852
rect 368204 264800 368256 264852
rect 421104 264800 421156 264852
rect 45008 264732 45060 264784
rect 130936 264732 130988 264784
rect 208032 264732 208084 264784
rect 214656 264732 214708 264784
rect 218520 264732 218572 264784
rect 221004 264732 221056 264784
rect 373080 264732 373132 264784
rect 374460 264732 374512 264784
rect 429752 264732 429804 264784
rect 43536 264664 43588 264716
rect 128360 264664 128412 264716
rect 207848 264664 207900 264716
rect 250444 264664 250496 264716
rect 362592 264664 362644 264716
rect 418436 264664 418488 264716
rect 45192 264596 45244 264648
rect 133420 264596 133472 264648
rect 217232 264596 217284 264648
rect 220912 264596 220964 264648
rect 224224 264596 224276 264648
rect 274180 264596 274232 264648
rect 365536 264596 365588 264648
rect 468484 264596 468536 264648
rect 45100 264528 45152 264580
rect 135904 264528 135956 264580
rect 214840 264528 214892 264580
rect 280804 264528 280856 264580
rect 375012 264528 375064 264580
rect 480904 264528 480956 264580
rect 46204 264460 46256 264512
rect 138480 264460 138532 264512
rect 216220 264460 216272 264512
rect 285956 264460 286008 264512
rect 366824 264460 366876 264512
rect 473452 264460 473504 264512
rect 48136 264392 48188 264444
rect 143540 264392 143592 264444
rect 210792 264392 210844 264444
rect 283380 264392 283432 264444
rect 363880 264392 363932 264444
rect 470968 264392 471020 264444
rect 43444 264324 43496 264376
rect 140872 264324 140924 264376
rect 209412 264324 209464 264376
rect 290924 264324 290976 264376
rect 372344 264324 372396 264376
rect 483388 264324 483440 264376
rect 45284 264256 45336 264308
rect 145932 264256 145984 264308
rect 203708 264256 203760 264308
rect 288164 264256 288216 264308
rect 369492 264256 369544 264308
rect 485964 264256 486016 264308
rect 45376 264188 45428 264240
rect 148508 264188 148560 264240
rect 200948 264188 201000 264240
rect 293408 264188 293460 264240
rect 356888 264188 356940 264240
rect 475844 264188 475896 264240
rect 46388 264120 46440 264172
rect 62212 264120 62264 264172
rect 213000 264120 213052 264172
rect 224224 264120 224276 264172
rect 370964 264120 371016 264172
rect 423496 264120 423548 264172
rect 46480 264052 46532 264104
rect 62120 264052 62172 264104
rect 214656 264052 214708 264104
rect 220820 264052 220872 264104
rect 62212 263712 62264 263764
rect 89996 263712 90048 263764
rect 58900 263644 58952 263696
rect 62304 263644 62356 263696
rect 92388 263644 92440 263696
rect 211620 263644 211672 263696
rect 214288 263644 214340 263696
rect 62120 263576 62172 263628
rect 91284 263576 91336 263628
rect 212356 263576 212408 263628
rect 213000 263576 213052 263628
rect 373908 263644 373960 263696
rect 374368 263644 374420 263696
rect 433340 263644 433392 263696
rect 273260 263576 273312 263628
rect 279240 263576 279292 263628
rect 357716 263576 357768 263628
rect 359280 263576 359332 263628
rect 371792 263576 371844 263628
rect 373632 263576 373684 263628
rect 432236 263576 432288 263628
rect 54484 263508 54536 263560
rect 120908 263508 120960 263560
rect 155960 263508 156012 263560
rect 204352 263508 204404 263560
rect 210700 263508 210752 263560
rect 308404 263508 308456 263560
rect 362500 263508 362552 263560
rect 453396 263508 453448 263560
rect 57796 263440 57848 263492
rect 123484 263440 123536 263492
rect 158536 263440 158588 263492
rect 205640 263440 205692 263492
rect 212264 263440 212316 263492
rect 305828 263440 305880 263492
rect 368112 263440 368164 263492
rect 455788 263440 455840 263492
rect 53104 263372 53156 263424
rect 115940 263372 115992 263424
rect 150992 263372 151044 263424
rect 197636 263372 197688 263424
rect 205088 263372 205140 263424
rect 268292 263372 268344 263424
rect 370872 263372 370924 263424
rect 451004 263372 451056 263424
rect 54576 263304 54628 263356
rect 118056 263304 118108 263356
rect 161112 263304 161164 263356
rect 207112 263304 207164 263356
rect 214748 263304 214800 263356
rect 276112 263304 276164 263356
rect 364064 263304 364116 263356
rect 443460 263304 443512 263356
rect 53012 263236 53064 263288
rect 113364 263236 113416 263288
rect 166080 263236 166132 263288
rect 210056 263236 210108 263288
rect 210608 263236 210660 263288
rect 270868 263236 270920 263288
rect 361304 263236 361356 263288
rect 438400 263236 438452 263288
rect 53380 263168 53432 263220
rect 108212 263168 108264 263220
rect 163504 263168 163556 263220
rect 197728 263168 197780 263220
rect 209320 263168 209372 263220
rect 265900 263168 265952 263220
rect 372252 263168 372304 263220
rect 448244 263168 448296 263220
rect 51632 263100 51684 263152
rect 105636 263100 105688 263152
rect 200856 263100 200908 263152
rect 256148 263100 256200 263152
rect 365352 263100 365404 263152
rect 435916 263100 435968 263152
rect 51816 263032 51868 263084
rect 103520 263032 103572 263084
rect 206560 263032 206612 263084
rect 260932 263032 260984 263084
rect 373540 263032 373592 263084
rect 440884 263032 440936 263084
rect 503536 263032 503588 263084
rect 517612 263032 517664 263084
rect 50252 262964 50304 263016
rect 101036 262964 101088 263016
rect 183376 262964 183428 263016
rect 201592 262964 201644 263016
rect 218980 262964 219032 263016
rect 273352 262964 273404 263016
rect 343548 262964 343600 263016
rect 357440 262964 357492 263016
rect 369308 262964 369360 263016
rect 433524 262964 433576 263016
rect 50344 262896 50396 262948
rect 98092 262896 98144 262948
rect 183468 262896 183520 262948
rect 202972 262896 203024 262948
rect 212172 262896 212224 262948
rect 263600 262896 263652 262948
rect 369400 262896 369452 262948
rect 410708 262896 410760 262948
rect 503628 262896 503680 262948
rect 517888 262896 517940 262948
rect 50436 262828 50488 262880
rect 96068 262828 96120 262880
rect 114376 262828 114428 262880
rect 196900 262828 196952 262880
rect 202236 262828 202288 262880
rect 253572 262828 253624 262880
rect 343456 262828 343508 262880
rect 360292 262828 360344 262880
rect 374828 262828 374880 262880
rect 413652 262828 413704 262880
rect 49148 262760 49200 262812
rect 93584 262760 93636 262812
rect 207940 262760 207992 262812
rect 258356 262760 258408 262812
rect 379060 262760 379112 262812
rect 415768 262760 415820 262812
rect 55772 262692 55824 262744
rect 90732 262692 90784 262744
rect 215024 262692 215076 262744
rect 247684 262692 247736 262744
rect 374920 262692 374972 262744
rect 408316 262692 408368 262744
rect 54668 262624 54720 262676
rect 88340 262624 88392 262676
rect 96528 262624 96580 262676
rect 101772 262624 101824 262676
rect 210332 262624 210384 262676
rect 213276 262624 213328 262676
rect 100024 262420 100076 262472
rect 116216 262420 116268 262472
rect 511908 262420 511960 262472
rect 517520 262420 517572 262472
rect 89720 262352 89772 262404
rect 109316 262352 109368 262404
rect 213276 262216 213328 262268
rect 272064 262216 272116 262268
rect 378692 262216 378744 262268
rect 379980 262216 380032 262268
rect 415860 262216 415912 262268
rect 425704 262216 425756 262268
rect 428280 262216 428332 262268
rect 206652 262148 206704 262200
rect 325792 262148 325844 262200
rect 365444 262148 365496 262200
rect 430948 262148 431000 262200
rect 205180 262080 205232 262132
rect 323032 262080 323084 262132
rect 374920 262080 374972 262132
rect 375840 262080 375892 262132
rect 376300 262080 376352 262132
rect 428188 262080 428240 262132
rect 211712 262012 211764 262064
rect 212908 262012 212960 262064
rect 373172 262012 373224 262064
rect 376392 262012 376444 262064
rect 378600 262012 378652 262064
rect 379244 262012 379296 262064
rect 426440 262012 426492 262064
rect 372988 261944 373040 261996
rect 376300 261944 376352 261996
rect 379612 261944 379664 261996
rect 396172 261944 396224 261996
rect 212908 261536 212960 261588
rect 269764 261536 269816 261588
rect 375840 261536 375892 261588
rect 393412 261536 393464 261588
rect 208952 261468 209004 261520
rect 212816 261468 212868 261520
rect 271236 261468 271288 261520
rect 380348 261468 380400 261520
rect 425244 261468 425296 261520
rect 379336 260992 379388 261044
rect 389180 260992 389232 261044
rect 376300 260924 376352 260976
rect 388444 260924 388496 260976
rect 52828 260856 52880 260908
rect 57980 260856 58032 260908
rect 59728 260788 59780 260840
rect 118700 260788 118752 260840
rect 213552 260788 213604 260840
rect 214380 260788 214432 260840
rect 214840 260788 214892 260840
rect 376392 260856 376444 260908
rect 390560 260856 390612 260908
rect 244372 260788 244424 260840
rect 375012 260788 375064 260840
rect 375196 260788 375248 260840
rect 375932 260788 375984 260840
rect 377036 260788 377088 260840
rect 100760 260720 100812 260772
rect 213092 260720 213144 260772
rect 214748 260720 214800 260772
rect 243084 260720 243136 260772
rect 435180 260788 435232 260840
rect 388444 260720 388496 260772
rect 421748 260720 421800 260772
rect 50528 260652 50580 260704
rect 84200 260652 84252 260704
rect 389180 260652 389232 260704
rect 419816 260652 419868 260704
rect 51724 260584 51776 260636
rect 84752 260584 84804 260636
rect 390560 260584 390612 260636
rect 419356 260584 419408 260636
rect 53196 260516 53248 260568
rect 54576 260516 54628 260568
rect 87604 260516 87656 260568
rect 393412 260516 393464 260568
rect 418160 260516 418212 260568
rect 55772 260448 55824 260500
rect 88616 260448 88668 260500
rect 49056 260380 49108 260432
rect 89720 260380 89772 260432
rect 57980 260312 58032 260364
rect 102324 260312 102376 260364
rect 52920 260244 52972 260296
rect 54300 260244 54352 260296
rect 99472 260244 99524 260296
rect 45468 260176 45520 260228
rect 49056 260176 49108 260228
rect 51632 260176 51684 260228
rect 105084 260176 105136 260228
rect 377036 260176 377088 260228
rect 423956 260176 424008 260228
rect 42248 260108 42300 260160
rect 46204 260108 46256 260160
rect 108028 260108 108080 260160
rect 214748 260108 214800 260160
rect 236000 260108 236052 260160
rect 379612 260108 379664 260160
rect 427452 260108 427504 260160
rect 53288 260040 53340 260092
rect 85948 260040 86000 260092
rect 54392 259972 54444 260024
rect 64880 259972 64932 260024
rect 43720 259360 43772 259412
rect 57980 259360 58032 259412
rect 46664 259292 46716 259344
rect 55772 259292 55824 259344
rect 43628 259224 43680 259276
rect 51632 259224 51684 259276
rect 372436 244196 372488 244248
rect 374552 244196 374604 244248
rect 440148 244196 440200 244248
rect 516692 244196 516744 244248
rect 371056 243652 371108 243704
rect 373540 243652 373592 243704
rect 398840 243652 398892 243704
rect 374552 243584 374604 243636
rect 374828 243584 374880 243636
rect 401600 243584 401652 243636
rect 368388 243516 368440 243568
rect 373448 243516 373500 243568
rect 400220 243516 400272 243568
rect 356888 242632 356940 242684
rect 361580 242632 361632 242684
rect 196716 242088 196768 242140
rect 201500 242088 201552 242140
rect 54392 241544 54444 241596
rect 64880 241544 64932 241596
rect 53012 241476 53064 241528
rect 66076 241476 66128 241528
rect 46112 241408 46164 241460
rect 46296 241408 46348 241460
rect 47860 241408 47912 241460
rect 48044 241408 48096 241460
rect 357256 241476 357308 241528
rect 360200 241476 360252 241528
rect 47492 241340 47544 241392
rect 48136 241340 48188 241392
rect 99380 241408 99432 241460
rect 210976 241408 211028 241460
rect 214288 241408 214340 241460
rect 214656 241408 214708 241460
rect 216772 241408 216824 241460
rect 240140 241408 240192 241460
rect 275928 241408 275980 241460
rect 356612 241408 356664 241460
rect 374460 241408 374512 241460
rect 375196 241408 375248 241460
rect 375748 241408 375800 241460
rect 376484 241408 376536 241460
rect 81440 241340 81492 241392
rect 219532 241340 219584 241392
rect 221188 241340 221240 241392
rect 253940 241340 253992 241392
rect 277308 241340 277360 241392
rect 356980 241340 357032 241392
rect 46296 241272 46348 241324
rect 78680 241272 78732 241324
rect 213000 241272 213052 241324
rect 214932 241272 214984 241324
rect 247132 241272 247184 241324
rect 278688 241272 278740 241324
rect 357532 241272 357584 241324
rect 376484 241272 376536 241324
rect 377496 241272 377548 241324
rect 378600 241408 378652 241460
rect 379888 241408 379940 241460
rect 412732 241408 412784 241460
rect 438768 241408 438820 241460
rect 516600 241408 516652 241460
rect 378048 241340 378100 241392
rect 378692 241340 378744 241392
rect 408500 241340 408552 241392
rect 379428 241272 379480 241324
rect 407212 241272 407264 241324
rect 47584 241204 47636 241256
rect 80060 241204 80112 241256
rect 219624 241204 219676 241256
rect 220268 241204 220320 241256
rect 251180 241204 251232 241256
rect 339408 241204 339460 241256
rect 357256 241204 357308 241256
rect 377588 241204 377640 241256
rect 379796 241204 379848 241256
rect 411260 241204 411312 241256
rect 48136 241136 48188 241188
rect 77300 241136 77352 241188
rect 219900 241136 219952 241188
rect 220636 241136 220688 241188
rect 251272 241136 251324 241188
rect 373816 241136 373868 241188
rect 404360 241136 404412 241188
rect 66260 241068 66312 241120
rect 96620 241068 96672 241120
rect 219808 241068 219860 241120
rect 220084 241068 220136 241120
rect 249800 241068 249852 241120
rect 377680 241068 377732 241120
rect 379704 241068 379756 241120
rect 409880 241068 409932 241120
rect 180156 241000 180208 241052
rect 196624 241000 196676 241052
rect 220728 241000 220780 241052
rect 248420 241000 248472 241052
rect 376668 241000 376720 241052
rect 402980 241000 403032 241052
rect 183376 240932 183428 240984
rect 200120 240932 200172 240984
rect 210884 240932 210936 240984
rect 237380 240932 237432 240984
rect 377496 240932 377548 240984
rect 403072 240932 403124 240984
rect 503628 240932 503680 240984
rect 517888 240932 517940 240984
rect 179328 240864 179380 240916
rect 196716 240864 196768 240916
rect 213368 240864 213420 240916
rect 218980 240864 219032 240916
rect 245660 240864 245712 240916
rect 343456 240864 343508 240916
rect 359464 240864 359516 240916
rect 372528 240864 372580 240916
rect 379060 240864 379112 240916
rect 405740 240864 405792 240916
rect 500776 240864 500828 240916
rect 517704 240864 517756 240916
rect 183468 240796 183520 240848
rect 201500 240796 201552 240848
rect 214288 240796 214340 240848
rect 244280 240796 244332 240848
rect 340052 240796 340104 240848
rect 356888 240796 356940 240848
rect 375104 240796 375156 240848
rect 67548 240728 67600 240780
rect 98000 240728 98052 240780
rect 209504 240728 209556 240780
rect 210792 240728 210844 240780
rect 241520 240728 241572 240780
rect 351552 240728 351604 240780
rect 358084 240728 358136 240780
rect 375656 240728 375708 240780
rect 376668 240728 376720 240780
rect 378692 240796 378744 240848
rect 411352 240796 411404 240848
rect 499028 240796 499080 240848
rect 517796 240796 517848 240848
rect 379428 240728 379480 240780
rect 379888 240728 379940 240780
rect 414020 240728 414072 240780
rect 218336 240660 218388 240712
rect 219348 240660 219400 240712
rect 252652 240660 252704 240712
rect 369676 240660 369728 240712
rect 372528 240660 372580 240712
rect 397460 240660 397512 240712
rect 213552 240524 213604 240576
rect 216312 240524 216364 240576
rect 238760 240592 238812 240644
rect 374552 240592 374604 240644
rect 396172 240592 396224 240644
rect 511908 240592 511960 240644
rect 517520 240592 517572 240644
rect 375196 240456 375248 240508
rect 396080 240456 396132 240508
rect 216312 240388 216364 240440
rect 219716 240388 219768 240440
rect 220728 240388 220780 240440
rect 217600 240252 217652 240304
rect 220268 240252 220320 240304
rect 190920 240184 190972 240236
rect 198004 240184 198056 240236
rect 219348 240184 219400 240236
rect 220636 240184 220688 240236
rect 50620 240048 50672 240100
rect 53104 240048 53156 240100
rect 58992 240048 59044 240100
rect 62304 240048 62356 240100
rect 214932 240048 214984 240100
rect 215300 240048 215352 240100
rect 219900 240048 219952 240100
rect 221096 240048 221148 240100
rect 222108 240048 222160 240100
rect 267740 240048 267792 240100
rect 371148 240048 371200 240100
rect 373172 240048 373224 240100
rect 376576 240048 376628 240100
rect 436100 240048 436152 240100
rect 58808 239980 58860 240032
rect 62212 239980 62264 240032
rect 213644 239980 213696 240032
rect 215668 239980 215720 240032
rect 218612 239980 218664 240032
rect 219256 239980 219308 240032
rect 264980 239980 265032 240032
rect 375288 239980 375340 240032
rect 434720 239980 434772 240032
rect 55680 239912 55732 239964
rect 60740 239912 60792 239964
rect 216404 239912 216456 239964
rect 262220 239912 262272 239964
rect 378048 239912 378100 239964
rect 423680 239912 423732 239964
rect 219808 239844 219860 239896
rect 220820 239844 220872 239896
rect 221096 239844 221148 239896
rect 266452 239844 266504 239896
rect 369768 239844 369820 239896
rect 379704 239844 379756 239896
rect 425704 239844 425756 239896
rect 53104 239776 53156 239828
rect 67548 239776 67600 239828
rect 217232 239776 217284 239828
rect 217968 239776 218020 239828
rect 219164 239776 219216 239828
rect 220728 239776 220780 239828
rect 222108 239776 222160 239828
rect 222200 239776 222252 239828
rect 266360 239776 266412 239828
rect 57152 239708 57204 239760
rect 82084 239708 82136 239760
rect 215300 239708 215352 239760
rect 259552 239708 259604 239760
rect 53840 239640 53892 239692
rect 100024 239640 100076 239692
rect 219624 239640 219676 239692
rect 220912 239640 220964 239692
rect 263600 239640 263652 239692
rect 60648 239572 60700 239624
rect 107660 239572 107712 239624
rect 217048 239572 217100 239624
rect 219072 239572 219124 239624
rect 258172 239572 258224 239624
rect 58900 239504 58952 239556
rect 107752 239504 107804 239556
rect 215668 239504 215720 239556
rect 256700 239504 256752 239556
rect 50804 239436 50856 239488
rect 110420 239436 110472 239488
rect 218520 239436 218572 239488
rect 259460 239436 259512 239488
rect 51816 239368 51868 239420
rect 113180 239368 113232 239420
rect 216220 239368 216272 239420
rect 260840 239368 260892 239420
rect 373172 239368 373224 239420
rect 430672 239368 430724 239420
rect 217968 239300 218020 239352
rect 255320 239300 255372 239352
rect 57244 239232 57296 239284
rect 62120 239232 62172 239284
rect 220820 239232 220872 239284
rect 222108 239232 222160 239284
rect 375932 239232 375984 239284
rect 376576 239232 376628 239284
rect 372436 238756 372488 238808
rect 375288 238756 375340 238808
rect 46848 238688 46900 238740
rect 50804 238688 50856 238740
rect 214472 238688 214524 238740
rect 216220 238688 216272 238740
rect 42340 238620 42392 238672
rect 46756 238620 46808 238672
rect 51816 238620 51868 238672
rect 215208 238620 215260 238672
rect 218520 238620 218572 238672
rect 47952 238552 48004 238604
rect 60648 238552 60700 238604
rect 53840 238484 53892 238536
rect 43812 238416 43864 238468
rect 57152 238416 57204 238468
rect 50344 237396 50396 237448
rect 50804 237396 50856 237448
rect 51540 237396 51592 237448
rect 51816 237396 51868 237448
rect 53840 237396 53892 237448
rect 54484 237396 54536 237448
rect 56968 235968 57020 236020
rect 59728 235968 59780 236020
rect 2872 169668 2924 169720
rect 4804 169668 4856 169720
rect 207756 165520 207808 165572
rect 216680 165520 216732 165572
rect 362408 165520 362460 165572
rect 376944 165520 376996 165572
rect 377772 165112 377824 165164
rect 377956 165112 378008 165164
rect 203616 164160 203668 164212
rect 217048 164160 217100 164212
rect 367836 164160 367888 164212
rect 376760 164160 376812 164212
rect 198004 163480 198056 163532
rect 216680 163480 216732 163532
rect 358084 163480 358136 163532
rect 376944 163480 376996 163532
rect 377772 156612 377824 156664
rect 377956 156612 378008 156664
rect 42432 154640 42484 154692
rect 163320 154640 163372 154692
rect 43904 154572 43956 154624
rect 165896 154572 165948 154624
rect 50344 154504 50396 154556
rect 51816 154504 51868 154556
rect 56968 154504 57020 154556
rect 59360 154504 59412 154556
rect 358268 154504 358320 154556
rect 418436 154504 418488 154556
rect 50712 154436 50764 154488
rect 96068 154436 96120 154488
rect 358360 154436 358412 154488
rect 421012 154436 421064 154488
rect 49516 154368 49568 154420
rect 98460 154368 98512 154420
rect 357624 154368 357676 154420
rect 360292 154368 360344 154420
rect 362316 154368 362368 154420
rect 425980 154368 426032 154420
rect 438860 154368 438912 154420
rect 516600 154368 516652 154420
rect 52092 154300 52144 154352
rect 101036 154300 101088 154352
rect 365260 154300 365312 154352
rect 443460 154300 443512 154352
rect 53564 154232 53616 154284
rect 105820 154232 105872 154284
rect 206468 154232 206520 154284
rect 261024 154232 261076 154284
rect 372160 154232 372212 154284
rect 475844 154232 475896 154284
rect 56324 154164 56376 154216
rect 138388 154164 138440 154216
rect 202144 154164 202196 154216
rect 273536 154164 273588 154216
rect 373356 154164 373408 154216
rect 478420 154164 478472 154216
rect 52184 154096 52236 154148
rect 108212 154096 108264 154148
rect 113364 154096 113416 154148
rect 114468 154096 114520 154148
rect 196808 154096 196860 154148
rect 204996 154096 205048 154148
rect 293316 154096 293368 154148
rect 366640 154096 366692 154148
rect 473452 154096 473504 154148
rect 59268 154028 59320 154080
rect 143540 154028 143592 154080
rect 198096 154028 198148 154080
rect 288164 154028 288216 154080
rect 369216 154028 369268 154080
rect 480812 154028 480864 154080
rect 46388 153960 46440 154012
rect 52184 153960 52236 154012
rect 59912 153960 59964 154012
rect 145932 153960 145984 154012
rect 206376 153960 206428 154012
rect 298468 153960 298520 154012
rect 356796 153960 356848 154012
rect 470876 153960 470928 154012
rect 510528 153960 510580 154012
rect 517520 153960 517572 154012
rect 60004 153892 60056 153944
rect 150900 153892 150952 153944
rect 210516 153892 210568 153944
rect 303436 153892 303488 153944
rect 368020 153892 368072 153944
rect 483204 153892 483256 153944
rect 59176 153824 59228 153876
rect 153292 153824 153344 153876
rect 209228 153824 209280 153876
rect 308404 153824 308456 153876
rect 370780 153824 370832 153876
rect 485964 153824 486016 153876
rect 366548 153756 366600 153808
rect 423404 153756 423456 153808
rect 51816 153348 51868 153400
rect 111156 153348 111208 153400
rect 59360 153280 59412 153332
rect 118700 153280 118752 153332
rect 52184 153212 52236 153264
rect 114744 153212 114796 153264
rect 197360 153212 197412 153264
rect 201500 153212 201552 153264
rect 373632 153212 373684 153264
rect 373816 153212 373868 153264
rect 431960 153212 432012 153264
rect 51908 153144 51960 153196
rect 155960 153144 156012 153196
rect 210424 153144 210476 153196
rect 300860 153144 300912 153196
rect 361120 153144 361172 153196
rect 455420 153144 455472 153196
rect 56140 153076 56192 153128
rect 135260 153076 135312 153128
rect 209044 153076 209096 153128
rect 285680 153076 285732 153128
rect 358452 153076 358504 153128
rect 447140 153076 447192 153128
rect 55956 153008 56008 153060
rect 132776 153008 132828 153060
rect 215944 153008 215996 153060
rect 289820 153008 289872 153060
rect 376116 153008 376168 153060
rect 458180 153008 458232 153060
rect 54852 152940 54904 152992
rect 129740 152940 129792 152992
rect 211988 152940 212040 152992
rect 277952 152940 278004 152992
rect 373264 152940 373316 152992
rect 452660 152940 452712 152992
rect 56416 152872 56468 152924
rect 128360 152872 128412 152924
rect 216128 152872 216180 152924
rect 280252 152872 280304 152924
rect 369124 152872 369176 152924
rect 445760 152872 445812 152924
rect 54760 152804 54812 152856
rect 125600 152804 125652 152856
rect 218888 152804 218940 152856
rect 282920 152804 282972 152856
rect 363788 152804 363840 152856
rect 440332 152804 440384 152856
rect 56048 152736 56100 152788
rect 122840 152736 122892 152788
rect 209136 152736 209188 152788
rect 268016 152736 268068 152788
rect 374644 152736 374696 152788
rect 449900 152736 449952 152788
rect 54944 152668 54996 152720
rect 120080 152668 120132 152720
rect 200764 152668 200816 152720
rect 255964 152668 256016 152720
rect 365168 152668 365220 152720
rect 434812 152668 434864 152720
rect 53472 152600 53524 152652
rect 117504 152600 117556 152652
rect 183468 152600 183520 152652
rect 197360 152600 197412 152652
rect 216036 152600 216088 152652
rect 265072 152600 265124 152652
rect 343548 152600 343600 152652
rect 357624 152600 357676 152652
rect 371976 152600 372028 152652
rect 437480 152600 437532 152652
rect 503628 152600 503680 152652
rect 517612 152600 517664 152652
rect 52000 152532 52052 152584
rect 113180 152532 113232 152584
rect 204904 152532 204956 152584
rect 253572 152532 253624 152584
rect 370688 152532 370740 152584
rect 433340 152532 433392 152584
rect 55864 152464 55916 152516
rect 115940 152464 115992 152516
rect 183468 152464 183520 152516
rect 200120 152464 200172 152516
rect 213184 152464 213236 152516
rect 258264 152464 258316 152516
rect 343548 152464 343600 152516
rect 359464 152464 359516 152516
rect 376208 152464 376260 152516
rect 415676 152464 415728 152516
rect 503628 152464 503680 152516
rect 517888 152464 517940 152516
rect 50896 152396 50948 152448
rect 103520 152396 103572 152448
rect 214564 152396 214616 152448
rect 250260 152396 250312 152448
rect 374736 152396 374788 152448
rect 413100 152396 413152 152448
rect 49240 152328 49292 152380
rect 89720 152328 89772 152380
rect 97264 152328 97316 152380
rect 100760 152328 100812 152380
rect 218796 152328 218848 152380
rect 247132 152328 247184 152380
rect 372068 152328 372120 152380
rect 409880 152328 409932 152380
rect 55036 152260 55088 152312
rect 88340 152260 88392 152312
rect 378876 152260 378928 152312
rect 407120 152260 407172 152312
rect 98644 151852 98696 151904
rect 104900 151852 104952 151904
rect 212264 151784 212316 151836
rect 219440 151784 219492 151836
rect 55680 151716 55732 151768
rect 57796 151716 57848 151768
rect 117412 151716 117464 151768
rect 212080 151716 212132 151768
rect 320180 151716 320232 151768
rect 375932 151716 375984 151768
rect 436192 151716 436244 151768
rect 53656 151648 53708 151700
rect 110420 151648 110472 151700
rect 219440 151648 219492 151700
rect 219808 151648 219860 151700
rect 267740 151648 267792 151700
rect 277400 151648 277452 151700
rect 278044 151648 278096 151700
rect 356980 151648 357032 151700
rect 379244 151648 379296 151700
rect 426532 151648 426584 151700
rect 54392 151580 54444 151632
rect 54944 151580 54996 151632
rect 98000 151580 98052 151632
rect 219900 151580 219952 151632
rect 266360 151580 266412 151632
rect 375840 151580 375892 151632
rect 218612 151512 218664 151564
rect 219256 151512 219308 151564
rect 264980 151512 265032 151564
rect 376392 151512 376444 151564
rect 380072 151512 380124 151564
rect 380808 151580 380860 151632
rect 427820 151580 427872 151632
rect 422300 151512 422352 151564
rect 216404 151444 216456 151496
rect 262220 151444 262272 151496
rect 53104 151376 53156 151428
rect 57060 151376 57112 151428
rect 96620 151376 96672 151428
rect 214932 151376 214984 151428
rect 259460 151376 259512 151428
rect 425060 151444 425112 151496
rect 60004 151308 60056 151360
rect 106372 151308 106424 151360
rect 216220 151308 216272 151360
rect 261208 151308 261260 151360
rect 379520 151308 379572 151360
rect 379796 151308 379848 151360
rect 52828 151240 52880 151292
rect 54852 151240 54904 151292
rect 100852 151240 100904 151292
rect 219624 151240 219676 151292
rect 263600 151240 263652 151292
rect 376300 151240 376352 151292
rect 420920 151376 420972 151428
rect 380164 151308 380216 151360
rect 418252 151308 418304 151360
rect 380072 151240 380124 151292
rect 418160 151240 418212 151292
rect 59268 151172 59320 151224
rect 106280 151172 106332 151224
rect 217140 151172 217192 151224
rect 258080 151172 258132 151224
rect 379704 151172 379756 151224
rect 423680 151172 423732 151224
rect 49056 151104 49108 151156
rect 55036 151104 55088 151156
rect 109132 151104 109184 151156
rect 219164 151104 219216 151156
rect 219808 151104 219860 151156
rect 266452 151104 266504 151156
rect 373172 151104 373224 151156
rect 375288 151104 375340 151156
rect 430580 151104 430632 151156
rect 46480 151036 46532 151088
rect 51908 151036 51960 151088
rect 111800 151036 111852 151088
rect 213276 151036 213328 151088
rect 216496 151036 216548 151088
rect 271880 151036 271932 151088
rect 372436 151036 372488 151088
rect 374460 151036 374512 151088
rect 433984 151036 434036 151088
rect 218520 150968 218572 151020
rect 218888 150968 218940 151020
rect 259552 150968 259604 151020
rect 379336 150968 379388 151020
rect 419540 150968 419592 151020
rect 374552 150900 374604 150952
rect 396080 150900 396132 150952
rect 375196 150832 375248 150884
rect 396172 150832 396224 150884
rect 374920 150764 374972 150816
rect 380164 150764 380216 150816
rect 58624 150628 58676 150680
rect 60004 150628 60056 150680
rect 375932 150492 375984 150544
rect 376668 150492 376720 150544
rect 377036 150492 377088 150544
rect 379704 150492 379756 150544
rect 214196 150424 214248 150476
rect 214932 150424 214984 150476
rect 216128 150424 216180 150476
rect 216404 150424 216456 150476
rect 376208 150424 376260 150476
rect 376392 150424 376444 150476
rect 379244 150424 379296 150476
rect 379428 150424 379480 150476
rect 47952 150356 48004 150408
rect 58624 150356 58676 150408
rect 59268 150356 59320 150408
rect 214748 150356 214800 150408
rect 236092 150356 236144 150408
rect 212816 149676 212868 149728
rect 214932 149676 214984 149728
rect 270500 149676 270552 149728
rect 52184 147024 52236 147076
rect 52092 146820 52144 146872
rect 51816 146752 51868 146804
rect 52184 146752 52236 146804
rect 54484 133832 54536 133884
rect 117320 133832 117372 133884
rect 212356 133832 212408 133884
rect 213368 133832 213420 133884
rect 213552 133832 213604 133884
rect 273260 133832 273312 133884
rect 378600 133832 378652 133884
rect 379152 133832 379204 133884
rect 48044 133764 48096 133816
rect 53656 133764 53708 133816
rect 56324 133764 56376 133816
rect 56968 133764 57020 133816
rect 103612 133764 103664 133816
rect 47768 133696 47820 133748
rect 53472 133696 53524 133748
rect 214656 133764 214708 133816
rect 240140 133764 240192 133816
rect 375012 133764 375064 133816
rect 436100 133832 436152 133884
rect 379336 133764 379388 133816
rect 434720 133764 434772 133816
rect 46296 133628 46348 133680
rect 54484 133492 54536 133544
rect 54760 133492 54812 133544
rect 238760 133696 238812 133748
rect 379152 133696 379204 133748
rect 412732 133696 412784 133748
rect 210792 133628 210844 133680
rect 215024 133628 215076 133680
rect 374828 133628 374880 133680
rect 401600 133628 401652 133680
rect 372436 133560 372488 133612
rect 373448 133560 373500 133612
rect 400220 133560 400272 133612
rect 80060 133492 80112 133544
rect 377680 133492 377732 133544
rect 379336 133492 379388 133544
rect 51908 133424 51960 133476
rect 78680 133424 78732 133476
rect 213644 133424 213696 133476
rect 214656 133424 214708 133476
rect 53656 133356 53708 133408
rect 81440 133356 81492 133408
rect 46204 133288 46256 133340
rect 59912 133288 59964 133340
rect 109040 133288 109092 133340
rect 51540 133220 51592 133272
rect 53564 133220 53616 133272
rect 114560 133220 114612 133272
rect 215024 133220 215076 133272
rect 241520 133220 241572 133272
rect 53288 133152 53340 133204
rect 114652 133152 114704 133204
rect 216496 133152 216548 133204
rect 278044 133152 278096 133204
rect 280068 133152 280120 133204
rect 306380 133152 306432 133204
rect 373540 133152 373592 133204
rect 375196 133152 375248 133204
rect 398840 133152 398892 133204
rect 373908 132472 373960 132524
rect 374828 132472 374880 132524
rect 306380 131792 306432 131844
rect 356980 131792 357032 131844
rect 356980 131588 357032 131640
rect 357716 131588 357768 131640
rect 191748 131112 191800 131164
rect 198004 131112 198056 131164
rect 213552 131112 213604 131164
rect 274732 131112 274784 131164
rect 55772 131044 55824 131096
rect 56416 131044 56468 131096
rect 56968 131044 57020 131096
rect 57244 131044 57296 131096
rect 59820 131044 59872 131096
rect 93860 131044 93912 131096
rect 179052 131044 179104 131096
rect 196716 131044 196768 131096
rect 216036 131044 216088 131096
rect 218980 131044 219032 131096
rect 245660 131044 245712 131096
rect 338488 131044 338540 131096
rect 360200 131044 360252 131096
rect 379980 131044 380032 131096
rect 415400 131044 415452 131096
rect 91100 130976 91152 131028
rect 179788 130976 179840 131028
rect 196624 130976 196676 131028
rect 219532 130976 219584 131028
rect 253940 130976 253992 131028
rect 340604 130976 340656 131028
rect 356888 130976 356940 131028
rect 377588 130976 377640 131028
rect 411260 130976 411312 131028
rect 500224 130976 500276 131028
rect 517704 130976 517756 131028
rect 56416 130908 56468 130960
rect 88432 130908 88484 130960
rect 218336 130908 218388 130960
rect 218796 130908 218848 130960
rect 252560 130908 252612 130960
rect 379336 130908 379388 130960
rect 411352 130908 411404 130960
rect 498752 130908 498804 130960
rect 517796 130908 517848 130960
rect 51724 130840 51776 130892
rect 84200 130840 84252 130892
rect 217600 130840 217652 130892
rect 251272 130840 251324 130892
rect 377680 130840 377732 130892
rect 409972 130840 410024 130892
rect 53380 130772 53432 130824
rect 85580 130772 85632 130824
rect 218980 130772 219032 130824
rect 219348 130772 219400 130824
rect 251180 130772 251232 130824
rect 376484 130772 376536 130824
rect 48964 130704 49016 130756
rect 55956 130704 56008 130756
rect 59084 130704 59136 130756
rect 91192 130704 91244 130756
rect 216312 130704 216364 130756
rect 248420 130704 248472 130756
rect 380072 130772 380124 130824
rect 408500 130772 408552 130824
rect 402980 130704 403032 130756
rect 58900 130636 58952 130688
rect 59268 130636 59320 130688
rect 89812 130636 89864 130688
rect 214656 130636 214708 130688
rect 244372 130636 244424 130688
rect 379060 130636 379112 130688
rect 405740 130636 405792 130688
rect 55956 130568 56008 130620
rect 82820 130568 82872 130620
rect 214472 130568 214524 130620
rect 242900 130568 242952 130620
rect 378692 130568 378744 130620
rect 379336 130568 379388 130620
rect 380256 130568 380308 130620
rect 403072 130568 403124 130620
rect 54484 130500 54536 130552
rect 84292 130500 84344 130552
rect 213000 130500 213052 130552
rect 219072 130500 219124 130552
rect 247040 130500 247092 130552
rect 375748 130500 375800 130552
rect 380072 130500 380124 130552
rect 380164 130500 380216 130552
rect 407212 130500 407264 130552
rect 55864 130432 55916 130484
rect 86960 130432 87012 130484
rect 183468 130432 183520 130484
rect 197452 130432 197504 130484
rect 214288 130432 214340 130484
rect 214656 130432 214708 130484
rect 215944 130432 215996 130484
rect 244280 130432 244332 130484
rect 278688 130432 278740 130484
rect 302240 130432 302292 130484
rect 343548 130432 343600 130484
rect 357440 130432 357492 130484
rect 373724 130432 373776 130484
rect 374736 130432 374788 130484
rect 404360 130432 404412 130484
rect 440148 130432 440200 130484
rect 466460 130432 466512 130484
rect 503628 130432 503680 130484
rect 517612 130432 517664 130484
rect 48872 130364 48924 130416
rect 59176 130364 59228 130416
rect 92480 130364 92532 130416
rect 198004 130364 198056 130416
rect 214564 130364 214616 130416
rect 215668 130364 215720 130416
rect 218520 130364 218572 130416
rect 256700 130364 256752 130416
rect 274732 130364 274784 130416
rect 300768 130364 300820 130416
rect 351736 130364 351788 130416
rect 358084 130364 358136 130416
rect 358728 130364 358780 130416
rect 510620 130364 510672 130416
rect 48136 130296 48188 130348
rect 51632 130296 51684 130348
rect 77300 130296 77352 130348
rect 215760 130296 215812 130348
rect 236000 130296 236052 130348
rect 372528 130296 372580 130348
rect 374828 130296 374880 130348
rect 397460 130296 397512 130348
rect 46572 130228 46624 130280
rect 54208 130228 54260 130280
rect 76012 130228 76064 130280
rect 218612 130228 218664 130280
rect 236092 130228 236144 130280
rect 378692 130228 378744 130280
rect 396172 130228 396224 130280
rect 48228 130160 48280 130212
rect 54668 130160 54720 130212
rect 75920 130160 75972 130212
rect 217232 130160 217284 130212
rect 255320 130160 255372 130212
rect 378600 130160 378652 130212
rect 396080 130160 396132 130212
rect 375104 130092 375156 130144
rect 378876 130092 378928 130144
rect 380164 130092 380216 130144
rect 375656 130024 375708 130076
rect 380256 130024 380308 130076
rect 376392 129820 376444 129872
rect 379060 129820 379112 129872
rect 219532 129752 219584 129804
rect 219716 129752 219768 129804
rect 374644 129752 374696 129804
rect 375656 129752 375708 129804
rect 375932 129752 375984 129804
rect 376484 129752 376536 129804
rect 378968 129752 379020 129804
rect 379980 129752 380032 129804
rect 50528 129684 50580 129736
rect 54484 129684 54536 129736
rect 54576 129684 54628 129736
rect 55864 129684 55916 129736
rect 213460 129684 213512 129736
rect 215944 129684 215996 129736
rect 300768 129684 300820 129736
rect 356612 129684 356664 129736
rect 373080 129684 373132 129736
rect 376116 129684 376168 129736
rect 376576 129684 376628 129736
rect 466460 129684 466512 129736
rect 516600 129684 516652 129736
rect 212908 129616 212960 129668
rect 215852 129616 215904 129668
rect 302240 129004 302292 129056
rect 356796 129004 356848 129056
rect 357532 129004 357584 129056
rect 375748 128664 375800 128716
rect 376576 128664 376628 128716
rect 215852 127576 215904 127628
rect 215944 127372 215996 127424
rect 2964 120028 3016 120080
rect 11704 120028 11756 120080
rect 57796 81404 57848 81456
rect 59360 81404 59412 81456
rect 366456 55156 366508 55208
rect 376944 55156 376996 55208
rect 214564 53116 214616 53168
rect 215208 53116 215260 53168
rect 216680 53116 216732 53168
rect 358728 53048 358780 53100
rect 376944 53048 376996 53100
rect 358084 52436 358136 52488
rect 358728 52436 358780 52488
rect 378692 44684 378744 44736
rect 397092 44684 397144 44736
rect 378600 44616 378652 44668
rect 396080 44616 396132 44668
rect 218612 44548 218664 44600
rect 236000 44548 236052 44600
rect 374644 44548 374696 44600
rect 403072 44548 403124 44600
rect 54208 44480 54260 44532
rect 77116 44480 77168 44532
rect 215760 44480 215812 44532
rect 237104 44480 237156 44532
rect 379888 44480 379940 44532
rect 414572 44480 414624 44532
rect 55956 44412 56008 44464
rect 83096 44412 83148 44464
rect 214472 44412 214524 44464
rect 243084 44412 243136 44464
rect 377220 44412 377272 44464
rect 416964 44412 417016 44464
rect 58992 44344 59044 44396
rect 101772 44344 101824 44396
rect 217232 44344 217284 44396
rect 255872 44344 255924 44396
rect 376208 44344 376260 44396
rect 419448 44344 419500 44396
rect 54852 44276 54904 44328
rect 100760 44276 100812 44328
rect 218520 44276 218572 44328
rect 256976 44276 257028 44328
rect 374920 44276 374972 44328
rect 418160 44276 418212 44328
rect 54392 44208 54444 44260
rect 143540 44208 143592 44260
rect 217140 44208 217192 44260
rect 258080 44208 258132 44260
rect 379704 44208 379756 44260
rect 423956 44208 424008 44260
rect 51448 44140 51500 44192
rect 145932 44140 145984 44192
rect 216128 44140 216180 44192
rect 262864 44140 262916 44192
rect 363604 44140 363656 44192
rect 410708 44140 410760 44192
rect 57888 44072 57940 44124
rect 215208 44072 215260 44124
rect 358084 44072 358136 44124
rect 376392 44072 376444 44124
rect 406476 44072 406528 44124
rect 3424 44004 3476 44056
rect 7564 44004 7616 44056
rect 54484 44004 54536 44056
rect 84200 44004 84252 44056
rect 215852 44004 215904 44056
rect 244280 44004 244332 44056
rect 374736 44004 374788 44056
rect 405464 44004 405516 44056
rect 59820 43936 59872 43988
rect 94504 43936 94556 43988
rect 218888 43936 218940 43988
rect 259460 43936 259512 43988
rect 379244 43936 379296 43988
rect 420644 43936 420696 43988
rect 57060 43868 57112 43920
rect 96988 43868 97040 43920
rect 219624 43868 219676 43920
rect 263876 43868 263928 43920
rect 376300 43868 376352 43920
rect 421748 43868 421800 43920
rect 54944 43800 54996 43852
rect 98092 43800 98144 43852
rect 216220 43800 216272 43852
rect 261760 43800 261812 43852
rect 379796 43800 379848 43852
rect 425244 43800 425296 43852
rect 56048 43732 56100 43784
rect 102784 43732 102836 43784
rect 214196 43732 214248 43784
rect 260656 43732 260708 43784
rect 279240 43732 279292 43784
rect 356980 43732 357032 43784
rect 375840 43732 375892 43784
rect 422852 43732 422904 43784
rect 56324 43664 56376 43716
rect 103888 43664 103940 43716
rect 212448 43664 212500 43716
rect 308496 43664 308548 43716
rect 356704 43664 356756 43716
rect 425980 43664 426032 43716
rect 53288 43596 53340 43648
rect 113272 43596 113324 43648
rect 213736 43596 213788 43648
rect 315856 43596 315908 43648
rect 366364 43596 366416 43648
rect 458456 43596 458508 43648
rect 42524 43528 42576 43580
rect 115940 43528 115992 43580
rect 219256 43528 219308 43580
rect 421012 43528 421064 43580
rect 56232 43460 56284 43512
rect 158444 43460 158496 43512
rect 198648 43460 198700 43512
rect 300860 43460 300912 43512
rect 358176 43460 358228 43512
rect 455880 43460 455932 43512
rect 49608 43392 49660 43444
rect 160836 43392 160888 43444
rect 218980 43392 219032 43444
rect 428188 43392 428240 43444
rect 439228 43392 439280 43444
rect 516600 43392 516652 43444
rect 378876 43324 378928 43376
rect 407580 43324 407632 43376
rect 375932 43256 375984 43308
rect 404176 43256 404228 43308
rect 57244 42780 57296 42832
rect 57888 42780 57940 42832
rect 50988 42712 51040 42764
rect 155960 42712 156012 42764
rect 183468 42712 183520 42764
rect 197452 42712 197504 42764
rect 209596 42712 209648 42764
rect 320916 42712 320968 42764
rect 343180 42712 343232 42764
rect 357624 42712 357676 42764
rect 378508 42712 378560 42764
rect 485964 42712 486016 42764
rect 503260 42712 503312 42764
rect 517612 42712 517664 42764
rect 52276 42644 52328 42696
rect 135904 42644 135956 42696
rect 183192 42644 183244 42696
rect 197360 42644 197412 42696
rect 218244 42644 218296 42696
rect 325884 42644 325936 42696
rect 343456 42644 343508 42696
rect 357440 42644 357492 42696
rect 365076 42644 365128 42696
rect 453396 42644 453448 42696
rect 503536 42644 503588 42696
rect 517520 42644 517572 42696
rect 53748 42576 53800 42628
rect 133420 42576 133472 42628
rect 216588 42576 216640 42628
rect 318340 42576 318392 42628
rect 360936 42576 360988 42628
rect 448244 42576 448296 42628
rect 56508 42508 56560 42560
rect 128360 42508 128412 42560
rect 211068 42508 211120 42560
rect 310980 42508 311032 42560
rect 364984 42508 365036 42560
rect 445852 42508 445904 42560
rect 55128 42440 55180 42492
rect 118240 42440 118292 42492
rect 213828 42440 213880 42492
rect 313372 42440 313424 42492
rect 367744 42440 367796 42492
rect 443460 42440 443512 42492
rect 52368 42372 52420 42424
rect 113180 42372 113232 42424
rect 215116 42372 215168 42424
rect 298468 42372 298520 42424
rect 361028 42372 361080 42424
rect 435916 42372 435968 42424
rect 43996 42304 44048 42356
rect 96252 42304 96304 42356
rect 209688 42304 209740 42356
rect 293316 42304 293368 42356
rect 370504 42304 370556 42356
rect 440884 42304 440936 42356
rect 59912 42236 59964 42288
rect 108580 42236 108632 42288
rect 218428 42236 218480 42288
rect 302516 42236 302568 42288
rect 371884 42236 371936 42288
rect 438492 42236 438544 42288
rect 56140 42168 56192 42220
rect 95884 42168 95936 42220
rect 211804 42168 211856 42220
rect 276112 42168 276164 42220
rect 278320 42168 278372 42220
rect 356796 42168 356848 42220
rect 378784 42168 378836 42220
rect 430948 42168 431000 42220
rect 50160 42100 50212 42152
rect 88340 42100 88392 42152
rect 218704 42100 218756 42152
rect 268200 42100 268252 42152
rect 363696 42100 363748 42152
rect 413652 42100 413704 42152
rect 54668 42032 54720 42084
rect 76012 42032 76064 42084
rect 211896 42032 211948 42084
rect 260932 42032 260984 42084
rect 379612 42032 379664 42084
rect 427636 42032 427688 42084
rect 378968 41964 379020 42016
rect 415492 41964 415544 42016
rect 52092 41352 52144 41404
rect 115756 41352 115808 41404
rect 219992 41352 220044 41404
rect 408316 41352 408368 41404
rect 57796 41284 57848 41336
rect 119068 41284 119120 41336
rect 216496 41284 216548 41336
rect 276940 41284 276992 41336
rect 376116 41284 376168 41336
rect 429660 41284 429712 41336
rect 53564 41216 53616 41268
rect 114192 41216 114244 41268
rect 214380 41216 214432 41268
rect 273260 41216 273312 41268
rect 379428 41216 379480 41268
rect 426440 41216 426492 41268
rect 42616 41148 42668 41200
rect 93676 41148 93728 41200
rect 214932 41148 214984 41200
rect 271236 41148 271288 41200
rect 379152 41148 379204 41200
rect 413284 41148 413336 41200
rect 58624 41080 58676 41132
rect 107016 41080 107068 41132
rect 212264 41080 212316 41132
rect 268476 41080 268528 41132
rect 377680 41080 377732 41132
rect 409972 41080 410024 41132
rect 60004 41012 60056 41064
rect 106372 41012 106424 41064
rect 219348 41012 219400 41064
rect 265164 41012 265216 41064
rect 373908 41012 373960 41064
rect 401692 41012 401744 41064
rect 51724 40944 51776 40996
rect 85396 40944 85448 40996
rect 218796 40944 218848 40996
rect 253388 40944 253440 40996
rect 374828 40944 374880 40996
rect 398196 40944 398248 40996
rect 53380 40876 53432 40928
rect 86500 40876 86552 40928
rect 219072 40876 219124 40928
rect 251180 40876 251232 40928
rect 59084 40808 59136 40860
rect 92388 40808 92440 40860
rect 216036 40808 216088 40860
rect 246396 40808 246448 40860
rect 55864 40740 55916 40792
rect 87604 40740 87656 40792
rect 214656 40740 214708 40792
rect 245292 40740 245344 40792
rect 51632 40672 51684 40724
rect 78220 40672 78272 40724
rect 213368 40672 213420 40724
rect 239128 40672 239180 40724
rect 53472 40604 53524 40656
rect 80428 40604 80480 40656
rect 215024 40604 215076 40656
rect 241612 40604 241664 40656
rect 54760 39992 54812 40044
rect 116308 39992 116360 40044
rect 213644 39992 213696 40044
rect 240508 39992 240560 40044
rect 375196 39992 375248 40044
rect 399392 39992 399444 40044
rect 52000 39924 52052 39976
rect 111892 39924 111944 39976
rect 214840 39924 214892 39976
rect 238116 39924 238168 39976
rect 376668 39924 376720 39976
rect 436376 39924 436428 39976
rect 52184 39856 52236 39908
rect 111156 39856 111208 39908
rect 216404 39856 216456 39908
rect 272156 39856 272208 39908
rect 374460 39856 374512 39908
rect 434628 39856 434680 39908
rect 55036 39788 55088 39840
rect 109316 39788 109368 39840
rect 215944 39788 215996 39840
rect 269764 39788 269816 39840
rect 373816 39788 373868 39840
rect 432144 39788 432196 39840
rect 44088 39720 44140 39772
rect 90732 39720 90784 39772
rect 219808 39720 219860 39772
rect 266636 39720 266688 39772
rect 375288 39720 375340 39772
rect 431132 39720 431184 39772
rect 56968 39652 57020 39704
rect 91284 39652 91336 39704
rect 219900 39652 219952 39704
rect 266360 39652 266412 39704
rect 377588 39652 377640 39704
rect 411904 39652 411956 39704
rect 59176 39584 59228 39636
rect 93308 39584 93360 39636
rect 219716 39584 219768 39636
rect 254124 39584 254176 39636
rect 379336 39584 379388 39636
rect 411260 39584 411312 39636
rect 56416 39516 56468 39568
rect 88616 39516 88668 39568
rect 217600 39516 217652 39568
rect 251732 39516 251784 39568
rect 376576 39516 376628 39568
rect 408684 39516 408736 39568
rect 59268 39448 59320 39500
rect 89996 39448 90048 39500
rect 216312 39448 216364 39500
rect 248604 39448 248656 39500
rect 372436 39448 372488 39500
rect 400312 39448 400364 39500
rect 53656 39380 53708 39432
rect 81808 39380 81860 39432
rect 219164 39380 219216 39432
rect 247684 39380 247736 39432
rect 375012 39380 375064 39432
rect 435180 39380 435232 39432
rect 51908 39312 51960 39364
rect 78772 39312 78824 39364
rect 213552 39312 213604 39364
rect 274732 39312 274784 39364
rect 212356 39244 212408 39296
rect 273536 39244 273588 39296
rect 2780 31696 2832 31748
rect 580448 31696 580500 31748
rect 1676 3476 1728 3528
rect 2780 3476 2832 3528
rect 572 3408 624 3460
rect 57244 3408 57296 3460
<< metal2 >>
rect 7626 703520 7738 704960
rect 22990 703520 23102 704960
rect 38354 703520 38466 704960
rect 53718 703520 53830 704960
rect 69082 703520 69194 704960
rect 84446 703520 84558 704960
rect 99810 703520 99922 704960
rect 115174 703520 115286 704960
rect 130538 703520 130650 704960
rect 145902 703520 146014 704960
rect 161266 703520 161378 704960
rect 176630 703520 176742 704960
rect 191994 703520 192106 704960
rect 207358 703520 207470 704960
rect 222722 703520 222834 704960
rect 238086 703520 238198 704960
rect 253450 703520 253562 704960
rect 268814 703520 268926 704960
rect 284178 703520 284290 704960
rect 299634 703520 299746 704960
rect 314998 703520 315110 704960
rect 330362 703520 330474 704960
rect 345726 703520 345838 704960
rect 361090 703520 361202 704960
rect 375392 703582 376340 703610
rect 38396 701010 38424 703520
rect 38384 701004 38436 701010
rect 38384 700946 38436 700952
rect 38396 699718 38424 700946
rect 69124 700330 69152 703520
rect 99852 701010 99880 703520
rect 130580 702434 130608 703520
rect 129752 702406 130608 702434
rect 99840 701004 99892 701010
rect 99840 700946 99892 700952
rect 69112 700324 69164 700330
rect 69112 700266 69164 700272
rect 37924 699712 37976 699718
rect 37924 699654 37976 699660
rect 38384 699712 38436 699718
rect 38384 699654 38436 699660
rect 3422 685128 3478 685137
rect 3422 685063 3478 685072
rect 3436 684554 3464 685063
rect 3424 684548 3476 684554
rect 3424 684490 3476 684496
rect 37936 660346 37964 699654
rect 59268 697604 59320 697610
rect 59268 697546 59320 697552
rect 2780 660340 2832 660346
rect 2780 660282 2832 660288
rect 37924 660340 37976 660346
rect 37924 660282 37976 660288
rect 2792 659977 2820 660282
rect 2778 659968 2834 659977
rect 2778 659903 2834 659912
rect 2792 609657 2820 659903
rect 40684 645992 40736 645998
rect 40684 645934 40736 645940
rect 3422 634808 3478 634817
rect 3422 634743 3478 634752
rect 2778 609648 2834 609657
rect 2778 609583 2834 609592
rect 2792 559337 2820 609583
rect 3436 569226 3464 634743
rect 3514 584488 3570 584497
rect 3514 584423 3570 584432
rect 3528 575482 3556 584423
rect 3516 575476 3568 575482
rect 3516 575418 3568 575424
rect 7564 570648 7616 570654
rect 7564 570590 7616 570596
rect 3424 569220 3476 569226
rect 3424 569162 3476 569168
rect 2778 559328 2834 559337
rect 2778 559263 2834 559272
rect 2792 509153 2820 559263
rect 3422 554840 3478 554849
rect 3422 554775 3478 554784
rect 3436 521665 3464 554775
rect 3422 521656 3478 521665
rect 3422 521591 3478 521600
rect 2778 509144 2834 509153
rect 2778 509079 2834 509088
rect 2792 458833 2820 509079
rect 3608 472660 3660 472666
rect 3608 472602 3660 472608
rect 3516 471980 3568 471986
rect 3516 471922 3568 471928
rect 3528 471345 3556 471922
rect 3514 471336 3570 471345
rect 3514 471271 3570 471280
rect 3620 470594 3648 472602
rect 3528 470566 3648 470594
rect 2778 458824 2834 458833
rect 2778 458759 2834 458768
rect 2792 408513 2820 458759
rect 3528 451274 3556 470566
rect 4804 469872 4856 469878
rect 4804 469814 4856 469820
rect 3436 451246 3556 451274
rect 3148 422272 3200 422278
rect 3148 422214 3200 422220
rect 3160 421161 3188 422214
rect 3146 421152 3202 421161
rect 3146 421087 3202 421096
rect 2778 408504 2834 408513
rect 2778 408439 2834 408448
rect 2792 358329 2820 408439
rect 2778 358320 2834 358329
rect 2778 358255 2834 358264
rect 2792 308009 2820 358255
rect 2778 308000 2834 308009
rect 2778 307935 2834 307944
rect 2792 257689 2820 307935
rect 2778 257680 2834 257689
rect 2778 257615 2834 257624
rect 2792 207369 2820 257615
rect 2778 207360 2834 207369
rect 2778 207295 2834 207304
rect 2792 157185 2820 207295
rect 2872 169720 2924 169726
rect 2870 169688 2872 169697
rect 2924 169688 2926 169697
rect 2870 169623 2926 169632
rect 2778 157176 2834 157185
rect 2778 157111 2834 157120
rect 2792 106865 2820 157111
rect 2964 120080 3016 120086
rect 2964 120022 3016 120028
rect 2976 119377 3004 120022
rect 2962 119368 3018 119377
rect 2962 119303 3018 119312
rect 2778 106856 2834 106865
rect 2778 106791 2834 106800
rect 2792 69193 2820 106791
rect 3436 81705 3464 451246
rect 3516 371204 3568 371210
rect 3516 371146 3568 371152
rect 3528 370841 3556 371146
rect 3514 370832 3570 370841
rect 3514 370767 3570 370776
rect 4816 169726 4844 469814
rect 4804 169720 4856 169726
rect 4804 169662 4856 169668
rect 3422 81696 3478 81705
rect 3422 81631 3478 81640
rect 2778 69184 2834 69193
rect 2778 69119 2834 69128
rect 2792 31754 2820 69119
rect 7576 44062 7604 570590
rect 11704 567248 11756 567254
rect 11704 567190 11756 567196
rect 11716 120086 11744 567190
rect 18604 468512 18656 468518
rect 18604 468454 18656 468460
rect 18616 422278 18644 468454
rect 18604 422272 18656 422278
rect 18604 422214 18656 422220
rect 40696 371210 40724 645934
rect 56508 640620 56560 640626
rect 56508 640562 56560 640568
rect 54944 640552 54996 640558
rect 54944 640494 54996 640500
rect 54852 640484 54904 640490
rect 54852 640426 54904 640432
rect 54864 574938 54892 640426
rect 54852 574932 54904 574938
rect 54852 574874 54904 574880
rect 54956 557122 54984 640494
rect 55128 640416 55180 640422
rect 55128 640358 55180 640364
rect 55036 640348 55088 640354
rect 55036 640290 55088 640296
rect 55048 557326 55076 640290
rect 55140 557462 55168 640358
rect 56324 637832 56376 637838
rect 56324 637774 56376 637780
rect 55128 557456 55180 557462
rect 55128 557398 55180 557404
rect 55036 557320 55088 557326
rect 55036 557262 55088 557268
rect 54944 557116 54996 557122
rect 54944 557058 54996 557064
rect 56336 556918 56364 637774
rect 56416 637696 56468 637702
rect 56416 637638 56468 637644
rect 56428 557258 56456 637638
rect 56520 557394 56548 640562
rect 57796 637900 57848 637906
rect 57796 637842 57848 637848
rect 57426 635624 57482 635633
rect 57426 635559 57482 635568
rect 57242 602304 57298 602313
rect 57242 602239 57298 602248
rect 57150 586664 57206 586673
rect 57150 586599 57206 586608
rect 57058 580544 57114 580553
rect 57058 580479 57114 580488
rect 57072 567934 57100 580479
rect 57164 573578 57192 586599
rect 57256 575550 57284 602239
rect 57440 600302 57468 635559
rect 57702 629504 57758 629513
rect 57702 629439 57758 629448
rect 57610 626784 57666 626793
rect 57610 626719 57666 626728
rect 57518 608424 57574 608433
rect 57518 608359 57574 608368
rect 57428 600296 57480 600302
rect 57428 600238 57480 600244
rect 57334 598904 57390 598913
rect 57334 598839 57390 598848
rect 57244 575544 57296 575550
rect 57244 575486 57296 575492
rect 57152 573572 57204 573578
rect 57152 573514 57204 573520
rect 57348 570790 57376 598839
rect 57426 596184 57482 596193
rect 57426 596119 57482 596128
rect 57336 570784 57388 570790
rect 57336 570726 57388 570732
rect 57060 567928 57112 567934
rect 57060 567870 57112 567876
rect 57440 558210 57468 596119
rect 57532 559774 57560 608359
rect 57624 574870 57652 626719
rect 57612 574864 57664 574870
rect 57612 574806 57664 574812
rect 57716 565146 57744 629439
rect 57704 565140 57756 565146
rect 57704 565082 57756 565088
rect 57520 559768 57572 559774
rect 57520 559710 57572 559716
rect 57428 558204 57480 558210
rect 57428 558146 57480 558152
rect 56508 557388 56560 557394
rect 56508 557330 56560 557336
rect 56416 557252 56468 557258
rect 56416 557194 56468 557200
rect 56324 556912 56376 556918
rect 56324 556854 56376 556860
rect 57808 556850 57836 637842
rect 59176 637628 59228 637634
rect 59176 637570 59228 637576
rect 59082 632904 59138 632913
rect 59082 632839 59138 632848
rect 58898 623384 58954 623393
rect 58898 623319 58954 623328
rect 58530 617264 58586 617273
rect 58530 617199 58586 617208
rect 57886 611144 57942 611153
rect 57886 611079 57942 611088
rect 57900 576230 57928 611079
rect 58438 590064 58494 590073
rect 58438 589999 58494 590008
rect 57888 576224 57940 576230
rect 57888 576166 57940 576172
rect 57796 556844 57848 556850
rect 57796 556786 57848 556792
rect 57900 528554 57928 576166
rect 58452 575278 58480 589999
rect 58440 575272 58492 575278
rect 58440 575214 58492 575220
rect 58544 562426 58572 617199
rect 58806 605024 58862 605033
rect 58806 604959 58862 604968
rect 58624 600296 58676 600302
rect 58624 600238 58676 600244
rect 58532 562420 58584 562426
rect 58532 562362 58584 562368
rect 58636 557054 58664 600238
rect 58714 583944 58770 583953
rect 58714 583879 58770 583888
rect 58728 559570 58756 583879
rect 58820 574326 58848 604959
rect 58808 574320 58860 574326
rect 58808 574262 58860 574268
rect 58912 572014 58940 623319
rect 58990 620664 59046 620673
rect 58990 620599 59046 620608
rect 58900 572008 58952 572014
rect 58900 571950 58952 571956
rect 59004 566574 59032 620599
rect 59096 569430 59124 632839
rect 59084 569424 59136 569430
rect 59084 569366 59136 569372
rect 58992 566568 59044 566574
rect 58992 566510 59044 566516
rect 58716 559564 58768 559570
rect 58716 559506 58768 559512
rect 58624 557048 58676 557054
rect 58624 556990 58676 556996
rect 59188 556782 59216 637570
rect 59280 614553 59308 697546
rect 129752 650690 129780 702406
rect 161308 701010 161336 703520
rect 161296 701004 161348 701010
rect 161296 700946 161348 700952
rect 192036 683114 192064 703520
rect 222764 701010 222792 703520
rect 222752 701004 222804 701010
rect 222752 700946 222804 700952
rect 253492 700398 253520 703520
rect 284220 701010 284248 703520
rect 284208 701004 284260 701010
rect 284208 700946 284260 700952
rect 253480 700392 253532 700398
rect 253480 700334 253532 700340
rect 305644 700392 305696 700398
rect 305644 700334 305696 700340
rect 304264 700324 304316 700330
rect 304264 700266 304316 700272
rect 191852 683086 192064 683114
rect 137560 658300 137612 658306
rect 137560 658242 137612 658248
rect 129740 650684 129792 650690
rect 129740 650626 129792 650632
rect 136548 640892 136600 640898
rect 136548 640834 136600 640840
rect 134892 640824 134944 640830
rect 134892 640766 134944 640772
rect 100576 640756 100628 640762
rect 100576 640698 100628 640704
rect 124496 640756 124548 640762
rect 124496 640698 124548 640704
rect 77392 640620 77444 640626
rect 77392 640562 77444 640568
rect 69020 638988 69072 638994
rect 69020 638930 69072 638936
rect 69032 638044 69060 638930
rect 77404 638044 77432 640562
rect 80612 640552 80664 640558
rect 80612 640494 80664 640500
rect 80624 638044 80652 640494
rect 88984 640484 89036 640490
rect 88984 640426 89036 640432
rect 88996 638044 89024 640426
rect 92204 640416 92256 640422
rect 92204 640358 92256 640364
rect 92216 638044 92244 640358
rect 94780 640348 94832 640354
rect 94780 640290 94832 640296
rect 94792 638044 94820 640290
rect 100588 638044 100616 640698
rect 115388 640688 115440 640694
rect 115388 640630 115440 640636
rect 112168 640620 112220 640626
rect 112168 640562 112220 640568
rect 109592 640552 109644 640558
rect 109592 640494 109644 640500
rect 106372 640484 106424 640490
rect 106372 640426 106424 640432
rect 103796 640416 103848 640422
rect 103796 640358 103848 640364
rect 103808 638044 103836 640358
rect 106384 638044 106412 640426
rect 109604 638044 109632 640494
rect 112180 638044 112208 640562
rect 115400 638044 115428 640630
rect 122840 640552 122892 640558
rect 122840 640494 122892 640500
rect 121460 640484 121512 640490
rect 121460 640426 121512 640432
rect 120816 640416 120868 640422
rect 120816 640358 120868 640364
rect 71240 637906 71622 637922
rect 71228 637900 71622 637906
rect 71280 637894 71622 637900
rect 71228 637842 71280 637848
rect 65524 637832 65576 637838
rect 65576 637780 65826 637786
rect 65524 637774 65826 637780
rect 59360 637764 59412 637770
rect 65536 637758 65826 637774
rect 97920 637770 98026 637786
rect 97908 637764 98026 637770
rect 59360 637706 59412 637712
rect 97960 637758 98026 637764
rect 97908 637706 97960 637712
rect 59266 614544 59322 614553
rect 59266 614479 59322 614488
rect 59266 592784 59322 592793
rect 59266 592719 59322 592728
rect 59280 573510 59308 592719
rect 59268 573504 59320 573510
rect 59268 573446 59320 573452
rect 59372 557534 59400 637706
rect 62948 637696 63000 637702
rect 86776 637696 86828 637702
rect 63000 637644 63250 637650
rect 62948 637638 63250 637644
rect 62960 637622 63250 637638
rect 74644 637634 74842 637650
rect 74632 637628 74842 637634
rect 74684 637622 74842 637628
rect 83214 637634 83504 637650
rect 86434 637644 86776 637650
rect 86434 637638 86828 637644
rect 83214 637628 83516 637634
rect 83214 637622 83464 637628
rect 74632 637570 74684 637576
rect 86434 637622 86816 637638
rect 117990 637634 118280 637650
rect 117990 637628 118292 637634
rect 117990 637622 118240 637628
rect 83464 637570 83516 637576
rect 118240 637570 118292 637576
rect 59464 637350 60030 637378
rect 120566 637350 120764 637378
rect 59464 573918 59492 637350
rect 59542 577788 59598 577797
rect 59542 577723 59598 577732
rect 59452 573912 59504 573918
rect 59452 573854 59504 573860
rect 59556 563786 59584 577723
rect 60372 575544 60424 575550
rect 60372 575486 60424 575492
rect 60016 571402 60044 575076
rect 60004 571396 60056 571402
rect 60004 571338 60056 571344
rect 59544 563780 59596 563786
rect 59544 563722 59596 563728
rect 59372 557506 60320 557534
rect 59176 556776 59228 556782
rect 59176 556718 59228 556724
rect 60292 554963 60320 557506
rect 60384 557190 60412 575486
rect 62396 575272 62448 575278
rect 62396 575214 62448 575220
rect 60924 574320 60976 574326
rect 60924 574262 60976 574268
rect 60372 557184 60424 557190
rect 60372 557126 60424 557132
rect 60936 554963 60964 574262
rect 61384 571396 61436 571402
rect 61384 571338 61436 571344
rect 61396 561134 61424 571338
rect 61384 561128 61436 561134
rect 61384 561070 61436 561076
rect 61660 557524 61712 557530
rect 61660 557466 61712 557472
rect 61672 554963 61700 557466
rect 62408 554963 62436 575214
rect 106280 575136 106332 575142
rect 62592 572218 62620 575076
rect 64892 575062 65182 575090
rect 63500 574796 63552 574802
rect 63500 574738 63552 574744
rect 63224 573912 63276 573918
rect 63224 573854 63276 573860
rect 62580 572212 62632 572218
rect 62580 572154 62632 572160
rect 63132 562352 63184 562358
rect 63132 562294 63184 562300
rect 63144 554963 63172 562294
rect 63236 556986 63264 573854
rect 63512 557534 63540 574738
rect 64512 573368 64564 573374
rect 64512 573310 64564 573316
rect 63512 557506 63816 557534
rect 63224 556980 63276 556986
rect 63224 556922 63276 556928
rect 63788 554963 63816 557506
rect 64524 554963 64552 573310
rect 64892 557530 64920 575062
rect 67640 573436 67692 573442
rect 67640 573378 67692 573384
rect 65984 570716 66036 570722
rect 65984 570658 66036 570664
rect 65248 566500 65300 566506
rect 65248 566442 65300 566448
rect 64880 557524 64932 557530
rect 64880 557466 64932 557472
rect 65260 554963 65288 566442
rect 65996 554963 66024 570658
rect 66720 563712 66772 563718
rect 66720 563654 66772 563660
rect 66732 554963 66760 563654
rect 67652 557534 67680 573378
rect 68388 572150 68416 575076
rect 68836 573504 68888 573510
rect 68836 573446 68888 573452
rect 68376 572144 68428 572150
rect 68376 572086 68428 572092
rect 67652 557506 68140 557534
rect 67364 557456 67416 557462
rect 67364 557398 67416 557404
rect 67376 554963 67404 557398
rect 68112 554963 68140 557506
rect 68376 557456 68428 557462
rect 68376 557398 68428 557404
rect 68388 557054 68416 557398
rect 68376 557048 68428 557054
rect 68376 556990 68428 556996
rect 68468 557048 68520 557054
rect 68468 556990 68520 556996
rect 68480 556782 68508 556990
rect 68468 556776 68520 556782
rect 68468 556718 68520 556724
rect 68848 554963 68876 573446
rect 70964 572082 70992 575076
rect 71044 572212 71096 572218
rect 71044 572154 71096 572160
rect 70952 572076 71004 572082
rect 70952 572018 71004 572024
rect 69020 569288 69072 569294
rect 69020 569230 69072 569236
rect 69032 562290 69060 569230
rect 70952 567860 71004 567866
rect 70952 567802 71004 567808
rect 69020 562284 69072 562290
rect 69020 562226 69072 562232
rect 70308 562284 70360 562290
rect 70308 562226 70360 562232
rect 69572 561060 69624 561066
rect 69572 561002 69624 561008
rect 69584 554963 69612 561002
rect 70320 554963 70348 562226
rect 70964 554963 70992 567802
rect 71056 565214 71084 572154
rect 74184 571402 74212 575076
rect 74540 572280 74592 572286
rect 74540 572222 74592 572228
rect 72424 571396 72476 571402
rect 72424 571338 72476 571344
rect 74172 571396 74224 571402
rect 74172 571338 74224 571344
rect 71044 565208 71096 565214
rect 71044 565150 71096 565156
rect 71688 560992 71740 560998
rect 71688 560934 71740 560940
rect 71700 554963 71728 560934
rect 72436 554963 72464 571338
rect 74552 562290 74580 572222
rect 74632 572008 74684 572014
rect 74632 571950 74684 571956
rect 74540 562284 74592 562290
rect 74540 562226 74592 562232
rect 73160 559700 73212 559706
rect 73160 559642 73212 559648
rect 73172 554963 73200 559642
rect 73804 556844 73856 556850
rect 73804 556786 73856 556792
rect 73816 554963 73844 556786
rect 74644 555234 74672 571950
rect 76760 571402 76788 575076
rect 78680 574932 78732 574938
rect 78680 574874 78732 574880
rect 76840 572008 76892 572014
rect 76840 571950 76892 571956
rect 76748 571396 76800 571402
rect 76748 571338 76800 571344
rect 76852 567194 76880 571950
rect 76760 567166 76880 567194
rect 75276 562284 75328 562290
rect 75276 562226 75328 562232
rect 74568 555206 74672 555234
rect 74568 554948 74596 555206
rect 75288 554963 75316 562226
rect 76012 556980 76064 556986
rect 76012 556922 76064 556928
rect 76024 554963 76052 556922
rect 76760 554963 76788 567166
rect 76840 565140 76892 565146
rect 76840 565082 76892 565088
rect 76852 556986 76880 565082
rect 78692 562290 78720 574874
rect 78864 573504 78916 573510
rect 78864 573446 78916 573452
rect 78680 562284 78732 562290
rect 78680 562226 78732 562232
rect 77392 557456 77444 557462
rect 77392 557398 77444 557404
rect 76840 556980 76892 556986
rect 76840 556922 76892 556928
rect 77404 554963 77432 557398
rect 78128 556844 78180 556850
rect 78128 556786 78180 556792
rect 78140 554963 78168 556786
rect 78876 554963 78904 573446
rect 79980 569362 80008 575076
rect 81716 573572 81768 573578
rect 81716 573514 81768 573520
rect 79968 569356 80020 569362
rect 79968 569298 80020 569304
rect 80336 565140 80388 565146
rect 80336 565082 80388 565088
rect 79600 562284 79652 562290
rect 79600 562226 79652 562232
rect 79612 554963 79640 562226
rect 80348 554963 80376 565082
rect 80980 563848 81032 563854
rect 80980 563790 81032 563796
rect 80992 554963 81020 563790
rect 81728 554963 81756 573514
rect 82556 572354 82584 575076
rect 83188 574864 83240 574870
rect 83188 574806 83240 574812
rect 82544 572348 82596 572354
rect 82544 572290 82596 572296
rect 82452 559632 82504 559638
rect 82452 559574 82504 559580
rect 82464 554963 82492 559574
rect 83200 554963 83228 574806
rect 85776 572218 85804 575076
rect 88156 573640 88208 573646
rect 88156 573582 88208 573588
rect 86960 573572 87012 573578
rect 86960 573514 87012 573520
rect 85764 572212 85816 572218
rect 85764 572154 85816 572160
rect 83464 571396 83516 571402
rect 83464 571338 83516 571344
rect 83476 557530 83504 571338
rect 84568 566704 84620 566710
rect 84568 566646 84620 566652
rect 83464 557524 83516 557530
rect 83464 557466 83516 557472
rect 83924 557388 83976 557394
rect 83924 557330 83976 557336
rect 83936 554963 83964 557330
rect 84580 554963 84608 566646
rect 86040 562488 86092 562494
rect 86040 562430 86092 562436
rect 85304 557320 85356 557326
rect 85304 557262 85356 557268
rect 85316 554963 85344 557262
rect 86052 554963 86080 562430
rect 86972 557534 87000 573514
rect 86776 557524 86828 557530
rect 86972 557506 87460 557534
rect 86776 557466 86828 557472
rect 86788 554963 86816 557466
rect 87432 554963 87460 557506
rect 88168 554963 88196 573582
rect 88352 565282 88380 575076
rect 88984 572348 89036 572354
rect 88984 572290 89036 572296
rect 88340 565276 88392 565282
rect 88340 565218 88392 565224
rect 88248 559768 88300 559774
rect 88248 559710 88300 559716
rect 88260 556306 88288 559710
rect 88892 557252 88944 557258
rect 88892 557194 88944 557200
rect 88248 556300 88300 556306
rect 88248 556242 88300 556248
rect 88904 554963 88932 557194
rect 88996 556510 89024 572290
rect 91572 571402 91600 575076
rect 93860 574864 93912 574870
rect 93860 574806 93912 574812
rect 91560 571396 91612 571402
rect 91560 571338 91612 571344
rect 93124 571396 93176 571402
rect 93124 571338 93176 571344
rect 89812 570784 89864 570790
rect 89812 570726 89864 570732
rect 89628 563916 89680 563922
rect 89628 563858 89680 563864
rect 88984 556504 89036 556510
rect 88984 556446 89036 556452
rect 89640 554963 89668 563858
rect 89824 562358 89852 570726
rect 92572 569424 92624 569430
rect 92572 569366 92624 569372
rect 89812 562352 89864 562358
rect 89812 562294 89864 562300
rect 91008 562352 91060 562358
rect 91008 562294 91060 562300
rect 90364 556504 90416 556510
rect 90364 556446 90416 556452
rect 90376 554963 90404 556446
rect 91020 554963 91048 562294
rect 91744 556300 91796 556306
rect 91744 556242 91796 556248
rect 91756 554963 91784 556242
rect 92584 555234 92612 569366
rect 93136 557122 93164 571338
rect 93872 557534 93900 574806
rect 94148 571470 94176 575076
rect 97368 572286 97396 575076
rect 98184 575000 98236 575006
rect 98184 574942 98236 574948
rect 97448 574932 97500 574938
rect 97448 574874 97500 574880
rect 97356 572280 97408 572286
rect 97356 572222 97408 572228
rect 94136 571464 94188 571470
rect 94136 571406 94188 571412
rect 94596 570852 94648 570858
rect 94596 570794 94648 570800
rect 93872 557506 93992 557534
rect 93032 557116 93084 557122
rect 93032 557058 93084 557064
rect 93124 557116 93176 557122
rect 93124 557058 93176 557064
rect 93044 557002 93072 557058
rect 93044 556974 93256 557002
rect 92508 555206 92612 555234
rect 92508 554948 92536 555206
rect 93228 554963 93256 556974
rect 93964 554963 93992 557506
rect 94608 554963 94636 570794
rect 95332 557252 95384 557258
rect 95332 557194 95384 557200
rect 95344 554963 95372 557194
rect 96804 557116 96856 557122
rect 96804 557058 96856 557064
rect 96068 556232 96120 556238
rect 96068 556174 96120 556180
rect 96080 554963 96108 556174
rect 96816 554963 96844 557058
rect 97460 554963 97488 574874
rect 98196 554963 98224 574942
rect 99944 572286 99972 575076
rect 100392 575068 100444 575074
rect 100392 575010 100444 575016
rect 99932 572280 99984 572286
rect 99932 572222 99984 572228
rect 99196 558204 99248 558210
rect 99196 558146 99248 558152
rect 99288 558204 99340 558210
rect 99288 558146 99340 558152
rect 99208 557122 99236 558146
rect 99196 557116 99248 557122
rect 99196 557058 99248 557064
rect 98920 556912 98972 556918
rect 98920 556854 98972 556860
rect 98932 554963 98960 556854
rect 99300 556238 99328 558146
rect 99656 557048 99708 557054
rect 99656 556990 99708 556996
rect 99288 556232 99340 556238
rect 99288 556174 99340 556180
rect 99668 554963 99696 556990
rect 100404 554963 100432 575010
rect 101404 571464 101456 571470
rect 101404 571406 101456 571412
rect 100760 571396 100812 571402
rect 100760 571338 100812 571344
rect 100772 562426 100800 571338
rect 101036 563780 101088 563786
rect 101036 563722 101088 563728
rect 100760 562420 100812 562426
rect 100760 562362 100812 562368
rect 101048 554963 101076 563722
rect 101416 557462 101444 571406
rect 103164 571402 103192 575076
rect 104912 575062 105754 575090
rect 106280 575078 106332 575084
rect 103152 571396 103204 571402
rect 103152 571338 103204 571344
rect 101496 567928 101548 567934
rect 101496 567870 101548 567876
rect 101404 557456 101456 557462
rect 101404 557398 101456 557404
rect 101508 556374 101536 567870
rect 104624 565276 104676 565282
rect 104624 565218 104676 565224
rect 101772 562420 101824 562426
rect 101772 562362 101824 562368
rect 101496 556368 101548 556374
rect 101496 556310 101548 556316
rect 101784 554963 101812 562362
rect 102508 562352 102560 562358
rect 102508 562294 102560 562300
rect 102520 554963 102548 562294
rect 103980 556912 104032 556918
rect 103980 556854 104032 556860
rect 103244 556368 103296 556374
rect 103244 556310 103296 556316
rect 103256 554963 103284 556310
rect 103992 554963 104020 556854
rect 104636 554963 104664 565218
rect 104912 563922 104940 575062
rect 105544 572144 105596 572150
rect 105544 572086 105596 572092
rect 104900 563916 104952 563922
rect 104900 563858 104952 563864
rect 105360 561128 105412 561134
rect 105360 561070 105412 561076
rect 105372 554963 105400 561070
rect 105556 556782 105584 572086
rect 106292 562358 106320 575078
rect 108304 572212 108356 572218
rect 108304 572154 108356 572160
rect 106924 571396 106976 571402
rect 106924 571338 106976 571344
rect 106280 562352 106332 562358
rect 106280 562294 106332 562300
rect 106936 559706 106964 571338
rect 108212 566568 108264 566574
rect 108212 566510 108264 566516
rect 107568 562352 107620 562358
rect 107568 562294 107620 562300
rect 106924 559700 106976 559706
rect 106924 559642 106976 559648
rect 106096 557456 106148 557462
rect 106096 557398 106148 557404
rect 105544 556776 105596 556782
rect 105544 556718 105596 556724
rect 106108 554963 106136 557398
rect 106832 557048 106884 557054
rect 106832 556990 106884 556996
rect 106844 554963 106872 556990
rect 107580 554963 107608 562294
rect 108224 554963 108252 566510
rect 108316 556374 108344 572154
rect 108396 572076 108448 572082
rect 108396 572018 108448 572024
rect 108408 557462 108436 572018
rect 108960 571402 108988 575076
rect 110524 575062 111550 575090
rect 114664 575062 114770 575090
rect 110420 572076 110472 572082
rect 110420 572018 110472 572024
rect 108948 571396 109000 571402
rect 108948 571338 109000 571344
rect 109684 565208 109736 565214
rect 109684 565150 109736 565156
rect 108396 557456 108448 557462
rect 108396 557398 108448 557404
rect 108948 556776 109000 556782
rect 108948 556718 109000 556724
rect 108304 556368 108356 556374
rect 108304 556310 108356 556316
rect 108960 554963 108988 556718
rect 109696 554963 109724 565150
rect 110432 554963 110460 572018
rect 110524 562222 110552 575062
rect 112536 573708 112588 573714
rect 112536 573650 112588 573656
rect 110512 562216 110564 562222
rect 110512 562158 110564 562164
rect 111064 559564 111116 559570
rect 111064 559506 111116 559512
rect 111076 554963 111104 559506
rect 111800 556368 111852 556374
rect 111800 556310 111852 556316
rect 111812 554963 111840 556310
rect 112548 554963 112576 573650
rect 113272 571668 113324 571674
rect 113272 571610 113324 571616
rect 113284 554963 113312 571610
rect 114664 561066 114692 575062
rect 115480 572280 115532 572286
rect 115480 572222 115532 572228
rect 114744 569356 114796 569362
rect 114744 569298 114796 569304
rect 114652 561060 114704 561066
rect 114652 561002 114704 561008
rect 114756 557534 114784 569298
rect 114756 557506 115428 557534
rect 114652 557456 114704 557462
rect 114652 557398 114704 557404
rect 114008 557184 114060 557190
rect 114008 557126 114060 557132
rect 114020 554963 114048 557126
rect 114664 554963 114692 557398
rect 115400 554963 115428 557506
rect 115492 556238 115520 572222
rect 117332 572014 117360 575076
rect 119712 572144 119764 572150
rect 119712 572086 119764 572092
rect 117320 572008 117372 572014
rect 117320 571950 117372 571956
rect 116584 571396 116636 571402
rect 116584 571338 116636 571344
rect 116596 559638 116624 571338
rect 116584 559632 116636 559638
rect 116584 559574 116636 559580
rect 116860 557116 116912 557122
rect 116860 557058 116912 557064
rect 118240 557116 118292 557122
rect 118240 557058 118292 557064
rect 115480 556232 115532 556238
rect 115480 556174 115532 556180
rect 116124 556232 116176 556238
rect 116124 556174 116176 556180
rect 116136 554963 116164 556174
rect 116872 554963 116900 557058
rect 117596 556980 117648 556986
rect 117596 556922 117648 556928
rect 117608 554963 117636 556922
rect 118252 554963 118280 557058
rect 118976 556980 119028 556986
rect 118976 556922 119028 556928
rect 118988 554963 119016 556922
rect 119724 554963 119752 572086
rect 120552 571402 120580 575076
rect 120736 572082 120764 637350
rect 120724 572076 120776 572082
rect 120724 572018 120776 572024
rect 120540 571396 120592 571402
rect 120540 571338 120592 571344
rect 120448 559564 120500 559570
rect 120448 559506 120500 559512
rect 120460 554963 120488 559506
rect 120828 556850 120856 640358
rect 120908 637628 120960 637634
rect 120908 637570 120960 637576
rect 120920 573646 120948 637570
rect 120998 597680 121054 597689
rect 120998 597615 121054 597624
rect 120908 573640 120960 573646
rect 120908 573582 120960 573588
rect 121012 563854 121040 597615
rect 121090 579864 121146 579873
rect 121090 579799 121146 579808
rect 121104 571674 121132 579799
rect 121182 577144 121238 577153
rect 121182 577079 121238 577088
rect 121092 571668 121144 571674
rect 121092 571610 121144 571616
rect 121000 563848 121052 563854
rect 121000 563790 121052 563796
rect 121196 563718 121224 577079
rect 121472 573578 121500 640426
rect 121644 637696 121696 637702
rect 121644 637638 121696 637644
rect 121550 589384 121606 589393
rect 121550 589319 121606 589328
rect 121564 575074 121592 589319
rect 121552 575068 121604 575074
rect 121552 575010 121604 575016
rect 121460 573572 121512 573578
rect 121460 573514 121512 573520
rect 121184 563712 121236 563718
rect 121184 563654 121236 563660
rect 121552 563712 121604 563718
rect 121552 563654 121604 563660
rect 120816 556844 120868 556850
rect 120816 556786 120868 556792
rect 121092 556232 121144 556238
rect 121092 556174 121144 556180
rect 121564 556186 121592 563654
rect 121656 557054 121684 637638
rect 122194 628824 122250 628833
rect 122194 628759 122250 628768
rect 121826 626104 121882 626113
rect 121826 626039 121882 626048
rect 121734 622704 121790 622713
rect 121734 622639 121790 622648
rect 121748 560998 121776 622639
rect 121840 573442 121868 626039
rect 121918 619984 121974 619993
rect 121918 619919 121974 619928
rect 121828 573436 121880 573442
rect 121828 573378 121880 573384
rect 121932 570722 121960 619919
rect 122010 613864 122066 613873
rect 122010 613799 122066 613808
rect 121920 570716 121972 570722
rect 121920 570658 121972 570664
rect 122024 565146 122052 613799
rect 122102 595504 122158 595513
rect 122102 595439 122158 595448
rect 122116 566710 122144 595439
rect 122104 566704 122156 566710
rect 122104 566646 122156 566652
rect 122012 565140 122064 565146
rect 122012 565082 122064 565088
rect 122104 565140 122156 565146
rect 122104 565082 122156 565088
rect 121736 560992 121788 560998
rect 121736 560934 121788 560940
rect 121644 557048 121696 557054
rect 121644 556990 121696 556996
rect 122116 556238 122144 565082
rect 122208 562494 122236 628759
rect 122286 585984 122342 585993
rect 122286 585919 122342 585928
rect 122300 573510 122328 585919
rect 122852 575006 122880 640494
rect 124220 640416 124272 640422
rect 124220 640358 124272 640364
rect 122930 634944 122986 634953
rect 122930 634879 122986 634888
rect 122840 575000 122892 575006
rect 122840 574942 122892 574948
rect 122288 573504 122340 573510
rect 122288 573446 122340 573452
rect 122944 573374 122972 634879
rect 123022 632224 123078 632233
rect 123022 632159 123078 632168
rect 123036 573714 123064 632159
rect 123206 616584 123262 616593
rect 123206 616519 123262 616528
rect 123114 610464 123170 610473
rect 123114 610399 123170 610408
rect 123024 573708 123076 573714
rect 123024 573650 123076 573656
rect 122932 573368 122984 573374
rect 122932 573310 122984 573316
rect 122840 570784 122892 570790
rect 122840 570726 122892 570732
rect 122564 566568 122616 566574
rect 122564 566510 122616 566516
rect 122196 562488 122248 562494
rect 122196 562430 122248 562436
rect 122104 556232 122156 556238
rect 121104 554963 121132 556174
rect 121564 556158 121868 556186
rect 122104 556174 122156 556180
rect 121840 554963 121868 556158
rect 122576 554963 122604 566510
rect 122852 557534 122880 570726
rect 123128 558210 123156 610399
rect 123220 567866 123248 616519
rect 123298 607744 123354 607753
rect 123298 607679 123354 607688
rect 123312 570858 123340 607679
rect 124126 604344 124182 604353
rect 124126 604279 124182 604288
rect 124140 603158 124168 604279
rect 124128 603152 124180 603158
rect 124128 603094 124180 603100
rect 123390 601624 123446 601633
rect 123390 601559 123446 601568
rect 123300 570852 123352 570858
rect 123300 570794 123352 570800
rect 123208 567860 123260 567866
rect 123208 567802 123260 567808
rect 123404 566506 123432 601559
rect 123482 592104 123538 592113
rect 123482 592039 123538 592048
rect 123496 569294 123524 592039
rect 123574 583264 123630 583273
rect 123574 583199 123630 583208
rect 123588 574802 123616 583199
rect 123576 574796 123628 574802
rect 123576 574738 123628 574744
rect 123484 569288 123536 569294
rect 123484 569230 123536 569236
rect 123392 566500 123444 566506
rect 123392 566442 123444 566448
rect 124232 562358 124260 640358
rect 124312 638988 124364 638994
rect 124312 638930 124364 638936
rect 124220 562352 124272 562358
rect 124220 562294 124272 562300
rect 124036 560992 124088 560998
rect 124036 560934 124088 560940
rect 123116 558204 123168 558210
rect 123116 558146 123168 558152
rect 122852 557506 123340 557534
rect 123312 554963 123340 557506
rect 124048 554963 124076 560934
rect 124324 557190 124352 638930
rect 124404 637764 124456 637770
rect 124404 637706 124456 637712
rect 124312 557184 124364 557190
rect 124312 557126 124364 557132
rect 124416 556918 124444 637706
rect 124508 574870 124536 640698
rect 124588 640688 124640 640694
rect 124588 640630 124640 640636
rect 124600 575142 124628 640630
rect 124680 640620 124732 640626
rect 124680 640562 124732 640568
rect 124588 575136 124640 575142
rect 124588 575078 124640 575084
rect 124692 574938 124720 640562
rect 133880 640348 133932 640354
rect 133880 640290 133932 640296
rect 133144 639056 133196 639062
rect 133144 638998 133196 639004
rect 126244 638036 126296 638042
rect 126244 637978 126296 637984
rect 125600 592068 125652 592074
rect 125600 592010 125652 592016
rect 124680 574932 124732 574938
rect 124680 574874 124732 574880
rect 124496 574864 124548 574870
rect 124496 574806 124548 574812
rect 125612 562358 125640 592010
rect 126152 573572 126204 573578
rect 126152 573514 126204 573520
rect 125416 562352 125468 562358
rect 125416 562294 125468 562300
rect 125600 562352 125652 562358
rect 125600 562294 125652 562300
rect 124680 559632 124732 559638
rect 124680 559574 124732 559580
rect 124404 556912 124456 556918
rect 124404 556854 124456 556860
rect 124692 554963 124720 559574
rect 125428 554963 125456 562294
rect 126164 554963 126192 573514
rect 126256 557122 126284 637978
rect 132500 622464 132552 622470
rect 132500 622406 132552 622412
rect 130384 589348 130436 589354
rect 130384 589290 130436 589296
rect 129740 574932 129792 574938
rect 129740 574874 129792 574880
rect 129004 573640 129056 573646
rect 129004 573582 129056 573588
rect 127624 562420 127676 562426
rect 127624 562362 127676 562368
rect 126888 562352 126940 562358
rect 126888 562294 126940 562300
rect 126244 557116 126296 557122
rect 126244 557058 126296 557064
rect 126900 554963 126928 562294
rect 127636 554963 127664 562362
rect 128268 558204 128320 558210
rect 128268 558146 128320 558152
rect 128280 554963 128308 558146
rect 129016 554963 129044 573582
rect 129752 554963 129780 574874
rect 129832 572212 129884 572218
rect 129832 572154 129884 572160
rect 129844 557534 129872 572154
rect 130396 559570 130424 589290
rect 130384 559564 130436 559570
rect 130384 559506 130436 559512
rect 131212 558272 131264 558278
rect 131212 558214 131264 558220
rect 129844 557506 130516 557534
rect 130488 554963 130516 557506
rect 131224 554963 131252 558214
rect 132512 557534 132540 622406
rect 132684 572008 132736 572014
rect 132684 571950 132736 571956
rect 131856 557524 131908 557530
rect 132512 557506 132632 557534
rect 131856 557466 131908 557472
rect 131868 554963 131896 557466
rect 132604 554963 132632 557506
rect 132696 556186 132724 571950
rect 133156 557530 133184 638998
rect 133892 557534 133920 640290
rect 134524 604512 134576 604518
rect 134524 604454 134576 604460
rect 134156 572076 134208 572082
rect 134156 572018 134208 572024
rect 133144 557524 133196 557530
rect 133892 557506 134104 557534
rect 133144 557466 133196 557472
rect 132696 556158 133368 556186
rect 133340 554963 133368 556158
rect 134076 554963 134104 557506
rect 134168 556186 134196 572018
rect 134536 556986 134564 604454
rect 134616 603152 134668 603158
rect 134616 603094 134668 603100
rect 134628 575414 134656 603094
rect 134616 575408 134668 575414
rect 134616 575350 134668 575356
rect 134904 574802 134932 640766
rect 134984 640620 135036 640626
rect 134984 640562 135036 640568
rect 134996 574870 135024 640562
rect 135260 638988 135312 638994
rect 135260 638930 135312 638936
rect 135168 637968 135220 637974
rect 135168 637910 135220 637916
rect 135076 637832 135128 637838
rect 135076 637774 135128 637780
rect 134984 574864 135036 574870
rect 134984 574806 135036 574812
rect 134892 574796 134944 574802
rect 134892 574738 134944 574744
rect 135088 557122 135116 637774
rect 135180 557190 135208 637910
rect 135272 564942 135300 638930
rect 136456 637900 136508 637906
rect 136456 637842 136508 637848
rect 135352 618248 135404 618254
rect 135352 618190 135404 618196
rect 135364 576854 135392 618190
rect 135364 576826 135484 576854
rect 135260 564936 135312 564942
rect 135260 564878 135312 564884
rect 135168 557184 135220 557190
rect 135168 557126 135220 557132
rect 135076 557116 135128 557122
rect 135076 557058 135128 557064
rect 134524 556980 134576 556986
rect 134524 556922 134576 556928
rect 134168 556158 134748 556186
rect 134720 554963 134748 556158
rect 135456 554963 135484 576826
rect 136180 564936 136232 564942
rect 136180 564878 136232 564884
rect 136192 554963 136220 564878
rect 136468 556918 136496 637842
rect 136560 557054 136588 640834
rect 137282 635624 137338 635633
rect 137282 635559 137338 635568
rect 136638 623384 136694 623393
rect 136638 623319 136694 623328
rect 136652 622470 136680 623319
rect 136640 622464 136692 622470
rect 136640 622406 136692 622412
rect 137098 620664 137154 620673
rect 137098 620599 137154 620608
rect 137006 617264 137062 617273
rect 137006 617199 137062 617208
rect 136638 592784 136694 592793
rect 136638 592719 136694 592728
rect 136652 592074 136680 592719
rect 136640 592068 136692 592074
rect 136640 592010 136692 592016
rect 136638 590064 136694 590073
rect 136638 589999 136694 590008
rect 136652 589354 136680 589999
rect 136640 589348 136692 589354
rect 136640 589290 136692 589296
rect 137020 573374 137048 617199
rect 137008 573368 137060 573374
rect 137008 573310 137060 573316
rect 137112 567866 137140 620599
rect 137296 618254 137324 635559
rect 137284 618248 137336 618254
rect 137284 618190 137336 618196
rect 137572 614553 137600 658242
rect 191852 649330 191880 683086
rect 291200 650072 291252 650078
rect 291200 650014 291252 650020
rect 191840 649324 191892 649330
rect 191840 649266 191892 649272
rect 280988 648780 281040 648786
rect 280988 648722 281040 648728
rect 217784 648644 217836 648650
rect 217784 648586 217836 648592
rect 149060 640892 149112 640898
rect 149060 640834 149112 640840
rect 140320 640824 140372 640830
rect 140320 640766 140372 640772
rect 139860 640756 139912 640762
rect 139860 640698 139912 640704
rect 137836 640688 137888 640694
rect 137836 640630 137888 640636
rect 137652 640484 137704 640490
rect 137652 640426 137704 640432
rect 137558 614544 137614 614553
rect 137558 614479 137614 614488
rect 137282 611144 137338 611153
rect 137282 611079 137338 611088
rect 137296 576230 137324 611079
rect 137374 605024 137430 605033
rect 137374 604959 137430 604968
rect 137388 604518 137416 604959
rect 137376 604512 137428 604518
rect 137376 604454 137428 604460
rect 137374 602304 137430 602313
rect 137374 602239 137430 602248
rect 137284 576224 137336 576230
rect 137284 576166 137336 576172
rect 137388 575550 137416 602239
rect 137466 596184 137522 596193
rect 137466 596119 137522 596128
rect 137376 575544 137428 575550
rect 137376 575486 137428 575492
rect 137100 567860 137152 567866
rect 137100 567802 137152 567808
rect 137480 562290 137508 596119
rect 137664 575142 137692 640426
rect 137742 629504 137798 629513
rect 137742 629439 137798 629448
rect 137652 575136 137704 575142
rect 137652 575078 137704 575084
rect 137468 562284 137520 562290
rect 137468 562226 137520 562232
rect 136916 559700 136968 559706
rect 136916 559642 136968 559648
rect 136548 557048 136600 557054
rect 136548 556990 136600 556996
rect 136456 556912 136508 556918
rect 136456 556854 136508 556860
rect 136928 554963 136956 559642
rect 137756 556986 137784 629439
rect 137848 557326 137876 640630
rect 139216 640552 139268 640558
rect 139216 640494 139268 640500
rect 138664 637764 138716 637770
rect 138664 637706 138716 637712
rect 137928 637628 137980 637634
rect 137928 637570 137980 637576
rect 137940 611153 137968 637570
rect 137926 611144 137982 611153
rect 137926 611079 137982 611088
rect 137926 583944 137982 583953
rect 137926 583879 137982 583888
rect 137940 570722 137968 583879
rect 138570 580544 138626 580553
rect 138570 580479 138626 580488
rect 138478 577824 138534 577833
rect 138478 577759 138534 577768
rect 137928 570716 137980 570722
rect 137928 570658 137980 570664
rect 138296 569424 138348 569430
rect 138296 569366 138348 569372
rect 137836 557320 137888 557326
rect 137836 557262 137888 557268
rect 137744 556980 137796 556986
rect 137744 556922 137796 556928
rect 137652 556300 137704 556306
rect 137652 556242 137704 556248
rect 137664 554963 137692 556242
rect 138308 554963 138336 569366
rect 138492 569294 138520 577759
rect 138480 569288 138532 569294
rect 138480 569230 138532 569236
rect 138584 566506 138612 580479
rect 138572 566500 138624 566506
rect 138572 566442 138624 566448
rect 138480 562488 138532 562494
rect 138480 562430 138532 562436
rect 138492 556186 138520 562430
rect 138676 556306 138704 637706
rect 138756 637696 138808 637702
rect 138756 637638 138808 637644
rect 138768 557394 138796 637638
rect 139122 632904 139178 632913
rect 139122 632839 139178 632848
rect 139030 626784 139086 626793
rect 139030 626719 139086 626728
rect 138938 608424 138994 608433
rect 138938 608359 138994 608368
rect 138846 598904 138902 598913
rect 138846 598839 138902 598848
rect 138860 575006 138888 598839
rect 138848 575000 138900 575006
rect 138848 574942 138900 574948
rect 138952 558346 138980 608359
rect 139044 574258 139072 626719
rect 139032 574252 139084 574258
rect 139032 574194 139084 574200
rect 139136 573442 139164 632839
rect 139228 575278 139256 640494
rect 139306 586664 139362 586673
rect 139306 586599 139362 586608
rect 139320 576854 139348 586599
rect 139320 576826 139440 576854
rect 139216 575272 139268 575278
rect 139216 575214 139268 575220
rect 139124 573436 139176 573442
rect 139124 573378 139176 573384
rect 138940 558340 138992 558346
rect 138940 558282 138992 558288
rect 139412 557534 139440 576826
rect 139872 575210 139900 640698
rect 140332 640626 140360 640766
rect 140228 640620 140280 640626
rect 140228 640562 140280 640568
rect 140320 640620 140372 640626
rect 140320 640562 140372 640568
rect 140240 640490 140268 640562
rect 140136 640484 140188 640490
rect 140136 640426 140188 640432
rect 140228 640484 140280 640490
rect 140228 640426 140280 640432
rect 140148 640354 140176 640426
rect 140044 640348 140096 640354
rect 140044 640290 140096 640296
rect 140136 640348 140188 640354
rect 140136 640290 140188 640296
rect 140056 638044 140084 640290
rect 149072 638044 149100 640834
rect 213920 640824 213972 640830
rect 213920 640766 213972 640772
rect 157432 640756 157484 640762
rect 157432 640698 157484 640704
rect 212540 640756 212592 640762
rect 212540 640698 212592 640704
rect 151636 639056 151688 639062
rect 151636 638998 151688 639004
rect 151648 638044 151676 638998
rect 157444 638044 157472 640698
rect 160652 640688 160704 640694
rect 160652 640630 160704 640636
rect 160664 638044 160692 640630
rect 166448 640620 166500 640626
rect 166448 640562 166500 640568
rect 166460 638044 166488 640562
rect 174820 640552 174872 640558
rect 174820 640494 174872 640500
rect 189632 640552 189684 640558
rect 189632 640494 189684 640500
rect 205640 640552 205692 640558
rect 205640 640494 205692 640500
rect 172244 640416 172296 640422
rect 172244 640358 172296 640364
rect 172256 638044 172284 640358
rect 174832 638044 174860 640494
rect 180616 640484 180668 640490
rect 180616 640426 180668 640432
rect 177868 638042 178066 638058
rect 180628 638044 180656 640426
rect 186412 640348 186464 640354
rect 186412 640290 186464 640296
rect 183836 638988 183888 638994
rect 183836 638930 183888 638936
rect 183848 638044 183876 638930
rect 186424 638044 186452 640290
rect 189644 638044 189672 640494
rect 192208 640416 192260 640422
rect 192208 640358 192260 640364
rect 204352 640416 204404 640422
rect 204352 640358 204404 640364
rect 192220 638044 192248 640358
rect 195428 640348 195480 640354
rect 195428 640290 195480 640296
rect 200856 640348 200908 640354
rect 200856 640290 200908 640296
rect 195440 638044 195468 640290
rect 177856 638036 178066 638042
rect 177908 638030 178066 638036
rect 177856 637978 177908 637984
rect 145564 637968 145616 637974
rect 145616 637916 145866 637922
rect 145564 637910 145866 637916
rect 145576 637894 145866 637910
rect 154592 637906 154882 637922
rect 154580 637900 154882 637906
rect 154632 637894 154882 637900
rect 154580 637842 154632 637848
rect 162860 637832 162912 637838
rect 162912 637780 163254 637786
rect 162860 637774 163254 637780
rect 162872 637758 163254 637774
rect 168760 637770 169050 637786
rect 168748 637764 169050 637770
rect 168800 637758 169050 637764
rect 168748 637706 168800 637712
rect 142988 637696 143040 637702
rect 198280 637696 198332 637702
rect 143040 637644 143290 637650
rect 142988 637638 143290 637644
rect 143000 637622 143290 637638
rect 198030 637644 198280 637650
rect 198030 637638 198332 637644
rect 198030 637622 198320 637638
rect 200606 637350 200712 637378
rect 140136 575544 140188 575550
rect 140136 575486 140188 575492
rect 139860 575204 139912 575210
rect 139860 575146 139912 575152
rect 139504 575062 140070 575090
rect 139504 561066 139532 575062
rect 140148 567194 140176 575486
rect 142160 575272 142212 575278
rect 142160 575214 142212 575220
rect 140780 575204 140832 575210
rect 140780 575146 140832 575152
rect 139872 567166 140176 567194
rect 139492 561060 139544 561066
rect 139492 561002 139544 561008
rect 139412 557506 139808 557534
rect 138756 557388 138808 557394
rect 138756 557330 138808 557336
rect 138664 556300 138716 556306
rect 138664 556242 138716 556248
rect 138492 556158 139072 556186
rect 139044 554963 139072 556158
rect 139780 554963 139808 557506
rect 139872 557258 139900 567166
rect 140792 562358 140820 575146
rect 141240 574252 141292 574258
rect 141240 574194 141292 574200
rect 140780 562352 140832 562358
rect 140780 562294 140832 562300
rect 140504 561128 140556 561134
rect 140504 561070 140556 561076
rect 139860 557252 139912 557258
rect 139860 557194 139912 557200
rect 140516 554963 140544 561070
rect 141252 554963 141280 574194
rect 141884 562352 141936 562358
rect 141884 562294 141936 562300
rect 141896 554963 141924 562294
rect 142172 562222 142200 575214
rect 164332 575204 164384 575210
rect 164332 575146 164384 575152
rect 145472 575136 145524 575142
rect 142264 575062 142646 575090
rect 145472 575078 145524 575084
rect 142264 563786 142292 575062
rect 143540 572416 143592 572422
rect 143540 572358 143592 572364
rect 142620 565208 142672 565214
rect 142620 565150 142672 565156
rect 142252 563780 142304 563786
rect 142252 563722 142304 563728
rect 142160 562216 142212 562222
rect 142160 562158 142212 562164
rect 142632 554963 142660 565150
rect 143552 562290 143580 572358
rect 145208 572150 145236 575076
rect 145196 572144 145248 572150
rect 145196 572086 145248 572092
rect 144092 563916 144144 563922
rect 144092 563858 144144 563864
rect 143540 562284 143592 562290
rect 143540 562226 143592 562232
rect 143356 562216 143408 562222
rect 143356 562158 143408 562164
rect 143368 554963 143396 562158
rect 144104 554963 144132 563858
rect 144736 562284 144788 562290
rect 144736 562226 144788 562232
rect 144748 554963 144776 562226
rect 145484 554963 145512 575078
rect 148428 572490 148456 575076
rect 149152 575000 149204 575006
rect 149152 574942 149204 574948
rect 148416 572484 148468 572490
rect 148416 572426 148468 572432
rect 147680 572348 147732 572354
rect 147680 572290 147732 572296
rect 147692 562290 147720 572290
rect 147772 572144 147824 572150
rect 147772 572086 147824 572092
rect 147680 562284 147732 562290
rect 147680 562226 147732 562232
rect 146944 557388 146996 557394
rect 146944 557330 146996 557336
rect 146208 556844 146260 556850
rect 146208 556786 146260 556792
rect 146220 554963 146248 556786
rect 146956 554963 146984 557330
rect 147784 555234 147812 572086
rect 148324 562284 148376 562290
rect 148324 562226 148376 562232
rect 147708 555206 147812 555234
rect 147708 554948 147736 555206
rect 148336 554963 148364 562226
rect 149164 555234 149192 574942
rect 150624 573436 150676 573442
rect 150624 573378 150676 573384
rect 149796 558340 149848 558346
rect 149796 558282 149848 558288
rect 149088 555206 149192 555234
rect 149088 554948 149116 555206
rect 149808 554963 149836 558282
rect 150636 555234 150664 573378
rect 151004 572558 151032 575076
rect 151912 574864 151964 574870
rect 151912 574806 151964 574812
rect 150992 572552 151044 572558
rect 150992 572494 151044 572500
rect 151268 557320 151320 557326
rect 151268 557262 151320 557268
rect 150560 555206 150664 555234
rect 150560 554948 150588 555206
rect 151280 554963 151308 557262
rect 151924 554963 151952 574806
rect 154224 572218 154252 575076
rect 156236 575068 156288 575074
rect 156236 575010 156288 575016
rect 154580 575000 154632 575006
rect 154580 574942 154632 574948
rect 154212 572212 154264 572218
rect 154212 572154 154264 572160
rect 154592 562290 154620 574942
rect 154856 572280 154908 572286
rect 154856 572222 154908 572228
rect 154580 562284 154632 562290
rect 154580 562226 154632 562232
rect 152648 558340 152700 558346
rect 152648 558282 152700 558288
rect 152660 554963 152688 558282
rect 153384 557252 153436 557258
rect 153384 557194 153436 557200
rect 153396 554963 153424 557194
rect 154120 556232 154172 556238
rect 154120 556174 154172 556180
rect 154132 554963 154160 556174
rect 154868 554963 154896 572222
rect 155500 562284 155552 562290
rect 155500 562226 155552 562232
rect 155512 554963 155540 562226
rect 156248 554963 156276 575010
rect 156800 572422 156828 575076
rect 159364 572484 159416 572490
rect 159364 572426 159416 572432
rect 156788 572416 156840 572422
rect 156788 572358 156840 572364
rect 158720 572212 158772 572218
rect 158720 572154 158772 572160
rect 157984 566704 158036 566710
rect 157984 566646 158036 566652
rect 156972 557184 157024 557190
rect 156972 557126 157024 557132
rect 156984 554963 157012 557126
rect 157708 556912 157760 556918
rect 157708 556854 157760 556860
rect 157720 554963 157748 556854
rect 157996 556238 158024 566646
rect 158732 563446 158760 572154
rect 159088 569288 159140 569294
rect 159088 569230 159140 569236
rect 158720 563440 158772 563446
rect 158720 563382 158772 563388
rect 158352 556912 158404 556918
rect 158352 556854 158404 556860
rect 157984 556232 158036 556238
rect 157984 556174 158036 556180
rect 158364 554963 158392 556854
rect 159100 554963 159128 569230
rect 159376 557326 159404 572426
rect 160020 572422 160048 575076
rect 161940 574796 161992 574802
rect 161940 574738 161992 574744
rect 160560 573368 160612 573374
rect 160560 573310 160612 573316
rect 160008 572416 160060 572422
rect 160008 572358 160060 572364
rect 159824 563440 159876 563446
rect 159824 563382 159876 563388
rect 159364 557320 159416 557326
rect 159364 557262 159416 557268
rect 159836 554963 159864 563382
rect 160572 554963 160600 573310
rect 160744 572552 160796 572558
rect 160744 572494 160796 572500
rect 160652 566500 160704 566506
rect 160652 566442 160704 566448
rect 160664 556186 160692 566442
rect 160756 557190 160784 572494
rect 160744 557184 160796 557190
rect 160744 557126 160796 557132
rect 160664 556158 161336 556186
rect 161308 554963 161336 556158
rect 161952 554963 161980 574738
rect 162596 572354 162624 575076
rect 162584 572348 162636 572354
rect 162584 572290 162636 572296
rect 164344 562290 164372 575146
rect 183468 575136 183520 575142
rect 164884 572416 164936 572422
rect 164884 572358 164936 572364
rect 164332 562284 164384 562290
rect 164332 562226 164384 562232
rect 163412 561060 163464 561066
rect 163412 561002 163464 561008
rect 162676 556300 162728 556306
rect 162676 556242 162728 556248
rect 162688 554963 162716 556242
rect 163424 554963 163452 561002
rect 164896 557394 164924 572358
rect 165816 571402 165844 575076
rect 165804 571396 165856 571402
rect 165804 571338 165856 571344
rect 167828 571396 167880 571402
rect 167828 571338 167880 571344
rect 166264 567860 166316 567866
rect 166264 567802 166316 567808
rect 165528 562284 165580 562290
rect 165528 562226 165580 562232
rect 164884 557388 164936 557394
rect 164884 557330 164936 557336
rect 164148 557252 164200 557258
rect 164148 557194 164200 557200
rect 164160 554963 164188 557194
rect 164884 557116 164936 557122
rect 164884 557058 164936 557064
rect 164896 554963 164924 557058
rect 165540 554963 165568 562226
rect 166276 554963 166304 567802
rect 167736 563780 167788 563786
rect 167736 563722 167788 563728
rect 167000 557320 167052 557326
rect 167000 557262 167052 557268
rect 167012 554963 167040 557262
rect 167748 554963 167776 563722
rect 167840 556238 167868 571338
rect 168392 556306 168420 575076
rect 171612 572286 171640 575076
rect 171600 572280 171652 572286
rect 171600 572222 171652 572228
rect 174188 571402 174216 575076
rect 177408 572014 177436 575076
rect 179524 575062 179998 575090
rect 183468 575078 183520 575084
rect 179420 574796 179472 574802
rect 179420 574738 179472 574744
rect 177396 572008 177448 572014
rect 177396 571950 177448 571956
rect 171784 571396 171836 571402
rect 171784 571338 171836 571344
rect 174176 571396 174228 571402
rect 174176 571338 174228 571344
rect 168472 570852 168524 570858
rect 168472 570794 168524 570800
rect 168380 556300 168432 556306
rect 168380 556242 168432 556248
rect 167828 556232 167880 556238
rect 167828 556174 167880 556180
rect 168484 555234 168512 570794
rect 169116 570716 169168 570722
rect 169116 570658 169168 570664
rect 168408 555206 168512 555234
rect 168408 554948 168436 555206
rect 169128 554963 169156 570658
rect 170588 567996 170640 568002
rect 170588 567938 170640 567944
rect 169852 556232 169904 556238
rect 169852 556174 169904 556180
rect 169864 554963 169892 556174
rect 170600 554963 170628 567938
rect 171796 557258 171824 571338
rect 177028 565276 177080 565282
rect 177028 565218 177080 565224
rect 173164 562352 173216 562358
rect 173164 562294 173216 562300
rect 171784 557252 171836 557258
rect 171784 557194 171836 557200
rect 172704 557184 172756 557190
rect 172704 557126 172756 557132
rect 171968 557116 172020 557122
rect 171968 557058 172020 557064
rect 171324 557048 171376 557054
rect 171324 556990 171376 556996
rect 171336 554963 171364 556990
rect 171980 554963 172008 557058
rect 172716 554963 172744 557126
rect 173176 556442 173204 562294
rect 173440 557388 173492 557394
rect 173440 557330 173492 557336
rect 173164 556436 173216 556442
rect 173164 556378 173216 556384
rect 173452 554963 173480 557330
rect 176292 557116 176344 557122
rect 176292 557058 176344 557064
rect 175556 556980 175608 556986
rect 175556 556922 175608 556928
rect 174912 556436 174964 556442
rect 174912 556378 174964 556384
rect 174176 556300 174228 556306
rect 174176 556242 174228 556248
rect 174188 554963 174216 556242
rect 174924 554963 174952 556378
rect 175568 554963 175596 556922
rect 176304 554963 176332 557058
rect 177040 554963 177068 565218
rect 177764 563984 177816 563990
rect 177764 563926 177816 563932
rect 177776 554963 177804 563926
rect 178500 561196 178552 561202
rect 178500 561138 178552 561144
rect 178512 554963 178540 561138
rect 179144 559564 179196 559570
rect 179144 559506 179196 559512
rect 179156 554963 179184 559506
rect 179432 556186 179460 574738
rect 179524 556306 179552 575062
rect 182272 573436 182324 573442
rect 182272 573378 182324 573384
rect 180800 573368 180852 573374
rect 180800 573310 180852 573316
rect 180616 570716 180668 570722
rect 180616 570658 180668 570664
rect 179512 556300 179564 556306
rect 179512 556242 179564 556248
rect 179432 556158 179920 556186
rect 179892 554963 179920 556158
rect 180628 554963 180656 570658
rect 180812 562358 180840 573310
rect 181352 569288 181404 569294
rect 181352 569230 181404 569236
rect 180800 562352 180852 562358
rect 180800 562294 180852 562300
rect 181364 554963 181392 569230
rect 181996 562352 182048 562358
rect 181996 562294 182048 562300
rect 182008 554963 182036 562294
rect 182284 557534 182312 573378
rect 183204 572218 183232 575076
rect 183192 572212 183244 572218
rect 183192 572154 183244 572160
rect 182284 557506 182772 557534
rect 182744 554963 182772 557506
rect 183480 554963 183508 575078
rect 185780 572150 185808 575076
rect 186320 573504 186372 573510
rect 186320 573446 186372 573452
rect 185768 572144 185820 572150
rect 185768 572086 185820 572092
rect 184204 571396 184256 571402
rect 184204 571338 184256 571344
rect 183560 567860 183612 567866
rect 183560 567802 183612 567808
rect 183572 557534 183600 567802
rect 184216 558278 184244 571338
rect 185584 562352 185636 562358
rect 185584 562294 185636 562300
rect 184940 559768 184992 559774
rect 184940 559710 184992 559716
rect 184204 558272 184256 558278
rect 184204 558214 184256 558220
rect 183572 557506 184244 557534
rect 184216 554963 184244 557506
rect 184952 554963 184980 559710
rect 185596 554963 185624 562294
rect 186332 554963 186360 573446
rect 188344 572212 188396 572218
rect 188344 572154 188396 572160
rect 187056 567928 187108 567934
rect 187056 567870 187108 567876
rect 187068 554963 187096 567870
rect 188068 566636 188120 566642
rect 188068 566578 188120 566584
rect 187792 557524 187844 557530
rect 187792 557466 187844 557472
rect 187804 554963 187832 557466
rect 188080 556866 188108 566578
rect 188356 557054 188384 572154
rect 189000 571402 189028 575076
rect 190564 575062 191590 575090
rect 194612 575062 194810 575090
rect 190460 572144 190512 572150
rect 190460 572086 190512 572092
rect 188988 571396 189040 571402
rect 188988 571338 189040 571344
rect 189172 563848 189224 563854
rect 189172 563790 189224 563796
rect 188344 557048 188396 557054
rect 188344 556990 188396 556996
rect 188080 556838 188568 556866
rect 188540 554963 188568 556838
rect 189184 554963 189212 563790
rect 189908 562624 189960 562630
rect 189908 562566 189960 562572
rect 189920 554963 189948 562566
rect 190472 560862 190500 572086
rect 190564 565146 190592 575062
rect 192760 572008 192812 572014
rect 192760 571950 192812 571956
rect 190644 565344 190696 565350
rect 190644 565286 190696 565292
rect 190552 565140 190604 565146
rect 190552 565082 190604 565088
rect 190460 560856 190512 560862
rect 190460 560798 190512 560804
rect 190656 554963 190684 565286
rect 192116 561264 192168 561270
rect 192116 561206 192168 561212
rect 191380 560856 191432 560862
rect 191380 560798 191432 560804
rect 191392 554963 191420 560798
rect 192128 554963 192156 561206
rect 192772 554963 192800 571950
rect 193220 570920 193272 570926
rect 193220 570862 193272 570868
rect 193232 559026 193260 570862
rect 193496 568064 193548 568070
rect 193496 568006 193548 568012
rect 193220 559020 193272 559026
rect 193220 558962 193272 558968
rect 193508 554963 193536 568006
rect 194612 562426 194640 575062
rect 197084 574864 197136 574870
rect 197084 574806 197136 574812
rect 195244 569356 195296 569362
rect 195244 569298 195296 569304
rect 194968 566500 195020 566506
rect 194968 566442 195020 566448
rect 194600 562420 194652 562426
rect 194600 562362 194652 562368
rect 194232 559020 194284 559026
rect 194232 558962 194284 558968
rect 194244 554963 194272 558962
rect 194980 554963 195008 566442
rect 195256 557530 195284 569298
rect 196348 565140 196400 565146
rect 196348 565082 196400 565088
rect 195244 557524 195296 557530
rect 195244 557466 195296 557472
rect 195612 556980 195664 556986
rect 195612 556922 195664 556928
rect 195624 554963 195652 556922
rect 196360 554963 196388 565082
rect 197096 554963 197124 574806
rect 197372 572082 197400 575076
rect 200592 572558 200620 575076
rect 198004 572552 198056 572558
rect 198004 572494 198056 572500
rect 200580 572552 200632 572558
rect 200580 572494 200632 572500
rect 197360 572076 197412 572082
rect 197360 572018 197412 572024
rect 197820 564052 197872 564058
rect 197820 563994 197872 564000
rect 197832 554963 197860 563994
rect 198016 561134 198044 572494
rect 200684 570858 200712 637350
rect 200762 613320 200818 613329
rect 200762 613255 200818 613264
rect 200672 570852 200724 570858
rect 200672 570794 200724 570800
rect 200776 569430 200804 613255
rect 200868 575210 200896 640290
rect 204260 638988 204312 638994
rect 204260 638930 204312 638936
rect 201500 637696 201552 637702
rect 201500 637638 201552 637644
rect 201038 592104 201094 592113
rect 201038 592039 201094 592048
rect 200948 575544 201000 575550
rect 200948 575486 201000 575492
rect 200856 575204 200908 575210
rect 200856 575146 200908 575152
rect 200764 569424 200816 569430
rect 200764 569366 200816 569372
rect 200672 563780 200724 563786
rect 200672 563722 200724 563728
rect 199200 562420 199252 562426
rect 199200 562362 199252 562368
rect 198004 561128 198056 561134
rect 198004 561070 198056 561076
rect 198556 561060 198608 561066
rect 198556 561002 198608 561008
rect 198568 554963 198596 561002
rect 199212 554963 199240 562362
rect 199936 557048 199988 557054
rect 199936 556990 199988 556996
rect 199948 554963 199976 556990
rect 200684 554963 200712 563722
rect 200960 556918 200988 575486
rect 201052 558210 201080 592039
rect 201130 583264 201186 583273
rect 201130 583199 201186 583208
rect 201144 563718 201172 583199
rect 201222 577144 201278 577153
rect 201222 577079 201278 577088
rect 201132 563712 201184 563718
rect 201132 563654 201184 563660
rect 201236 559638 201264 577079
rect 201224 559632 201276 559638
rect 201224 559574 201276 559580
rect 201040 558204 201092 558210
rect 201040 558146 201092 558152
rect 200948 556912 201000 556918
rect 200948 556854 201000 556860
rect 201512 556850 201540 637638
rect 201590 634944 201646 634953
rect 201590 634879 201646 634888
rect 201604 566574 201632 634879
rect 201774 632224 201830 632233
rect 201774 632159 201830 632168
rect 201682 628824 201738 628833
rect 201682 628759 201738 628768
rect 201592 566568 201644 566574
rect 201592 566510 201644 566516
rect 201696 563922 201724 628759
rect 201788 568002 201816 632159
rect 201958 626104 202014 626113
rect 201958 626039 202014 626048
rect 201866 619984 201922 619993
rect 201866 619919 201922 619928
rect 201776 567996 201828 568002
rect 201776 567938 201828 567944
rect 201684 563916 201736 563922
rect 201684 563858 201736 563864
rect 201880 560998 201908 619919
rect 201972 573578 202000 626039
rect 202970 622704 203026 622713
rect 202970 622639 203026 622648
rect 202878 607744 202934 607753
rect 202878 607679 202934 607688
rect 202142 601624 202198 601633
rect 202142 601559 202198 601568
rect 202050 595504 202106 595513
rect 202050 595439 202106 595448
rect 201960 573572 202012 573578
rect 201960 573514 202012 573520
rect 202064 565214 202092 595439
rect 202156 570790 202184 601559
rect 202234 585984 202290 585993
rect 202234 585919 202290 585928
rect 202144 570784 202196 570790
rect 202144 570726 202196 570732
rect 202052 565208 202104 565214
rect 202052 565150 202104 565156
rect 201868 560992 201920 560998
rect 201868 560934 201920 560940
rect 202248 559706 202276 585919
rect 202236 559700 202288 559706
rect 202236 559642 202288 559648
rect 202144 559632 202196 559638
rect 202144 559574 202196 559580
rect 201500 556844 201552 556850
rect 201500 556786 201552 556792
rect 201408 556300 201460 556306
rect 201408 556242 201460 556248
rect 201420 554963 201448 556242
rect 202156 554963 202184 559574
rect 202892 558346 202920 607679
rect 202984 574938 203012 622639
rect 203154 616584 203210 616593
rect 203154 616519 203210 616528
rect 203062 610464 203118 610473
rect 203062 610399 203118 610408
rect 202972 574932 203024 574938
rect 202972 574874 203024 574880
rect 203076 566710 203104 610399
rect 203168 573646 203196 616519
rect 203890 604344 203946 604353
rect 203890 604279 203946 604288
rect 203904 603158 203932 604279
rect 203892 603152 203944 603158
rect 203892 603094 203944 603100
rect 203246 598224 203302 598233
rect 203246 598159 203302 598168
rect 203156 573640 203208 573646
rect 203156 573582 203208 573588
rect 203064 566704 203116 566710
rect 203064 566646 203116 566652
rect 203260 562494 203288 598159
rect 203338 589384 203394 589393
rect 203338 589319 203394 589328
rect 203352 575550 203380 589319
rect 203430 579864 203486 579873
rect 203430 579799 203486 579808
rect 203340 575544 203392 575550
rect 203340 575486 203392 575492
rect 203444 572218 203472 579799
rect 203432 572212 203484 572218
rect 203432 572154 203484 572160
rect 203248 562488 203300 562494
rect 203248 562430 203300 562436
rect 202880 558340 202932 558346
rect 202880 558282 202932 558288
rect 202788 556368 202840 556374
rect 202788 556310 202840 556316
rect 202800 554963 202828 556310
rect 203524 556232 203576 556238
rect 203524 556174 203576 556180
rect 203536 554963 203564 556174
rect 204272 554963 204300 638930
rect 204364 575006 204392 640358
rect 204904 638036 204956 638042
rect 204904 637978 204956 637984
rect 204352 575000 204404 575006
rect 204352 574942 204404 574948
rect 204916 556238 204944 637978
rect 204996 622464 205048 622470
rect 204996 622406 205048 622412
rect 205008 565350 205036 622406
rect 205652 575074 205680 640494
rect 210424 639124 210476 639130
rect 210424 639066 210476 639072
rect 206284 639056 206336 639062
rect 206284 638998 206336 639004
rect 205640 575068 205692 575074
rect 205640 575010 205692 575016
rect 204996 565344 205048 565350
rect 204996 565286 205048 565292
rect 205732 562556 205784 562562
rect 205732 562498 205784 562504
rect 204996 556844 205048 556850
rect 204996 556786 205048 556792
rect 204904 556232 204956 556238
rect 204904 556174 204956 556180
rect 205008 554963 205036 556786
rect 205744 555234 205772 562498
rect 206296 556306 206324 638998
rect 208400 637900 208452 637906
rect 208400 637842 208452 637848
rect 206376 637832 206428 637838
rect 206376 637774 206428 637780
rect 206388 567194 206416 637774
rect 206468 634840 206520 634846
rect 206468 634782 206520 634788
rect 206480 568070 206508 634782
rect 207020 577516 207072 577522
rect 207020 577458 207072 577464
rect 207032 576854 207060 577458
rect 207032 576826 207888 576854
rect 206468 568064 206520 568070
rect 206468 568006 206520 568012
rect 206388 567166 206508 567194
rect 206376 565208 206428 565214
rect 206376 565150 206428 565156
rect 206284 556300 206336 556306
rect 206284 556242 206336 556248
rect 205668 555206 205772 555234
rect 205668 554948 205696 555206
rect 206388 554963 206416 565150
rect 206480 556986 206508 567166
rect 207112 560992 207164 560998
rect 207112 560934 207164 560940
rect 206468 556980 206520 556986
rect 206468 556922 206520 556928
rect 207124 554963 207152 560934
rect 207860 554963 207888 576826
rect 208412 562290 208440 637842
rect 208492 632120 208544 632126
rect 208492 632062 208544 632068
rect 208504 576854 208532 632062
rect 209044 589348 209096 589354
rect 209044 589290 209096 589296
rect 208504 576826 208624 576854
rect 208400 562284 208452 562290
rect 208400 562226 208452 562232
rect 208596 554963 208624 576826
rect 209056 561202 209084 589290
rect 209228 562284 209280 562290
rect 209228 562226 209280 562232
rect 209044 561196 209096 561202
rect 209044 561138 209096 561144
rect 209136 561128 209188 561134
rect 209136 561070 209188 561076
rect 209148 556374 209176 561070
rect 209136 556368 209188 556374
rect 209136 556310 209188 556316
rect 209240 554963 209268 562226
rect 210436 557054 210464 639066
rect 210516 637764 210568 637770
rect 210516 637706 210568 637712
rect 210528 557122 210556 637706
rect 211804 626612 211856 626618
rect 211804 626554 211856 626560
rect 211160 601724 211212 601730
rect 211160 601666 211212 601672
rect 210608 592068 210660 592074
rect 210608 592010 210660 592016
rect 210620 559774 210648 592010
rect 210700 586560 210752 586566
rect 210700 586502 210752 586508
rect 210712 564058 210740 586502
rect 211172 576854 211200 601666
rect 211172 576826 211476 576854
rect 210700 564052 210752 564058
rect 210700 563994 210752 564000
rect 210608 559768 210660 559774
rect 210608 559710 210660 559716
rect 210700 559700 210752 559706
rect 210700 559642 210752 559648
rect 210516 557116 210568 557122
rect 210516 557058 210568 557064
rect 210424 557048 210476 557054
rect 210424 556990 210476 556996
rect 209964 556300 210016 556306
rect 209964 556242 210016 556248
rect 209976 554963 210004 556242
rect 210712 554963 210740 559642
rect 211448 554963 211476 576826
rect 211816 562426 211844 626554
rect 212552 576854 212580 640698
rect 213184 637968 213236 637974
rect 213184 637910 213236 637916
rect 212552 576826 212948 576854
rect 212172 562488 212224 562494
rect 212172 562430 212224 562436
rect 211804 562420 211856 562426
rect 211804 562362 211856 562368
rect 212184 554963 212212 562430
rect 212816 558000 212868 558006
rect 212816 557942 212868 557948
rect 212828 554963 212856 557942
rect 212920 556186 212948 576826
rect 213196 556850 213224 637910
rect 213276 604512 213328 604518
rect 213276 604454 213328 604460
rect 213288 565282 213316 604454
rect 213932 566574 213960 640766
rect 214012 640484 214064 640490
rect 214012 640426 214064 640432
rect 214024 576854 214052 640426
rect 217324 640348 217376 640354
rect 217324 640290 217376 640296
rect 215300 639260 215352 639266
rect 215300 639202 215352 639208
rect 214564 597576 214616 597582
rect 214564 597518 214616 597524
rect 214024 576826 214328 576854
rect 213920 566568 213972 566574
rect 213920 566510 213972 566516
rect 213276 565276 213328 565282
rect 213276 565218 213328 565224
rect 213184 556844 213236 556850
rect 213184 556786 213236 556792
rect 212920 556158 213592 556186
rect 213564 554963 213592 556158
rect 214300 554963 214328 576826
rect 214576 560998 214604 597518
rect 215024 566568 215076 566574
rect 215024 566510 215076 566516
rect 214564 560992 214616 560998
rect 214564 560934 214616 560940
rect 215036 554963 215064 566510
rect 215312 557534 215340 639202
rect 215944 638172 215996 638178
rect 215944 638114 215996 638120
rect 215852 570784 215904 570790
rect 215852 570726 215904 570732
rect 215312 557506 215800 557534
rect 215772 554963 215800 557506
rect 215864 556186 215892 570726
rect 215956 556306 215984 638114
rect 216036 637696 216088 637702
rect 216036 637638 216088 637644
rect 216048 561270 216076 637638
rect 216678 635624 216734 635633
rect 216678 635559 216734 635568
rect 216692 634846 216720 635559
rect 216680 634840 216732 634846
rect 216680 634782 216732 634788
rect 216678 632904 216734 632913
rect 216678 632839 216734 632848
rect 216692 632126 216720 632839
rect 216680 632120 216732 632126
rect 216680 632062 216732 632068
rect 216678 626784 216734 626793
rect 216678 626719 216734 626728
rect 216692 626618 216720 626719
rect 216680 626612 216732 626618
rect 216680 626554 216732 626560
rect 216678 623384 216734 623393
rect 216678 623319 216734 623328
rect 216692 622470 216720 623319
rect 216680 622464 216732 622470
rect 216680 622406 216732 622412
rect 216678 605024 216734 605033
rect 216678 604959 216734 604968
rect 216692 604518 216720 604959
rect 216680 604512 216732 604518
rect 216680 604454 216732 604460
rect 216772 603152 216824 603158
rect 216772 603094 216824 603100
rect 216678 602304 216734 602313
rect 216678 602239 216734 602248
rect 216692 601730 216720 602239
rect 216680 601724 216732 601730
rect 216680 601666 216732 601672
rect 216678 592784 216734 592793
rect 216678 592719 216734 592728
rect 216692 592074 216720 592719
rect 216680 592068 216732 592074
rect 216680 592010 216732 592016
rect 216678 590064 216734 590073
rect 216678 589999 216734 590008
rect 216692 589354 216720 589999
rect 216680 589348 216732 589354
rect 216680 589290 216732 589296
rect 216678 586664 216734 586673
rect 216678 586599 216734 586608
rect 216692 586566 216720 586599
rect 216680 586560 216732 586566
rect 216680 586502 216732 586508
rect 216678 577824 216734 577833
rect 216678 577759 216734 577768
rect 216692 567194 216720 577759
rect 216784 575414 216812 603094
rect 217046 598904 217102 598913
rect 217046 598839 217102 598848
rect 217060 597582 217088 598839
rect 217048 597576 217100 597582
rect 217048 597518 217100 597524
rect 216772 575408 216824 575414
rect 216772 575350 216824 575356
rect 216692 567166 217180 567194
rect 216036 561264 216088 561270
rect 216036 561206 216088 561212
rect 215944 556300 215996 556306
rect 215944 556242 215996 556248
rect 215864 556158 216444 556186
rect 216416 554963 216444 556158
rect 217152 554963 217180 567166
rect 217336 562630 217364 640290
rect 217690 629504 217746 629513
rect 217690 629439 217746 629448
rect 217598 617264 217654 617273
rect 217598 617199 217654 617208
rect 217414 608424 217470 608433
rect 217414 608359 217470 608368
rect 217428 577522 217456 608359
rect 217416 577516 217468 577522
rect 217416 577458 217468 577464
rect 217324 562624 217376 562630
rect 217324 562566 217376 562572
rect 217612 557569 217640 617199
rect 217704 596018 217732 629439
rect 217796 614553 217824 648586
rect 280712 646672 280764 646678
rect 280712 646614 280764 646620
rect 218704 645924 218756 645930
rect 218704 645866 218756 645872
rect 217876 640688 217928 640694
rect 217876 640630 217928 640636
rect 217782 614544 217838 614553
rect 217782 614479 217838 614488
rect 217782 596184 217838 596193
rect 217782 596119 217838 596128
rect 217692 596012 217744 596018
rect 217692 595954 217744 595960
rect 217796 586514 217824 596119
rect 217704 586486 217824 586514
rect 217704 576230 217732 586486
rect 217692 576224 217744 576230
rect 217692 576166 217744 576172
rect 217888 574938 217916 640630
rect 217968 638104 218020 638110
rect 217968 638046 218020 638052
rect 217876 574932 217928 574938
rect 217876 574874 217928 574880
rect 217876 561196 217928 561202
rect 217876 561138 217928 561144
rect 217598 557560 217654 557569
rect 217598 557495 217654 557504
rect 217888 554963 217916 561138
rect 217980 557648 218008 638046
rect 218716 637634 218744 645866
rect 225788 640824 225840 640830
rect 225788 640766 225840 640772
rect 218888 640620 218940 640626
rect 218888 640562 218940 640568
rect 218796 640552 218848 640558
rect 218796 640494 218848 640500
rect 218704 637628 218756 637634
rect 218704 637570 218756 637576
rect 218716 611153 218744 637570
rect 218702 611144 218758 611153
rect 218702 611079 218758 611088
rect 218704 596012 218756 596018
rect 218704 595954 218756 595960
rect 218150 580544 218206 580553
rect 218150 580479 218206 580488
rect 218164 562426 218192 580479
rect 218152 562420 218204 562426
rect 218152 562362 218204 562368
rect 217980 557620 218100 557648
rect 217966 557560 218022 557569
rect 217966 557495 218022 557504
rect 217980 557054 218008 557495
rect 217968 557048 218020 557054
rect 217968 556990 218020 556996
rect 218072 556986 218100 557620
rect 218612 557048 218664 557054
rect 218612 556990 218664 556996
rect 218060 556980 218112 556986
rect 218060 556922 218112 556928
rect 218624 554963 218652 556990
rect 218716 556850 218744 595954
rect 218808 570926 218836 640494
rect 218900 575142 218928 640562
rect 219348 640416 219400 640422
rect 219348 640358 219400 640364
rect 219254 620664 219310 620673
rect 219254 620599 219310 620608
rect 219162 583944 219218 583953
rect 219162 583879 219218 583888
rect 218888 575136 218940 575142
rect 218888 575078 218940 575084
rect 218796 570920 218848 570926
rect 218796 570862 218848 570868
rect 219176 558278 219204 583879
rect 219268 573578 219296 620599
rect 219360 575006 219388 640358
rect 219624 639192 219676 639198
rect 219624 639134 219676 639140
rect 219348 575000 219400 575006
rect 219348 574942 219400 574948
rect 219256 573572 219308 573578
rect 219256 573514 219308 573520
rect 219256 562420 219308 562426
rect 219256 562362 219308 562368
rect 219164 558272 219216 558278
rect 219164 558214 219216 558220
rect 218704 556844 218756 556850
rect 218704 556786 218756 556792
rect 219268 554963 219296 562362
rect 219636 557534 219664 639134
rect 223764 638240 223816 638246
rect 223764 638182 223816 638188
rect 223776 638042 223804 638182
rect 225800 638044 225828 640766
rect 272156 640756 272208 640762
rect 272156 640698 272208 640704
rect 243176 640688 243228 640694
rect 243176 640630 243228 640636
rect 231584 640348 231636 640354
rect 231584 640290 231636 640296
rect 228732 638104 228784 638110
rect 228784 638052 229034 638058
rect 228732 638046 229034 638052
rect 223764 638036 223816 638042
rect 228744 638030 229034 638046
rect 231596 638044 231624 640290
rect 234804 639260 234856 639266
rect 234804 639202 234856 639208
rect 234816 638044 234844 639202
rect 237380 639124 237432 639130
rect 237380 639066 237432 639072
rect 237392 638044 237420 639066
rect 243188 638044 243216 640630
rect 252192 640620 252244 640626
rect 252192 640562 252244 640568
rect 246396 639192 246448 639198
rect 246396 639134 246448 639140
rect 246408 638044 246436 639134
rect 252204 638044 252232 640562
rect 263784 640552 263836 640558
rect 263784 640494 263836 640500
rect 254768 639056 254820 639062
rect 254768 638998 254820 639004
rect 254780 638044 254808 638998
rect 263796 638044 263824 640494
rect 269580 640484 269632 640490
rect 269580 640426 269632 640432
rect 266280 638042 266386 638058
rect 269592 638044 269620 640426
rect 272168 638044 272196 640698
rect 275376 640416 275428 640422
rect 275376 640358 275428 640364
rect 275388 638044 275416 640358
rect 277952 638988 278004 638994
rect 277952 638930 278004 638936
rect 277964 638044 277992 638930
rect 266268 638036 266386 638042
rect 223764 637978 223816 637984
rect 266320 638030 266386 638036
rect 266268 637978 266320 637984
rect 222844 637968 222896 637974
rect 260196 637968 260248 637974
rect 222896 637916 223238 637922
rect 222844 637910 223238 637916
rect 222856 637894 223238 637910
rect 240336 637906 240626 637922
rect 260248 637916 260590 637922
rect 260196 637910 260590 637916
rect 240324 637900 240626 637906
rect 240376 637894 240626 637900
rect 260208 637894 260590 637910
rect 240324 637842 240376 637848
rect 248696 637832 248748 637838
rect 248748 637780 248998 637786
rect 248696 637774 248998 637780
rect 248708 637758 248998 637774
rect 257632 637770 258014 637786
rect 257620 637764 258014 637770
rect 257672 637758 258014 637764
rect 257620 637706 257672 637712
rect 219716 637696 219768 637702
rect 219768 637644 220018 637650
rect 219716 637638 220018 637644
rect 219728 637622 220018 637638
rect 280724 637498 280752 646614
rect 280712 637492 280764 637498
rect 280712 637434 280764 637440
rect 280554 637350 280844 637378
rect 280712 637288 280764 637294
rect 280712 637230 280764 637236
rect 219900 576224 219952 576230
rect 219900 576166 219952 576172
rect 219912 567194 219940 576166
rect 220004 571402 220032 575076
rect 222200 574932 222252 574938
rect 222200 574874 222252 574880
rect 219992 571396 220044 571402
rect 219992 571338 220044 571344
rect 221464 571396 221516 571402
rect 221464 571338 221516 571344
rect 219912 567166 220124 567194
rect 219636 557506 220032 557534
rect 220004 554963 220032 557506
rect 220096 556918 220124 567166
rect 220728 565412 220780 565418
rect 220728 565354 220780 565360
rect 220084 556912 220136 556918
rect 220084 556854 220136 556860
rect 220740 554963 220768 565354
rect 221476 554963 221504 571338
rect 222212 562426 222240 574874
rect 222292 572212 222344 572218
rect 222292 572154 222344 572160
rect 222200 562420 222252 562426
rect 222200 562362 222252 562368
rect 222304 555234 222332 572154
rect 222580 571402 222608 575076
rect 223580 575000 223632 575006
rect 223580 574942 223632 574948
rect 222568 571396 222620 571402
rect 222568 571338 222620 571344
rect 222844 562420 222896 562426
rect 222844 562362 222896 562368
rect 222228 555206 222332 555234
rect 222228 554948 222256 555206
rect 222856 554963 222884 562362
rect 223592 554963 223620 574942
rect 224316 573572 224368 573578
rect 224316 573514 224368 573520
rect 224328 554963 224356 573514
rect 224960 571396 225012 571402
rect 224960 571338 225012 571344
rect 225052 571396 225104 571402
rect 225052 571338 225104 571344
rect 224972 562426 225000 571338
rect 224960 562420 225012 562426
rect 224960 562362 225012 562368
rect 225064 554963 225092 571338
rect 225156 563990 225184 575076
rect 227904 572076 227956 572082
rect 227904 572018 227956 572024
rect 226432 566704 226484 566710
rect 226432 566646 226484 566652
rect 225144 563984 225196 563990
rect 225144 563926 225196 563932
rect 225788 562420 225840 562426
rect 225788 562362 225840 562368
rect 225800 554963 225828 562362
rect 226444 554963 226472 566646
rect 227168 558272 227220 558278
rect 227168 558214 227220 558220
rect 227180 554963 227208 558214
rect 227916 554963 227944 572018
rect 228376 571402 228404 575076
rect 230768 575062 230966 575090
rect 233252 575062 234186 575090
rect 236012 575062 236762 575090
rect 238772 575062 239982 575090
rect 241532 575062 242558 575090
rect 229284 574932 229336 574938
rect 229284 574874 229336 574880
rect 228364 571396 228416 571402
rect 228364 571338 228416 571344
rect 228640 565344 228692 565350
rect 228640 565286 228692 565292
rect 228652 554963 228680 565286
rect 229296 554963 229324 574874
rect 230020 556980 230072 556986
rect 230020 556922 230072 556928
rect 230032 554963 230060 556922
rect 230768 554963 230796 575062
rect 232228 572280 232280 572286
rect 232228 572222 232280 572228
rect 231492 556980 231544 556986
rect 231492 556922 231544 556928
rect 231504 554963 231532 556922
rect 232240 554963 232268 572222
rect 233252 566642 233280 575062
rect 233240 566636 233292 566642
rect 233240 566578 233292 566584
rect 234344 563712 234396 563718
rect 234344 563654 234396 563660
rect 232872 556912 232924 556918
rect 232872 556854 232924 556860
rect 232884 554963 232912 556854
rect 233608 556844 233660 556850
rect 233608 556786 233660 556792
rect 233620 554963 233648 556786
rect 234356 554963 234384 563654
rect 236012 561134 236040 575062
rect 236000 561128 236052 561134
rect 236000 561070 236052 561076
rect 235080 560992 235132 560998
rect 235080 560934 235132 560940
rect 235092 554963 235120 560934
rect 237932 559904 237984 559910
rect 237932 559846 237984 559852
rect 237196 556844 237248 556850
rect 237196 556786 237248 556792
rect 236476 555212 236528 555218
rect 236476 555154 236528 555160
rect 235844 555082 235948 555098
rect 235844 555076 235960 555082
rect 235844 555070 235908 555076
rect 235844 554948 235872 555070
rect 235908 555018 235960 555024
rect 236488 554948 236516 555154
rect 237208 554963 237236 556786
rect 237944 554963 237972 559846
rect 238772 556986 238800 575062
rect 240784 573572 240836 573578
rect 240784 573514 240836 573520
rect 238760 556980 238812 556986
rect 238760 556922 238812 556928
rect 239404 556980 239456 556986
rect 239404 556922 239456 556928
rect 238668 556912 238720 556918
rect 238668 556854 238720 556860
rect 238680 554963 238708 556854
rect 239416 554963 239444 556922
rect 240048 556436 240100 556442
rect 240048 556378 240100 556384
rect 240060 554963 240088 556378
rect 240796 554963 240824 573514
rect 241532 565214 241560 575062
rect 245764 572082 245792 575076
rect 247144 575062 248354 575090
rect 251192 575062 251574 575090
rect 245752 572076 245804 572082
rect 245752 572018 245804 572024
rect 247040 572076 247092 572082
rect 247040 572018 247092 572024
rect 245108 566568 245160 566574
rect 245108 566510 245160 566516
rect 241520 565208 241572 565214
rect 241520 565150 241572 565156
rect 242900 565208 242952 565214
rect 242900 565150 242952 565156
rect 242256 559020 242308 559026
rect 242256 558962 242308 558968
rect 241518 556200 241574 556209
rect 241518 556135 241574 556144
rect 241532 554963 241560 556135
rect 242268 554963 242296 558962
rect 242912 554963 242940 565150
rect 244372 558340 244424 558346
rect 244372 558282 244424 558288
rect 243636 555280 243688 555286
rect 243636 555222 243688 555228
rect 243648 554963 243676 555222
rect 244384 554963 244412 558282
rect 245120 554963 245148 566510
rect 246488 565276 246540 565282
rect 246488 565218 246540 565224
rect 245844 557048 245896 557054
rect 245844 556990 245896 556996
rect 245856 554963 245884 556990
rect 246500 554963 246528 565218
rect 247052 562306 247080 572018
rect 247144 565418 247172 575062
rect 250076 569424 250128 569430
rect 250076 569366 250128 569372
rect 247132 565412 247184 565418
rect 247132 565354 247184 565360
rect 247052 562278 247356 562306
rect 247224 557660 247276 557666
rect 247224 557602 247276 557608
rect 247236 554963 247264 557602
rect 247328 557534 247356 562278
rect 247328 557506 248000 557534
rect 247972 554963 248000 557506
rect 248694 556744 248750 556753
rect 248694 556679 248750 556688
rect 248708 554963 248736 556679
rect 249448 555144 249500 555150
rect 249448 555086 249500 555092
rect 249460 554948 249488 555086
rect 250088 554963 250116 569366
rect 250812 562284 250864 562290
rect 250812 562226 250864 562232
rect 250824 554963 250852 562226
rect 251192 558210 251220 575062
rect 254136 572218 254164 575076
rect 254124 572212 254176 572218
rect 254124 572154 254176 572160
rect 257356 572150 257384 575076
rect 259932 572286 259960 575076
rect 259920 572280 259972 572286
rect 259920 572222 259972 572228
rect 257344 572144 257396 572150
rect 257344 572086 257396 572092
rect 262864 571464 262916 571470
rect 262864 571406 262916 571412
rect 260104 571396 260156 571402
rect 260104 571338 260156 571344
rect 259460 568064 259512 568070
rect 259460 568006 259512 568012
rect 255320 567996 255372 568002
rect 255320 567938 255372 567944
rect 255332 562426 255360 567938
rect 257988 566636 258040 566642
rect 257988 566578 258040 566584
rect 255320 562420 255372 562426
rect 255320 562362 255372 562368
rect 256516 562420 256568 562426
rect 256516 562362 256568 562368
rect 251548 561128 251600 561134
rect 251548 561070 251600 561076
rect 251180 558204 251232 558210
rect 251180 558146 251232 558152
rect 251560 554963 251588 561070
rect 253664 559768 253716 559774
rect 253664 559710 253716 559716
rect 252284 557728 252336 557734
rect 252284 557670 252336 557676
rect 252296 554963 252324 557670
rect 252928 557252 252980 557258
rect 252928 557194 252980 557200
rect 252940 554963 252968 557194
rect 253676 554963 253704 559710
rect 254400 557796 254452 557802
rect 254400 557738 254452 557744
rect 254412 554963 254440 557738
rect 255872 557184 255924 557190
rect 255872 557126 255924 557132
rect 255134 556472 255190 556481
rect 255134 556407 255190 556416
rect 255148 554963 255176 556407
rect 255884 554963 255912 557126
rect 256528 554963 256556 562362
rect 257252 557320 257304 557326
rect 257252 557262 257304 557268
rect 257264 554963 257292 557262
rect 258000 554963 258028 566578
rect 258722 556608 258778 556617
rect 258722 556543 258778 556552
rect 258736 554963 258764 556543
rect 259472 554963 259500 568006
rect 260116 561202 260144 571338
rect 260196 563916 260248 563922
rect 260196 563858 260248 563864
rect 260104 561196 260156 561202
rect 260104 561138 260156 561144
rect 260208 555234 260236 563858
rect 262876 562562 262904 571406
rect 263152 571402 263180 575076
rect 263692 572144 263744 572150
rect 263692 572086 263744 572092
rect 263140 571396 263192 571402
rect 263140 571338 263192 571344
rect 262864 562556 262916 562562
rect 262864 562498 262916 562504
rect 260840 558000 260892 558006
rect 260840 557942 260892 557948
rect 260132 555206 260236 555234
rect 260132 554948 260160 555206
rect 260852 554963 260880 557942
rect 261576 557116 261628 557122
rect 261576 557058 261628 557064
rect 261588 554963 261616 557058
rect 262312 556504 262364 556510
rect 262312 556446 262364 556452
rect 262324 554963 262352 556446
rect 263048 555416 263100 555422
rect 263048 555358 263100 555364
rect 263060 554963 263088 555358
rect 263704 554963 263732 572086
rect 265728 571470 265756 575076
rect 268016 572756 268068 572762
rect 268016 572698 268068 572704
rect 267004 572552 267056 572558
rect 267004 572494 267056 572500
rect 265716 571464 265768 571470
rect 265716 571406 265768 571412
rect 266636 569492 266688 569498
rect 266636 569434 266688 569440
rect 266544 566772 266596 566778
rect 266544 566714 266596 566720
rect 265900 558204 265952 558210
rect 265900 558146 265952 558152
rect 264428 558068 264480 558074
rect 264428 558010 264480 558016
rect 264440 554963 264468 558010
rect 265164 555348 265216 555354
rect 265164 555290 265216 555296
rect 265176 554963 265204 555290
rect 265912 554963 265940 558146
rect 266360 556436 266412 556442
rect 266360 556378 266412 556384
rect 266372 555490 266400 556378
rect 266360 555484 266412 555490
rect 266360 555426 266412 555432
rect 266556 554963 266584 566714
rect 266648 557534 266676 569434
rect 267016 563854 267044 572494
rect 267004 563848 267056 563854
rect 267004 563790 267056 563796
rect 266648 557506 267320 557534
rect 267292 554963 267320 557506
rect 268028 554963 268056 572698
rect 268948 572558 268976 575076
rect 268936 572552 268988 572558
rect 268936 572494 268988 572500
rect 269672 572212 269724 572218
rect 269672 572154 269724 572160
rect 269488 559836 269540 559842
rect 269488 559778 269540 559784
rect 268752 555552 268804 555558
rect 268752 555494 268804 555500
rect 268764 554963 268792 555494
rect 269500 554963 269528 559778
rect 269684 557534 269712 572154
rect 271524 571402 271552 575076
rect 274652 575062 274758 575090
rect 273260 575000 273312 575006
rect 273260 574942 273312 574948
rect 269764 571396 269816 571402
rect 269764 571338 269816 571344
rect 271512 571396 271564 571402
rect 271512 571338 271564 571344
rect 269776 559570 269804 571338
rect 273272 562358 273300 574942
rect 273260 562352 273312 562358
rect 273260 562294 273312 562300
rect 274456 562352 274508 562358
rect 274456 562294 274508 562300
rect 269764 559564 269816 559570
rect 269764 559506 269816 559512
rect 271604 558272 271656 558278
rect 271604 558214 271656 558220
rect 269684 557506 270172 557534
rect 270144 554963 270172 557506
rect 270868 556708 270920 556714
rect 270868 556650 270920 556656
rect 270880 554963 270908 556650
rect 271616 554963 271644 558214
rect 273076 558136 273128 558142
rect 273076 558078 273128 558084
rect 272340 557864 272392 557870
rect 272340 557806 272392 557812
rect 272352 554963 272380 557806
rect 273088 554963 273116 558078
rect 273720 557932 273772 557938
rect 273720 557874 273772 557880
rect 273732 554963 273760 557874
rect 274468 554963 274496 562294
rect 274652 562290 274680 575062
rect 277320 572014 277348 575076
rect 277308 572008 277360 572014
rect 277308 571950 277360 571956
rect 280540 571402 280568 575076
rect 278044 571396 278096 571402
rect 278044 571338 278096 571344
rect 280528 571396 280580 571402
rect 280528 571338 280580 571344
rect 275192 562352 275244 562358
rect 275192 562294 275244 562300
rect 274640 562284 274692 562290
rect 274640 562226 274692 562232
rect 275204 554963 275232 562294
rect 278056 561066 278084 571338
rect 278044 561060 278096 561066
rect 278044 561002 278096 561008
rect 279516 561060 279568 561066
rect 279516 561002 279568 561008
rect 277308 557456 277360 557462
rect 277308 557398 277360 557404
rect 275928 556776 275980 556782
rect 275928 556718 275980 556724
rect 275940 554963 275968 556718
rect 276572 556232 276624 556238
rect 276572 556174 276624 556180
rect 276584 554963 276612 556174
rect 277320 554963 277348 557398
rect 278044 557388 278096 557394
rect 278044 557330 278096 557336
rect 278056 554963 278084 557330
rect 278780 555620 278832 555626
rect 278780 555562 278832 555568
rect 278792 554963 278820 555562
rect 279528 554963 279556 561002
rect 280724 557534 280752 637230
rect 280816 566710 280844 637350
rect 280894 610056 280950 610065
rect 280894 609991 280950 610000
rect 280804 566704 280856 566710
rect 280804 566646 280856 566652
rect 280908 562494 280936 609991
rect 280896 562488 280948 562494
rect 280896 562430 280948 562436
rect 280724 557506 280936 557534
rect 280160 556572 280212 556578
rect 280160 556514 280212 556520
rect 280172 554963 280200 556514
rect 280908 554963 280936 557506
rect 281000 556986 281028 648722
rect 289820 648712 289872 648718
rect 289820 648654 289872 648660
rect 284944 647624 284996 647630
rect 284944 647566 284996 647572
rect 281078 647320 281134 647329
rect 281078 647255 281134 647264
rect 281092 557054 281120 647255
rect 282184 646264 282236 646270
rect 282184 646206 282236 646212
rect 281630 634944 281686 634953
rect 281630 634879 281686 634888
rect 281170 589384 281226 589393
rect 281170 589319 281226 589328
rect 281184 570790 281212 589319
rect 281644 583370 281672 634879
rect 282090 632224 282146 632233
rect 282090 632159 282146 632168
rect 281722 626104 281778 626113
rect 281722 626039 281778 626048
rect 281632 583364 281684 583370
rect 281632 583306 281684 583312
rect 281630 583264 281686 583273
rect 281630 583199 281686 583208
rect 281262 579864 281318 579873
rect 281262 579799 281318 579808
rect 281276 574938 281304 579799
rect 281538 577144 281594 577153
rect 281538 577079 281594 577088
rect 281264 574932 281316 574938
rect 281264 574874 281316 574880
rect 281552 573442 281580 577079
rect 281644 574802 281672 583199
rect 281632 574796 281684 574802
rect 281632 574738 281684 574744
rect 281540 573436 281592 573442
rect 281540 573378 281592 573384
rect 281172 570784 281224 570790
rect 281172 570726 281224 570732
rect 281736 567866 281764 626039
rect 281906 601624 281962 601633
rect 281906 601559 281962 601568
rect 281814 595504 281870 595513
rect 281814 595439 281870 595448
rect 281724 567860 281776 567866
rect 281724 567802 281776 567808
rect 281828 563786 281856 595439
rect 281920 569294 281948 601559
rect 281998 598224 282054 598233
rect 281998 598159 282054 598168
rect 282012 574870 282040 598159
rect 282000 574864 282052 574870
rect 282000 574806 282052 574812
rect 281908 569288 281960 569294
rect 281908 569230 281960 569236
rect 282104 565350 282132 632159
rect 282092 565344 282144 565350
rect 282092 565286 282144 565292
rect 281816 563780 281868 563786
rect 281816 563722 281868 563728
rect 282196 557122 282224 646206
rect 283470 628824 283526 628833
rect 283470 628759 283526 628768
rect 283010 622704 283066 622713
rect 283010 622639 283066 622648
rect 282918 592104 282974 592113
rect 282918 592039 282974 592048
rect 282276 583364 282328 583370
rect 282276 583306 282328 583312
rect 282288 570722 282316 583306
rect 282932 573510 282960 592039
rect 282920 573504 282972 573510
rect 282920 573446 282972 573452
rect 282276 570716 282328 570722
rect 282276 570658 282328 570664
rect 283024 569362 283052 622639
rect 283378 619984 283434 619993
rect 283378 619919 283434 619928
rect 283286 616584 283342 616593
rect 283286 616519 283342 616528
rect 283102 613864 283158 613873
rect 283102 613799 283158 613808
rect 283012 569356 283064 569362
rect 283012 569298 283064 569304
rect 283116 565146 283144 613799
rect 283194 607744 283250 607753
rect 283194 607679 283250 607688
rect 283104 565140 283156 565146
rect 283104 565082 283156 565088
rect 283208 559706 283236 607679
rect 283300 567934 283328 616519
rect 283392 573374 283420 619919
rect 283380 573368 283432 573374
rect 283380 573310 283432 573316
rect 283288 567928 283340 567934
rect 283288 567870 283340 567876
rect 283196 559700 283248 559706
rect 283196 559642 283248 559648
rect 283484 559638 283512 628759
rect 283654 604344 283710 604353
rect 283654 604279 283710 604288
rect 283668 603158 283696 604279
rect 283656 603152 283708 603158
rect 283656 603094 283708 603100
rect 283562 585984 283618 585993
rect 283562 585919 283618 585928
rect 283576 566506 283604 585919
rect 284956 566778 284984 647566
rect 288532 646400 288584 646406
rect 288532 646342 288584 646348
rect 288440 646060 288492 646066
rect 288440 646002 288492 646008
rect 287704 640348 287756 640354
rect 287704 640290 287756 640296
rect 286324 611380 286376 611386
rect 286324 611322 286376 611328
rect 286336 572218 286364 611322
rect 286416 597576 286468 597582
rect 286416 597518 286468 597524
rect 286428 575482 286456 597518
rect 286416 575476 286468 575482
rect 286416 575418 286468 575424
rect 286324 572212 286376 572218
rect 286324 572154 286376 572160
rect 284944 566772 284996 566778
rect 284944 566714 284996 566720
rect 283564 566500 283616 566506
rect 283564 566442 283616 566448
rect 283748 561876 283800 561882
rect 283748 561818 283800 561824
rect 283472 559632 283524 559638
rect 283472 559574 283524 559580
rect 282368 559564 282420 559570
rect 282368 559506 282420 559512
rect 282184 557116 282236 557122
rect 282184 557058 282236 557064
rect 281080 557048 281132 557054
rect 281080 556990 281132 556996
rect 280988 556980 281040 556986
rect 280988 556922 281040 556928
rect 281632 556436 281684 556442
rect 281632 556378 281684 556384
rect 281644 554963 281672 556378
rect 282380 554963 282408 559506
rect 283104 556368 283156 556374
rect 283104 556310 283156 556316
rect 283116 554963 283144 556310
rect 283760 554963 283788 561818
rect 286692 559428 286744 559434
rect 286692 559370 286744 559376
rect 285220 559292 285272 559298
rect 285220 559234 285272 559240
rect 284944 559224 284996 559230
rect 284944 559166 284996 559172
rect 284484 559156 284536 559162
rect 284484 559098 284536 559104
rect 284208 559088 284260 559094
rect 284208 559030 284260 559036
rect 284220 556850 284248 559030
rect 284208 556844 284260 556850
rect 284208 556786 284260 556792
rect 284496 554963 284524 559098
rect 284956 556918 284984 559166
rect 284944 556912 284996 556918
rect 284944 556854 284996 556860
rect 285232 554963 285260 559234
rect 285956 556640 286008 556646
rect 285956 556582 286008 556588
rect 285968 554963 285996 556582
rect 286704 554963 286732 559370
rect 287716 558278 287744 640290
rect 287796 621036 287848 621042
rect 287796 620978 287848 620984
rect 287808 561882 287836 620978
rect 287796 561876 287848 561882
rect 287796 561818 287848 561824
rect 288072 559360 288124 559366
rect 288072 559302 288124 559308
rect 287704 558272 287756 558278
rect 287704 558214 287756 558220
rect 287336 557592 287388 557598
rect 287336 557534 287388 557540
rect 287348 554963 287376 557534
rect 288084 554963 288112 559302
rect 288452 557534 288480 646002
rect 288544 576854 288572 646342
rect 289084 634840 289136 634846
rect 289084 634782 289136 634788
rect 288544 576826 289032 576854
rect 289004 557534 289032 576826
rect 289096 561066 289124 634782
rect 289176 586560 289228 586566
rect 289176 586502 289228 586508
rect 289188 563922 289216 586502
rect 289832 576854 289860 648654
rect 289832 576826 290228 576854
rect 289176 563916 289228 563922
rect 289176 563858 289228 563864
rect 289084 561060 289136 561066
rect 289084 561002 289136 561008
rect 288452 557506 288848 557534
rect 289004 557506 289584 557534
rect 288820 554963 288848 557506
rect 289556 554963 289584 557506
rect 290200 554963 290228 576826
rect 291212 557534 291240 650014
rect 298744 648032 298796 648038
rect 298744 647974 298796 647980
rect 296720 646604 296772 646610
rect 296720 646546 296772 646552
rect 291292 646468 291344 646474
rect 291292 646410 291344 646416
rect 291304 576854 291332 646410
rect 293960 646196 294012 646202
rect 293960 646138 294012 646144
rect 291304 576826 292436 576854
rect 291212 557506 291700 557534
rect 290922 556336 290978 556345
rect 290922 556271 290978 556280
rect 290936 554963 290964 556271
rect 291672 554963 291700 557506
rect 292408 554963 292436 576826
rect 293776 559496 293828 559502
rect 293776 559438 293828 559444
rect 293132 558952 293184 558958
rect 293132 558894 293184 558900
rect 293144 554963 293172 558894
rect 293788 554963 293816 559438
rect 293972 556306 294000 646138
rect 295984 615528 296036 615534
rect 295984 615470 296036 615476
rect 295996 569430 296024 615470
rect 296076 601724 296128 601730
rect 296076 601666 296128 601672
rect 295984 569424 296036 569430
rect 295984 569366 296036 569372
rect 296088 559570 296116 601666
rect 296076 559564 296128 559570
rect 296076 559506 296128 559512
rect 296732 556306 296760 646546
rect 298100 646536 298152 646542
rect 298100 646478 298152 646484
rect 296812 646128 296864 646134
rect 296812 646070 296864 646076
rect 293960 556300 294012 556306
rect 293960 556242 294012 556248
rect 295248 556300 295300 556306
rect 295248 556242 295300 556248
rect 296720 556300 296772 556306
rect 296720 556242 296772 556248
rect 294512 555688 294564 555694
rect 294512 555630 294564 555636
rect 294524 554963 294552 555630
rect 295260 554963 295288 556242
rect 295984 555756 296036 555762
rect 295984 555698 296036 555704
rect 295996 554963 296024 555698
rect 296824 555234 296852 646070
rect 298112 567194 298140 646478
rect 298756 569498 298784 647974
rect 302884 644496 302936 644502
rect 302884 644438 302936 644444
rect 300216 603152 300268 603158
rect 300216 603094 300268 603100
rect 300124 592068 300176 592074
rect 300124 592010 300176 592016
rect 298744 569492 298796 569498
rect 298744 569434 298796 569440
rect 298112 567166 298876 567194
rect 297364 556300 297416 556306
rect 297364 556242 297416 556248
rect 298100 556300 298152 556306
rect 298100 556242 298152 556248
rect 296748 555206 296852 555234
rect 296748 554948 296776 555206
rect 297376 554963 297404 556242
rect 298112 554963 298140 556242
rect 298848 554963 298876 567166
rect 300136 559842 300164 592010
rect 300228 584186 300256 603094
rect 300216 584180 300268 584186
rect 300216 584122 300268 584128
rect 302240 584180 302292 584186
rect 302240 584122 302292 584128
rect 302252 575414 302280 584122
rect 302240 575408 302292 575414
rect 302240 575350 302292 575356
rect 302252 574122 302280 575350
rect 302240 574116 302292 574122
rect 302240 574058 302292 574064
rect 302896 568070 302924 644438
rect 302976 574116 303028 574122
rect 302976 574058 303028 574064
rect 302884 568064 302936 568070
rect 302884 568006 302936 568012
rect 300124 559836 300176 559842
rect 300124 559778 300176 559784
rect 301504 558204 301556 558210
rect 301504 558146 301556 558152
rect 299572 556844 299624 556850
rect 299572 556786 299624 556792
rect 299584 554963 299612 556786
rect 300400 556776 300452 556782
rect 300400 556718 300452 556724
rect 300674 556744 300730 556753
rect 300216 556708 300268 556714
rect 300216 556650 300268 556656
rect 300124 556436 300176 556442
rect 300124 556378 300176 556384
rect 300136 533594 300164 556378
rect 300124 533588 300176 533594
rect 300124 533530 300176 533536
rect 300228 533526 300256 556650
rect 300308 556504 300360 556510
rect 300308 556446 300360 556452
rect 300216 533520 300268 533526
rect 300216 533462 300268 533468
rect 300320 533186 300348 556446
rect 300412 534206 300440 556718
rect 300674 556679 300730 556688
rect 300490 556472 300546 556481
rect 300490 556407 300546 556416
rect 300504 535226 300532 556407
rect 300492 535220 300544 535226
rect 300492 535162 300544 535168
rect 300688 535158 300716 556679
rect 300768 555620 300820 555626
rect 300768 555562 300820 555568
rect 300780 554742 300808 555562
rect 301412 555212 301464 555218
rect 301412 555154 301464 555160
rect 300768 554736 300820 554742
rect 300768 554678 300820 554684
rect 301424 550594 301452 555154
rect 301412 550588 301464 550594
rect 301412 550530 301464 550536
rect 300676 535152 300728 535158
rect 300676 535094 300728 535100
rect 300400 534200 300452 534206
rect 300400 534142 300452 534148
rect 300308 533180 300360 533186
rect 300308 533122 300360 533128
rect 301516 532370 301544 558146
rect 301688 557456 301740 557462
rect 301688 557398 301740 557404
rect 301596 556368 301648 556374
rect 301596 556310 301648 556316
rect 301608 533390 301636 556310
rect 301700 533458 301728 557398
rect 301780 557184 301832 557190
rect 301780 557126 301832 557132
rect 301688 533452 301740 533458
rect 301688 533394 301740 533400
rect 301596 533384 301648 533390
rect 301596 533326 301648 533332
rect 301792 533254 301820 557126
rect 301872 556232 301924 556238
rect 301872 556174 301924 556180
rect 301884 533322 301912 556174
rect 302884 555552 302936 555558
rect 302884 555494 302936 555500
rect 301964 555416 302016 555422
rect 301964 555358 302016 555364
rect 301872 533316 301924 533322
rect 301872 533258 301924 533264
rect 301780 533248 301832 533254
rect 301780 533190 301832 533196
rect 301504 532364 301556 532370
rect 301504 532306 301556 532312
rect 301976 531826 302004 555358
rect 302330 532536 302386 532545
rect 302330 532471 302386 532480
rect 301964 531820 302016 531826
rect 301964 531762 302016 531768
rect 302344 529242 302372 532471
rect 302896 532438 302924 555494
rect 302988 533866 303016 574058
rect 304276 564398 304304 700266
rect 304264 564392 304316 564398
rect 304264 564334 304316 564340
rect 304356 558068 304408 558074
rect 304356 558010 304408 558016
rect 304264 558000 304316 558006
rect 304264 557942 304316 557948
rect 303068 557320 303120 557326
rect 303068 557262 303120 557268
rect 303080 535090 303108 557262
rect 303158 556608 303214 556617
rect 303158 556543 303214 556552
rect 303172 535537 303200 556543
rect 303250 547496 303306 547505
rect 303250 547431 303306 547440
rect 303158 535528 303214 535537
rect 303158 535463 303214 535472
rect 303068 535084 303120 535090
rect 303068 535026 303120 535032
rect 302976 533860 303028 533866
rect 302976 533802 303028 533808
rect 302884 532432 302936 532438
rect 302884 532374 302936 532380
rect 302332 529236 302384 529242
rect 302332 529178 302384 529184
rect 57716 528526 57928 528554
rect 57716 525094 57744 528526
rect 42708 525088 42760 525094
rect 57704 525088 57756 525094
rect 42708 525030 42760 525036
rect 57702 525056 57704 525065
rect 57756 525056 57758 525065
rect 42338 486432 42394 486441
rect 42338 486367 42394 486376
rect 42248 483948 42300 483954
rect 42248 483890 42300 483896
rect 42156 468784 42208 468790
rect 42156 468726 42208 468732
rect 40684 371204 40736 371210
rect 40684 371146 40736 371152
rect 42168 264858 42196 468726
rect 42156 264852 42208 264858
rect 42156 264794 42208 264800
rect 42260 260166 42288 483890
rect 42248 260160 42300 260166
rect 42248 260102 42300 260108
rect 42352 238678 42380 486367
rect 42616 469124 42668 469130
rect 42616 469066 42668 469072
rect 42524 469056 42576 469062
rect 42524 468998 42576 469004
rect 42432 468988 42484 468994
rect 42432 468930 42484 468936
rect 42340 238672 42392 238678
rect 42340 238614 42392 238620
rect 42444 154698 42472 468930
rect 42432 154692 42484 154698
rect 42432 154634 42484 154640
rect 11704 120080 11756 120086
rect 11704 120022 11756 120028
rect 3424 44056 3476 44062
rect 3422 44024 3424 44033
rect 7564 44056 7616 44062
rect 3476 44024 3478 44033
rect 7564 43998 7616 44004
rect 3422 43959 3478 43968
rect 42536 43586 42564 468998
rect 42524 43580 42576 43586
rect 42524 43522 42576 43528
rect 42628 41206 42656 469066
rect 42720 382226 42748 525030
rect 57702 524991 57758 525000
rect 302988 517585 303016 533802
rect 303264 530602 303292 547431
rect 304276 532710 304304 557942
rect 304264 532704 304316 532710
rect 304264 532646 304316 532652
rect 304368 532234 304396 558010
rect 305656 534138 305684 700334
rect 315040 698970 315068 703520
rect 345768 701010 345796 703520
rect 345756 701004 345808 701010
rect 345756 700946 345808 700952
rect 315028 698964 315080 698970
rect 315028 698906 315080 698912
rect 316684 684548 316736 684554
rect 316684 684490 316736 684496
rect 312544 648100 312596 648106
rect 312544 648042 312596 648048
rect 309782 647456 309838 647465
rect 309782 647391 309838 647400
rect 307024 630692 307076 630698
rect 307024 630634 307076 630640
rect 305736 555280 305788 555286
rect 305736 555222 305788 555228
rect 305748 545086 305776 555222
rect 305736 545080 305788 545086
rect 305736 545022 305788 545028
rect 305644 534132 305696 534138
rect 305644 534074 305696 534080
rect 304356 532228 304408 532234
rect 304356 532170 304408 532176
rect 303252 530596 303304 530602
rect 303252 530538 303304 530544
rect 302974 517576 303030 517585
rect 302974 517511 303030 517520
rect 302882 502616 302938 502625
rect 302882 502551 302938 502560
rect 302896 502382 302924 502551
rect 302884 502376 302936 502382
rect 302884 502318 302936 502324
rect 60108 495094 60214 495122
rect 299782 495094 299888 495122
rect 56324 493400 56376 493406
rect 56324 493342 56376 493348
rect 51816 493332 51868 493338
rect 51816 493274 51868 493280
rect 50896 492516 50948 492522
rect 50896 492458 50948 492464
rect 50528 492448 50580 492454
rect 50528 492390 50580 492396
rect 49148 492108 49200 492114
rect 49148 492050 49200 492056
rect 43904 491972 43956 491978
rect 43904 491914 43956 491920
rect 43718 486840 43774 486849
rect 43718 486775 43774 486784
rect 43628 484016 43680 484022
rect 43628 483958 43680 483964
rect 43352 483744 43404 483750
rect 43352 483686 43404 483692
rect 42708 382220 42760 382226
rect 42708 382162 42760 382168
rect 43364 373862 43392 483686
rect 43536 468852 43588 468858
rect 43536 468794 43588 468800
rect 43444 468580 43496 468586
rect 43444 468522 43496 468528
rect 43352 373856 43404 373862
rect 43352 373798 43404 373804
rect 43456 264382 43484 468522
rect 43548 264722 43576 468794
rect 43536 264716 43588 264722
rect 43536 264658 43588 264664
rect 43444 264376 43496 264382
rect 43444 264318 43496 264324
rect 43640 259282 43668 483958
rect 43732 259418 43760 486775
rect 43810 486704 43866 486713
rect 43810 486639 43866 486648
rect 43720 259412 43772 259418
rect 43720 259354 43772 259360
rect 43628 259276 43680 259282
rect 43628 259218 43680 259224
rect 43824 238474 43852 486639
rect 43812 238468 43864 238474
rect 43812 238410 43864 238416
rect 43916 154630 43944 491914
rect 48228 489728 48280 489734
rect 48228 489670 48280 489676
rect 48044 489660 48096 489666
rect 48044 489602 48096 489608
rect 46572 489592 46624 489598
rect 46572 489534 46624 489540
rect 46296 489524 46348 489530
rect 46296 489466 46348 489472
rect 45468 484084 45520 484090
rect 45468 484026 45520 484032
rect 45376 468716 45428 468722
rect 45376 468658 45428 468664
rect 45284 468648 45336 468654
rect 45284 468590 45336 468596
rect 44088 468444 44140 468450
rect 44088 468386 44140 468392
rect 43996 460420 44048 460426
rect 43996 460362 44048 460368
rect 43904 154624 43956 154630
rect 43904 154566 43956 154572
rect 44008 42362 44036 460362
rect 43996 42356 44048 42362
rect 43996 42298 44048 42304
rect 42616 41200 42668 41206
rect 42616 41142 42668 41148
rect 44100 39778 44128 468386
rect 45192 466404 45244 466410
rect 45192 466346 45244 466352
rect 45100 466336 45152 466342
rect 45100 466278 45152 466284
rect 44732 465656 44784 465662
rect 44732 465598 44784 465604
rect 44640 462800 44692 462806
rect 44640 462742 44692 462748
rect 44652 371482 44680 462742
rect 44640 371476 44692 371482
rect 44640 371418 44692 371424
rect 44744 371414 44772 465598
rect 44824 465588 44876 465594
rect 44824 465530 44876 465536
rect 44732 371408 44784 371414
rect 44732 371350 44784 371356
rect 44836 371346 44864 465530
rect 44916 465520 44968 465526
rect 44916 465462 44968 465468
rect 44824 371340 44876 371346
rect 44824 371282 44876 371288
rect 44928 371278 44956 465462
rect 45008 460284 45060 460290
rect 45008 460226 45060 460232
rect 44916 371272 44968 371278
rect 44916 371214 44968 371220
rect 45020 264790 45048 460226
rect 45008 264784 45060 264790
rect 45008 264726 45060 264732
rect 45112 264586 45140 466278
rect 45204 264654 45232 466346
rect 45192 264648 45244 264654
rect 45192 264590 45244 264596
rect 45100 264580 45152 264586
rect 45100 264522 45152 264528
rect 45296 264314 45324 468590
rect 45284 264308 45336 264314
rect 45284 264250 45336 264256
rect 45388 264246 45416 468658
rect 45376 264240 45428 264246
rect 45376 264182 45428 264188
rect 45480 260234 45508 484026
rect 46112 483812 46164 483818
rect 46112 483754 46164 483760
rect 46020 483676 46072 483682
rect 46020 483618 46072 483624
rect 46032 385014 46060 483618
rect 46020 385008 46072 385014
rect 46020 384950 46072 384956
rect 46124 373522 46152 483754
rect 46204 468920 46256 468926
rect 46204 468862 46256 468868
rect 46112 373516 46164 373522
rect 46112 373458 46164 373464
rect 46112 371340 46164 371346
rect 46112 371282 46164 371288
rect 45468 260228 45520 260234
rect 45468 260170 45520 260176
rect 46124 241466 46152 371282
rect 46216 264518 46244 468862
rect 46308 276010 46336 489466
rect 46388 486804 46440 486810
rect 46388 486746 46440 486752
rect 46296 276004 46348 276010
rect 46296 275946 46348 275952
rect 46204 264512 46256 264518
rect 46204 264454 46256 264460
rect 46400 264178 46428 486746
rect 46480 486736 46532 486742
rect 46480 486678 46532 486684
rect 46388 264172 46440 264178
rect 46388 264114 46440 264120
rect 46492 264110 46520 486678
rect 46480 264104 46532 264110
rect 46480 264046 46532 264052
rect 46584 263265 46612 489534
rect 46846 489152 46902 489161
rect 46846 489087 46902 489096
rect 46664 486872 46716 486878
rect 46664 486814 46716 486820
rect 46570 263256 46626 263265
rect 46570 263191 46626 263200
rect 46478 260400 46534 260409
rect 46478 260335 46534 260344
rect 46204 260160 46256 260166
rect 46204 260102 46256 260108
rect 46386 260128 46442 260137
rect 46112 241460 46164 241466
rect 46112 241402 46164 241408
rect 46216 133346 46244 260102
rect 46386 260063 46442 260072
rect 46296 241460 46348 241466
rect 46296 241402 46348 241408
rect 46308 241330 46336 241402
rect 46296 241324 46348 241330
rect 46296 241266 46348 241272
rect 46308 133686 46336 241266
rect 46400 154018 46428 260063
rect 46388 154012 46440 154018
rect 46388 153954 46440 153960
rect 46492 151094 46520 260335
rect 46480 151088 46532 151094
rect 46480 151030 46532 151036
rect 46296 133680 46348 133686
rect 46296 133622 46348 133628
rect 46204 133340 46256 133346
rect 46204 133282 46256 133288
rect 46584 130286 46612 263191
rect 46676 259350 46704 486814
rect 46754 486568 46810 486577
rect 46754 486503 46810 486512
rect 46664 259344 46716 259350
rect 46664 259286 46716 259292
rect 46768 238678 46796 486503
rect 46860 238746 46888 489087
rect 47952 486532 48004 486538
rect 47952 486474 48004 486480
rect 47860 486464 47912 486470
rect 47860 486406 47912 486412
rect 47584 461644 47636 461650
rect 47584 461586 47636 461592
rect 47492 458312 47544 458318
rect 47492 458254 47544 458260
rect 47504 411262 47532 458254
rect 47596 412622 47624 461586
rect 47676 460216 47728 460222
rect 47676 460158 47728 460164
rect 47584 412616 47636 412622
rect 47584 412558 47636 412564
rect 47492 411256 47544 411262
rect 47492 411198 47544 411204
rect 47584 408536 47636 408542
rect 47584 408478 47636 408484
rect 47492 407176 47544 407182
rect 47492 407118 47544 407124
rect 47400 405748 47452 405754
rect 47400 405690 47452 405696
rect 47412 373998 47440 405690
rect 47504 375018 47532 407118
rect 47596 375086 47624 408478
rect 47584 375080 47636 375086
rect 47584 375022 47636 375028
rect 47492 375012 47544 375018
rect 47492 374954 47544 374960
rect 47400 373992 47452 373998
rect 47400 373934 47452 373940
rect 47492 371476 47544 371482
rect 47492 371418 47544 371424
rect 47504 241398 47532 371418
rect 47584 371408 47636 371414
rect 47584 371350 47636 371356
rect 47492 241392 47544 241398
rect 47492 241334 47544 241340
rect 47596 241262 47624 371350
rect 47688 371210 47716 460158
rect 47768 460080 47820 460086
rect 47768 460022 47820 460028
rect 47676 371204 47728 371210
rect 47676 371146 47728 371152
rect 47780 371142 47808 460022
rect 47872 373318 47900 486406
rect 47964 383654 47992 486474
rect 47952 383648 48004 383654
rect 47952 383590 48004 383596
rect 47952 380928 48004 380934
rect 47952 380870 48004 380876
rect 47860 373312 47912 373318
rect 47860 373254 47912 373260
rect 47860 371272 47912 371278
rect 47860 371214 47912 371220
rect 47768 371136 47820 371142
rect 47768 371078 47820 371084
rect 47872 241466 47900 371214
rect 47860 241460 47912 241466
rect 47860 241402 47912 241408
rect 47584 241256 47636 241262
rect 47584 241198 47636 241204
rect 47596 238754 47624 241198
rect 46848 238740 46900 238746
rect 47596 238726 47808 238754
rect 46848 238682 46900 238688
rect 46756 238672 46808 238678
rect 46756 238614 46808 238620
rect 47780 133754 47808 238726
rect 47964 238610 47992 380870
rect 48056 292534 48084 489602
rect 48136 469192 48188 469198
rect 48136 469134 48188 469140
rect 48044 292528 48096 292534
rect 48044 292470 48096 292476
rect 48148 264450 48176 469134
rect 48136 264444 48188 264450
rect 48136 264386 48188 264392
rect 48240 263129 48268 489670
rect 48964 489388 49016 489394
rect 48964 489330 49016 489336
rect 48688 489252 48740 489258
rect 48688 489194 48740 489200
rect 48700 373386 48728 489194
rect 48780 484220 48832 484226
rect 48780 484162 48832 484168
rect 48792 380934 48820 484162
rect 48872 483880 48924 483886
rect 48872 483822 48924 483828
rect 48780 380928 48832 380934
rect 48780 380870 48832 380876
rect 48884 373590 48912 483822
rect 48872 373584 48924 373590
rect 48872 373526 48924 373532
rect 48688 373380 48740 373386
rect 48688 373322 48740 373328
rect 48872 264988 48924 264994
rect 48872 264930 48924 264936
rect 48226 263120 48282 263129
rect 48226 263055 48282 263064
rect 48044 241460 48096 241466
rect 48044 241402 48096 241408
rect 47952 238604 48004 238610
rect 47952 238546 48004 238552
rect 47964 150414 47992 238546
rect 47952 150408 48004 150414
rect 47952 150350 48004 150356
rect 48056 133822 48084 241402
rect 48136 241392 48188 241398
rect 48136 241334 48188 241340
rect 48148 241194 48176 241334
rect 48136 241188 48188 241194
rect 48136 241130 48188 241136
rect 48044 133816 48096 133822
rect 48044 133758 48096 133764
rect 47768 133748 47820 133754
rect 47768 133690 47820 133696
rect 48148 130354 48176 241130
rect 48136 130348 48188 130354
rect 48136 130290 48188 130296
rect 46572 130280 46624 130286
rect 46572 130222 46624 130228
rect 48240 130218 48268 263055
rect 48884 130422 48912 264930
rect 48976 263401 49004 489330
rect 49054 489288 49110 489297
rect 49054 489223 49110 489232
rect 48962 263392 49018 263401
rect 48962 263327 49018 263336
rect 48976 130762 49004 263327
rect 49068 262857 49096 489223
rect 49054 262848 49110 262857
rect 49160 262818 49188 492050
rect 50540 491337 50568 492390
rect 50526 491328 50582 491337
rect 50526 491263 50582 491272
rect 50344 489864 50396 489870
rect 50344 489806 50396 489812
rect 49516 466132 49568 466138
rect 49516 466074 49568 466080
rect 49422 463040 49478 463049
rect 49422 462975 49478 462984
rect 49330 462904 49386 462913
rect 49330 462839 49386 462848
rect 49240 460896 49292 460902
rect 49240 460838 49292 460844
rect 49252 459649 49280 460838
rect 49238 459640 49294 459649
rect 49238 459575 49294 459584
rect 49240 456136 49292 456142
rect 49240 456078 49292 456084
rect 49054 262783 49110 262792
rect 49148 262812 49200 262818
rect 49148 262754 49200 262760
rect 49056 260432 49108 260438
rect 49056 260374 49108 260380
rect 49068 260234 49096 260374
rect 49056 260228 49108 260234
rect 49056 260170 49108 260176
rect 49068 151162 49096 260170
rect 49252 152386 49280 456078
rect 49344 152697 49372 462839
rect 49436 152969 49464 462975
rect 49528 154426 49556 466074
rect 50252 465792 50304 465798
rect 50252 465734 50304 465740
rect 49608 463548 49660 463554
rect 49608 463490 49660 463496
rect 49620 456142 49648 463490
rect 50160 460148 50212 460154
rect 50160 460090 50212 460096
rect 49608 456136 49660 456142
rect 49608 456078 49660 456084
rect 49606 381032 49662 381041
rect 49606 380967 49662 380976
rect 49516 154420 49568 154426
rect 49516 154362 49568 154368
rect 49422 152960 49478 152969
rect 49422 152895 49478 152904
rect 49330 152688 49386 152697
rect 49330 152623 49386 152632
rect 49240 152380 49292 152386
rect 49240 152322 49292 152328
rect 49056 151156 49108 151162
rect 49056 151098 49108 151104
rect 48964 130756 49016 130762
rect 48964 130698 49016 130704
rect 48872 130416 48924 130422
rect 48872 130358 48924 130364
rect 48228 130212 48280 130218
rect 48228 130154 48280 130160
rect 49620 43450 49648 380967
rect 49608 43444 49660 43450
rect 49608 43386 49660 43392
rect 50172 42158 50200 460090
rect 50264 263022 50292 465734
rect 50252 263016 50304 263022
rect 50252 262958 50304 262964
rect 50356 262954 50384 489806
rect 50526 489560 50582 489569
rect 50526 489495 50582 489504
rect 50436 489116 50488 489122
rect 50436 489058 50488 489064
rect 50344 262948 50396 262954
rect 50344 262890 50396 262896
rect 50448 262886 50476 489058
rect 50436 262880 50488 262886
rect 50436 262822 50488 262828
rect 50434 260808 50490 260817
rect 50434 260743 50490 260752
rect 50448 260273 50476 260743
rect 50540 260710 50568 489495
rect 50618 489424 50674 489433
rect 50618 489359 50674 489368
rect 50528 260704 50580 260710
rect 50528 260646 50580 260652
rect 50434 260264 50490 260273
rect 50434 260199 50490 260208
rect 50344 237448 50396 237454
rect 50344 237390 50396 237396
rect 50356 154562 50384 237390
rect 50344 154556 50396 154562
rect 50344 154498 50396 154504
rect 50448 130665 50476 260199
rect 50434 130656 50490 130665
rect 50434 130591 50490 130600
rect 50540 129742 50568 260646
rect 50632 240106 50660 489359
rect 50804 486600 50856 486606
rect 50804 486542 50856 486548
rect 50712 466200 50764 466206
rect 50712 466142 50764 466148
rect 50620 240100 50672 240106
rect 50620 240042 50672 240048
rect 50724 154494 50752 466142
rect 50816 411126 50844 486542
rect 50804 411120 50856 411126
rect 50804 411062 50856 411068
rect 50804 404388 50856 404394
rect 50804 404330 50856 404336
rect 50816 373969 50844 404330
rect 50802 373960 50858 373969
rect 50802 373895 50858 373904
rect 50804 239488 50856 239494
rect 50804 239430 50856 239436
rect 50816 238746 50844 239430
rect 50804 238740 50856 238746
rect 50804 238682 50856 238688
rect 50816 237454 50844 238682
rect 50804 237448 50856 237454
rect 50804 237390 50856 237396
rect 50712 154488 50764 154494
rect 50712 154430 50764 154436
rect 50908 152454 50936 492458
rect 51724 489456 51776 489462
rect 51724 489398 51776 489404
rect 51632 465724 51684 465730
rect 51632 465666 51684 465672
rect 50988 460828 51040 460834
rect 50988 460770 51040 460776
rect 51000 459649 51028 460770
rect 50986 459640 51042 459649
rect 50986 459575 51042 459584
rect 51540 459196 51592 459202
rect 51540 459138 51592 459144
rect 50988 403028 51040 403034
rect 50988 402970 51040 402976
rect 51000 375442 51028 402970
rect 51000 375414 51120 375442
rect 50986 375320 51042 375329
rect 50986 375255 51042 375264
rect 50896 152448 50948 152454
rect 50896 152390 50948 152396
rect 50528 129736 50580 129742
rect 50528 129678 50580 129684
rect 51000 42770 51028 375255
rect 51092 375057 51120 375414
rect 51078 375048 51134 375057
rect 51078 374983 51134 374992
rect 51552 264926 51580 459138
rect 51540 264920 51592 264926
rect 51540 264862 51592 264868
rect 51446 263664 51502 263673
rect 51446 263599 51502 263608
rect 51460 44198 51488 263599
rect 51644 263158 51672 465666
rect 51632 263152 51684 263158
rect 51632 263094 51684 263100
rect 51736 260642 51764 489398
rect 51828 263090 51856 493274
rect 53380 492176 53432 492182
rect 53380 492118 53432 492124
rect 52368 491768 52420 491774
rect 52368 491710 52420 491716
rect 52380 491337 52408 491710
rect 52366 491328 52422 491337
rect 52366 491263 52422 491272
rect 53196 487144 53248 487150
rect 53196 487086 53248 487092
rect 52092 466268 52144 466274
rect 52092 466210 52144 466216
rect 52000 463412 52052 463418
rect 52000 463354 52052 463360
rect 51908 460352 51960 460358
rect 51908 460294 51960 460300
rect 51816 263084 51868 263090
rect 51816 263026 51868 263032
rect 51724 260636 51776 260642
rect 51724 260578 51776 260584
rect 51632 260228 51684 260234
rect 51632 260170 51684 260176
rect 51644 259282 51672 260170
rect 51632 259276 51684 259282
rect 51632 259218 51684 259224
rect 51540 237448 51592 237454
rect 51540 237390 51592 237396
rect 51552 133278 51580 237390
rect 51540 133272 51592 133278
rect 51540 133214 51592 133220
rect 51644 132433 51672 259218
rect 51630 132424 51686 132433
rect 51630 132359 51686 132368
rect 51736 130898 51764 260578
rect 51816 239420 51868 239426
rect 51816 239362 51868 239368
rect 51828 238678 51856 239362
rect 51816 238672 51868 238678
rect 51816 238614 51868 238620
rect 51828 237454 51856 238614
rect 51816 237448 51868 237454
rect 51816 237390 51868 237396
rect 51816 154556 51868 154562
rect 51816 154498 51868 154504
rect 51828 153406 51856 154498
rect 51816 153400 51868 153406
rect 51816 153342 51868 153348
rect 51828 146810 51856 153342
rect 51920 153202 51948 460294
rect 51908 153196 51960 153202
rect 51908 153138 51960 153144
rect 52012 152590 52040 463354
rect 52104 154358 52132 466210
rect 52182 466032 52238 466041
rect 52182 465967 52238 465976
rect 52092 154352 52144 154358
rect 52092 154294 52144 154300
rect 52196 154154 52224 465967
rect 53104 465928 53156 465934
rect 53104 465870 53156 465876
rect 53012 463140 53064 463146
rect 53012 463082 53064 463088
rect 52828 463004 52880 463010
rect 52828 462946 52880 462952
rect 52276 460692 52328 460698
rect 52276 460634 52328 460640
rect 52288 459649 52316 460634
rect 52368 460488 52420 460494
rect 52368 460430 52420 460436
rect 52274 459640 52330 459649
rect 52274 459575 52330 459584
rect 52276 458924 52328 458930
rect 52276 458866 52328 458872
rect 52288 373794 52316 458866
rect 52276 373788 52328 373794
rect 52276 373730 52328 373736
rect 52274 372736 52330 372745
rect 52274 372671 52330 372680
rect 52184 154148 52236 154154
rect 52184 154090 52236 154096
rect 52184 154012 52236 154018
rect 52184 153954 52236 153960
rect 52196 153270 52224 153954
rect 52184 153264 52236 153270
rect 52184 153206 52236 153212
rect 52000 152584 52052 152590
rect 52000 152526 52052 152532
rect 51908 151088 51960 151094
rect 51908 151030 51960 151036
rect 51816 146804 51868 146810
rect 51816 146746 51868 146752
rect 51920 142154 51948 151030
rect 52196 147082 52224 153206
rect 52184 147076 52236 147082
rect 52184 147018 52236 147024
rect 52092 146872 52144 146878
rect 52092 146814 52144 146820
rect 51920 142126 52040 142154
rect 51908 133476 51960 133482
rect 51908 133418 51960 133424
rect 51724 130892 51776 130898
rect 51724 130834 51776 130840
rect 51632 130348 51684 130354
rect 51632 130290 51684 130296
rect 51448 44192 51500 44198
rect 51448 44134 51500 44140
rect 50988 42764 51040 42770
rect 50988 42706 51040 42712
rect 50160 42152 50212 42158
rect 50160 42094 50212 42100
rect 51644 40730 51672 130290
rect 51736 41002 51764 130834
rect 51724 40996 51776 41002
rect 51724 40938 51776 40944
rect 51632 40724 51684 40730
rect 51632 40666 51684 40672
rect 44088 39772 44140 39778
rect 44088 39714 44140 39720
rect 51920 39370 51948 133418
rect 52012 39982 52040 142126
rect 52104 41410 52132 146814
rect 52184 146804 52236 146810
rect 52184 146746 52236 146752
rect 52092 41404 52144 41410
rect 52092 41346 52144 41352
rect 52000 39976 52052 39982
rect 52000 39918 52052 39924
rect 52196 39914 52224 146746
rect 52288 42702 52316 372671
rect 52276 42696 52328 42702
rect 52276 42638 52328 42644
rect 52380 42430 52408 460430
rect 52736 459128 52788 459134
rect 52736 459070 52788 459076
rect 52748 451274 52776 459070
rect 52840 457722 52868 462946
rect 53024 457842 53052 463082
rect 53012 457836 53064 457842
rect 53012 457778 53064 457784
rect 52840 457694 53052 457722
rect 52748 451246 52960 451274
rect 52932 372230 52960 451246
rect 52920 372224 52972 372230
rect 52920 372166 52972 372172
rect 52920 370524 52972 370530
rect 52920 370466 52972 370472
rect 52932 320142 52960 370466
rect 52920 320136 52972 320142
rect 52920 320078 52972 320084
rect 52918 319968 52974 319977
rect 52918 319903 52974 319912
rect 52828 260908 52880 260914
rect 52828 260850 52880 260856
rect 52840 151298 52868 260850
rect 52932 260302 52960 319903
rect 53024 263294 53052 457694
rect 53116 263430 53144 465870
rect 53104 263424 53156 263430
rect 53104 263366 53156 263372
rect 53012 263288 53064 263294
rect 53012 263230 53064 263236
rect 53208 260574 53236 487086
rect 53288 487076 53340 487082
rect 53288 487018 53340 487024
rect 53196 260568 53248 260574
rect 53196 260510 53248 260516
rect 52920 260296 52972 260302
rect 52920 260238 52972 260244
rect 53300 260098 53328 487018
rect 53392 263226 53420 492118
rect 55036 491904 55088 491910
rect 55036 491846 55088 491852
rect 53748 491836 53800 491842
rect 53748 491778 53800 491784
rect 53562 466304 53618 466313
rect 53562 466239 53618 466248
rect 53472 460760 53524 460766
rect 53472 460702 53524 460708
rect 53484 459649 53512 460702
rect 53470 459640 53526 459649
rect 53470 459575 53526 459584
rect 53472 457836 53524 457842
rect 53472 457778 53524 457784
rect 53380 263220 53432 263226
rect 53380 263162 53432 263168
rect 53288 260092 53340 260098
rect 53288 260034 53340 260040
rect 53300 258074 53328 260034
rect 53300 258046 53420 258074
rect 53012 241528 53064 241534
rect 53012 241470 53064 241476
rect 52828 151292 52880 151298
rect 52828 151234 52880 151240
rect 53024 130937 53052 241470
rect 53104 240100 53156 240106
rect 53104 240042 53156 240048
rect 53116 239834 53144 240042
rect 53104 239828 53156 239834
rect 53104 239770 53156 239776
rect 53116 151434 53144 239770
rect 53104 151428 53156 151434
rect 53104 151370 53156 151376
rect 53288 133204 53340 133210
rect 53288 133146 53340 133152
rect 53010 130928 53066 130937
rect 53010 130863 53066 130872
rect 53300 43654 53328 133146
rect 53392 130830 53420 258046
rect 53484 152658 53512 457778
rect 53576 154290 53604 466239
rect 53654 466168 53710 466177
rect 53654 466103 53710 466112
rect 53564 154284 53616 154290
rect 53564 154226 53616 154232
rect 53472 152652 53524 152658
rect 53472 152594 53524 152600
rect 53668 151706 53696 466103
rect 53656 151700 53708 151706
rect 53656 151642 53708 151648
rect 53656 133816 53708 133822
rect 53656 133758 53708 133764
rect 53472 133748 53524 133754
rect 53472 133690 53524 133696
rect 53380 130824 53432 130830
rect 53380 130766 53432 130772
rect 53288 43648 53340 43654
rect 53288 43590 53340 43596
rect 52368 42424 52420 42430
rect 52368 42366 52420 42372
rect 53392 40934 53420 130766
rect 53380 40928 53432 40934
rect 53380 40870 53432 40876
rect 53484 40662 53512 133690
rect 53668 133414 53696 133758
rect 53656 133408 53708 133414
rect 53656 133350 53708 133356
rect 53564 133272 53616 133278
rect 53564 133214 53616 133220
rect 53576 41274 53604 133214
rect 53564 41268 53616 41274
rect 53564 41210 53616 41216
rect 53472 40656 53524 40662
rect 53472 40598 53524 40604
rect 52184 39908 52236 39914
rect 52184 39850 52236 39856
rect 53668 39438 53696 133350
rect 53760 42634 53788 491778
rect 54668 489048 54720 489054
rect 54668 488990 54720 488996
rect 54392 486668 54444 486674
rect 54392 486610 54444 486616
rect 54300 459060 54352 459066
rect 54300 459002 54352 459008
rect 54312 373250 54340 459002
rect 54300 373244 54352 373250
rect 54300 373186 54352 373192
rect 54404 373182 54432 486610
rect 54576 465996 54628 466002
rect 54576 465938 54628 465944
rect 54484 416696 54536 416702
rect 54484 416638 54536 416644
rect 54392 373176 54444 373182
rect 54392 373118 54444 373124
rect 54392 372224 54444 372230
rect 54392 372166 54444 372172
rect 54300 320136 54352 320142
rect 54300 320078 54352 320084
rect 54312 271182 54340 320078
rect 54300 271176 54352 271182
rect 54300 271118 54352 271124
rect 54300 260296 54352 260302
rect 54300 260238 54352 260244
rect 53840 239692 53892 239698
rect 53840 239634 53892 239640
rect 53852 238542 53880 239634
rect 53840 238536 53892 238542
rect 53840 238478 53892 238484
rect 53852 237454 53880 238478
rect 53840 237448 53892 237454
rect 53840 237390 53892 237396
rect 54208 130280 54260 130286
rect 54208 130222 54260 130228
rect 54220 44538 54248 130222
rect 54312 129577 54340 260238
rect 54404 260030 54432 372166
rect 54496 263566 54524 416638
rect 54484 263560 54536 263566
rect 54484 263502 54536 263508
rect 54588 263362 54616 465938
rect 54576 263356 54628 263362
rect 54576 263298 54628 263304
rect 54680 262682 54708 488990
rect 54944 463616 54996 463622
rect 54944 463558 54996 463564
rect 54852 463276 54904 463282
rect 54852 463218 54904 463224
rect 54760 463208 54812 463214
rect 54760 463150 54812 463156
rect 54668 262676 54720 262682
rect 54668 262618 54720 262624
rect 54576 260568 54628 260574
rect 54576 260510 54628 260516
rect 54392 260024 54444 260030
rect 54392 259966 54444 259972
rect 54392 241596 54444 241602
rect 54392 241538 54444 241544
rect 54404 151638 54432 241538
rect 54484 237448 54536 237454
rect 54484 237390 54536 237396
rect 54392 151632 54444 151638
rect 54392 151574 54444 151580
rect 54496 133890 54524 237390
rect 54484 133884 54536 133890
rect 54484 133826 54536 133832
rect 54496 133550 54524 133826
rect 54484 133544 54536 133550
rect 54484 133486 54536 133492
rect 54484 130552 54536 130558
rect 54484 130494 54536 130500
rect 54496 129742 54524 130494
rect 54588 129742 54616 260510
rect 54772 152862 54800 463150
rect 54864 152998 54892 463218
rect 54852 152992 54904 152998
rect 54852 152934 54904 152940
rect 54760 152856 54812 152862
rect 54760 152798 54812 152804
rect 54956 152726 54984 463558
rect 54944 152720 54996 152726
rect 54944 152662 54996 152668
rect 55048 152318 55076 491846
rect 55772 488980 55824 488986
rect 55772 488922 55824 488928
rect 55496 460624 55548 460630
rect 55496 460566 55548 460572
rect 55128 460556 55180 460562
rect 55128 460498 55180 460504
rect 55036 152312 55088 152318
rect 55036 152254 55088 152260
rect 54944 151632 54996 151638
rect 54944 151574 54996 151580
rect 54852 151292 54904 151298
rect 54852 151234 54904 151240
rect 54760 133544 54812 133550
rect 54760 133486 54812 133492
rect 54668 130212 54720 130218
rect 54668 130154 54720 130160
rect 54484 129736 54536 129742
rect 54390 129704 54446 129713
rect 54484 129678 54536 129684
rect 54576 129736 54628 129742
rect 54576 129678 54628 129684
rect 54390 129639 54446 129648
rect 54298 129568 54354 129577
rect 54298 129503 54354 129512
rect 54208 44532 54260 44538
rect 54208 44474 54260 44480
rect 54404 44266 54432 129639
rect 54392 44260 54444 44266
rect 54392 44202 54444 44208
rect 54496 44062 54524 129678
rect 54484 44056 54536 44062
rect 54484 43998 54536 44004
rect 53748 42628 53800 42634
rect 53748 42570 53800 42576
rect 54680 42090 54708 130154
rect 54668 42084 54720 42090
rect 54668 42026 54720 42032
rect 54772 40050 54800 133486
rect 54864 44334 54892 151234
rect 54852 44328 54904 44334
rect 54852 44270 54904 44276
rect 54956 43858 54984 151574
rect 55036 151156 55088 151162
rect 55036 151098 55088 151104
rect 54944 43852 54996 43858
rect 54944 43794 54996 43800
rect 54760 40044 54812 40050
rect 54760 39986 54812 39992
rect 55048 39846 55076 151098
rect 55140 42498 55168 460498
rect 55508 459649 55536 460566
rect 55494 459640 55550 459649
rect 55494 459575 55550 459584
rect 55680 411120 55732 411126
rect 55680 411062 55732 411068
rect 55692 373454 55720 411062
rect 55680 373448 55732 373454
rect 55680 373390 55732 373396
rect 55784 262750 55812 488922
rect 55956 463480 56008 463486
rect 55956 463422 56008 463428
rect 55864 462868 55916 462874
rect 55864 462810 55916 462816
rect 55772 262744 55824 262750
rect 55772 262686 55824 262692
rect 55772 260500 55824 260506
rect 55772 260442 55824 260448
rect 55784 259350 55812 260442
rect 55772 259344 55824 259350
rect 55772 259286 55824 259292
rect 55680 239964 55732 239970
rect 55680 239906 55732 239912
rect 55692 151774 55720 239906
rect 55680 151768 55732 151774
rect 55680 151710 55732 151716
rect 55784 131102 55812 259286
rect 55876 152522 55904 462810
rect 55968 153066 55996 463422
rect 56232 463344 56284 463350
rect 56232 463286 56284 463292
rect 56048 462936 56100 462942
rect 56048 462878 56100 462884
rect 55956 153060 56008 153066
rect 55956 153002 56008 153008
rect 56060 152794 56088 462878
rect 56244 460934 56272 463286
rect 56152 460906 56272 460934
rect 56152 153134 56180 460906
rect 56232 458992 56284 458998
rect 56232 458934 56284 458940
rect 56244 415410 56272 458934
rect 56232 415404 56284 415410
rect 56232 415346 56284 415352
rect 56232 408604 56284 408610
rect 56232 408546 56284 408552
rect 56244 373726 56272 408546
rect 56232 373720 56284 373726
rect 56232 373662 56284 373668
rect 56230 372736 56286 372745
rect 56230 372671 56286 372680
rect 56140 153128 56192 153134
rect 56140 153070 56192 153076
rect 56048 152788 56100 152794
rect 56048 152730 56100 152736
rect 55864 152516 55916 152522
rect 55864 152458 55916 152464
rect 55772 131096 55824 131102
rect 55772 131038 55824 131044
rect 56046 131064 56102 131073
rect 56046 130999 56102 131008
rect 55956 130756 56008 130762
rect 55956 130698 56008 130704
rect 55968 130626 55996 130698
rect 55956 130620 56008 130626
rect 55956 130562 56008 130568
rect 55864 130484 55916 130490
rect 55864 130426 55916 130432
rect 55876 129742 55904 130426
rect 55864 129736 55916 129742
rect 55864 129678 55916 129684
rect 55128 42492 55180 42498
rect 55128 42434 55180 42440
rect 55876 40798 55904 129678
rect 55968 44470 55996 130562
rect 55956 44464 56008 44470
rect 55956 44406 56008 44412
rect 56060 43790 56088 130999
rect 56138 130928 56194 130937
rect 56138 130863 56194 130872
rect 56152 130529 56180 130863
rect 56138 130520 56194 130529
rect 56138 130455 56194 130464
rect 56048 43784 56100 43790
rect 56048 43726 56100 43732
rect 56152 42226 56180 130455
rect 56244 43518 56272 372671
rect 56336 154222 56364 493342
rect 59268 492652 59320 492658
rect 59268 492594 59320 492600
rect 56416 492312 56468 492318
rect 56416 492254 56468 492260
rect 56324 154216 56376 154222
rect 56324 154158 56376 154164
rect 56428 152930 56456 492254
rect 57244 492244 57296 492250
rect 57244 492186 57296 492192
rect 56508 491700 56560 491706
rect 56508 491642 56560 491648
rect 56416 152924 56468 152930
rect 56416 152866 56468 152872
rect 56324 133816 56376 133822
rect 56324 133758 56376 133764
rect 56336 43722 56364 133758
rect 56416 131096 56468 131102
rect 56416 131038 56468 131044
rect 56428 130966 56456 131038
rect 56416 130960 56468 130966
rect 56416 130902 56468 130908
rect 56324 43716 56376 43722
rect 56324 43658 56376 43664
rect 56232 43512 56284 43518
rect 56232 43454 56284 43460
rect 56140 42220 56192 42226
rect 56140 42162 56192 42168
rect 55864 40792 55916 40798
rect 55864 40734 55916 40740
rect 55036 39840 55088 39846
rect 55036 39782 55088 39788
rect 56428 39574 56456 130902
rect 56520 42566 56548 491642
rect 57152 489320 57204 489326
rect 57152 489262 57204 489268
rect 57060 484356 57112 484362
rect 57060 484298 57112 484304
rect 56600 415404 56652 415410
rect 56600 415346 56652 415352
rect 56612 408610 56640 415346
rect 57072 408610 57100 484298
rect 56600 408604 56652 408610
rect 56600 408546 56652 408552
rect 57060 408604 57112 408610
rect 57060 408546 57112 408552
rect 57060 407516 57112 407522
rect 57060 407458 57112 407464
rect 56876 383648 56928 383654
rect 56876 383590 56928 383596
rect 56888 383081 56916 383590
rect 56874 383072 56930 383081
rect 56874 383007 56930 383016
rect 56968 382356 57020 382362
rect 56968 382298 57020 382304
rect 56980 374066 57008 382298
rect 56968 374060 57020 374066
rect 56968 374002 57020 374008
rect 57072 373658 57100 407458
rect 57164 383654 57192 489262
rect 57256 416702 57284 492186
rect 58992 490612 59044 490618
rect 58992 490554 59044 490560
rect 57704 487824 57756 487830
rect 57704 487766 57756 487772
rect 57612 482316 57664 482322
rect 57612 482258 57664 482264
rect 57520 467152 57572 467158
rect 57520 467094 57572 467100
rect 57428 465860 57480 465866
rect 57428 465802 57480 465808
rect 57336 461780 57388 461786
rect 57336 461722 57388 461728
rect 57244 416696 57296 416702
rect 57244 416638 57296 416644
rect 57244 412616 57296 412622
rect 57244 412558 57296 412564
rect 57256 412457 57284 412558
rect 57242 412448 57298 412457
rect 57242 412383 57298 412392
rect 57244 411256 57296 411262
rect 57242 411224 57244 411233
rect 57296 411224 57298 411233
rect 57242 411159 57298 411168
rect 57242 408640 57298 408649
rect 57242 408575 57298 408584
rect 57256 408542 57284 408575
rect 57244 408536 57296 408542
rect 57244 408478 57296 408484
rect 57242 407280 57298 407289
rect 57242 407215 57298 407224
rect 57256 407182 57284 407215
rect 57244 407176 57296 407182
rect 57244 407118 57296 407124
rect 57242 405784 57298 405793
rect 57242 405719 57244 405728
rect 57296 405719 57298 405728
rect 57244 405690 57296 405696
rect 57242 404424 57298 404433
rect 57242 404359 57244 404368
rect 57296 404359 57298 404368
rect 57244 404330 57296 404336
rect 57242 403064 57298 403073
rect 57242 402999 57244 403008
rect 57296 402999 57298 403008
rect 57244 402970 57296 402976
rect 57244 385008 57296 385014
rect 57242 384976 57244 384985
rect 57296 384976 57298 384985
rect 57242 384911 57298 384920
rect 57164 383626 57284 383654
rect 57152 383580 57204 383586
rect 57152 383522 57204 383528
rect 57164 377806 57192 383522
rect 57256 382362 57284 383626
rect 57244 382356 57296 382362
rect 57244 382298 57296 382304
rect 57244 382220 57296 382226
rect 57244 382162 57296 382168
rect 57152 377800 57204 377806
rect 57152 377742 57204 377748
rect 57060 373652 57112 373658
rect 57060 373594 57112 373600
rect 57152 346928 57204 346934
rect 57152 346870 57204 346876
rect 56782 301744 56838 301753
rect 56782 301679 56838 301688
rect 56598 300928 56654 300937
rect 56598 300863 56654 300872
rect 56612 191729 56640 300863
rect 56690 293992 56746 294001
rect 56690 293927 56746 293936
rect 56598 191720 56654 191729
rect 56598 191655 56654 191664
rect 56704 185473 56732 293927
rect 56796 193225 56824 301679
rect 57060 292528 57112 292534
rect 57060 292470 57112 292476
rect 56876 291916 56928 291922
rect 56876 291858 56928 291864
rect 56888 264217 56916 291858
rect 56874 264208 56930 264217
rect 56874 264143 56930 264152
rect 56968 236020 57020 236026
rect 56968 235962 57020 235968
rect 56782 193216 56838 193225
rect 56782 193151 56838 193160
rect 56782 191720 56838 191729
rect 56782 191655 56838 191664
rect 56796 190913 56824 191655
rect 56782 190904 56838 190913
rect 56782 190839 56838 190848
rect 56690 185464 56746 185473
rect 56690 185399 56746 185408
rect 56796 81433 56824 190839
rect 56874 187912 56930 187921
rect 56874 187847 56930 187856
rect 56782 81424 56838 81433
rect 56782 81359 56838 81368
rect 56888 78441 56916 187847
rect 56980 154562 57008 235962
rect 57072 183569 57100 292470
rect 57164 292262 57192 346870
rect 57152 292256 57204 292262
rect 57152 292198 57204 292204
rect 57256 273329 57284 382162
rect 57348 294953 57376 461722
rect 57440 297809 57468 465802
rect 57532 383466 57560 467094
rect 57624 383586 57652 482258
rect 57612 383580 57664 383586
rect 57612 383522 57664 383528
rect 57532 383438 57652 383466
rect 57518 383344 57574 383353
rect 57518 383279 57574 383288
rect 57532 382226 57560 383279
rect 57520 382220 57572 382226
rect 57520 382162 57572 382168
rect 57624 377890 57652 383438
rect 57532 377862 57652 377890
rect 57426 297800 57482 297809
rect 57426 297735 57482 297744
rect 57334 294944 57390 294953
rect 57334 294879 57390 294888
rect 57348 294001 57376 294879
rect 57334 293992 57390 294001
rect 57334 293927 57390 293936
rect 57334 292632 57390 292641
rect 57334 292567 57390 292576
rect 57348 292534 57376 292567
rect 57336 292528 57388 292534
rect 57336 292470 57388 292476
rect 57242 273320 57298 273329
rect 57242 273255 57298 273264
rect 57152 239760 57204 239766
rect 57152 239702 57204 239708
rect 57164 238474 57192 239702
rect 57244 239284 57296 239290
rect 57244 239226 57296 239232
rect 57152 238468 57204 238474
rect 57152 238410 57204 238416
rect 57164 237425 57192 238410
rect 57150 237416 57206 237425
rect 57150 237351 57206 237360
rect 57150 185736 57206 185745
rect 57150 185671 57206 185680
rect 57058 183560 57114 183569
rect 57058 183495 57114 183504
rect 56968 154556 57020 154562
rect 56968 154498 57020 154504
rect 57060 151428 57112 151434
rect 57060 151370 57112 151376
rect 56968 133816 57020 133822
rect 56966 133784 56968 133793
rect 57020 133784 57022 133793
rect 56966 133719 57022 133728
rect 56968 131096 57020 131102
rect 56968 131038 57020 131044
rect 56874 78432 56930 78441
rect 56874 78367 56930 78376
rect 56508 42560 56560 42566
rect 56508 42502 56560 42508
rect 56980 39710 57008 131038
rect 57072 43926 57100 151370
rect 57164 76673 57192 185671
rect 57256 131102 57284 239226
rect 57440 187921 57468 297735
rect 57532 296041 57560 377862
rect 57612 377800 57664 377806
rect 57612 377742 57664 377748
rect 57624 301753 57652 377742
rect 57610 301744 57666 301753
rect 57610 301679 57666 301688
rect 57716 300937 57744 487766
rect 58624 487008 58676 487014
rect 58624 486950 58676 486956
rect 57888 486260 57940 486266
rect 57888 486202 57940 486208
rect 57796 466064 57848 466070
rect 57796 466006 57848 466012
rect 57702 300928 57758 300937
rect 57702 300863 57758 300872
rect 57702 299432 57758 299441
rect 57702 299367 57758 299376
rect 57518 296032 57574 296041
rect 57518 295967 57574 295976
rect 57426 187912 57482 187921
rect 57426 187847 57482 187856
rect 57334 187776 57390 187785
rect 57334 187711 57390 187720
rect 57244 131096 57296 131102
rect 57244 131038 57296 131044
rect 57348 79393 57376 187711
rect 57532 185745 57560 295967
rect 57612 276004 57664 276010
rect 57612 275946 57664 275952
rect 57624 275641 57652 275946
rect 57610 275632 57666 275641
rect 57610 275567 57666 275576
rect 57610 193216 57666 193225
rect 57610 193151 57666 193160
rect 57624 191865 57652 193151
rect 57610 191856 57666 191865
rect 57610 191791 57666 191800
rect 57518 185736 57574 185745
rect 57518 185671 57574 185680
rect 57426 183560 57482 183569
rect 57426 183495 57482 183504
rect 57334 79384 57390 79393
rect 57334 79319 57390 79328
rect 57150 76664 57206 76673
rect 57150 76599 57206 76608
rect 57440 73817 57468 183495
rect 57624 82521 57652 191791
rect 57716 188737 57744 299367
rect 57808 263498 57836 466006
rect 57900 299441 57928 486202
rect 58532 483608 58584 483614
rect 58532 483550 58584 483556
rect 57980 408604 58032 408610
rect 57980 408546 58032 408552
rect 57886 299432 57942 299441
rect 57886 299367 57942 299376
rect 57992 291922 58020 408546
rect 58544 407794 58572 483550
rect 58532 407788 58584 407794
rect 58532 407730 58584 407736
rect 58636 370530 58664 486950
rect 58900 486396 58952 486402
rect 58900 486338 58952 486344
rect 58808 486328 58860 486334
rect 58808 486270 58860 486276
rect 58716 484288 58768 484294
rect 58716 484230 58768 484236
rect 58728 373930 58756 484230
rect 58820 374950 58848 486270
rect 58808 374944 58860 374950
rect 58808 374886 58860 374892
rect 58912 374882 58940 486338
rect 58900 374876 58952 374882
rect 58900 374818 58952 374824
rect 58716 373924 58768 373930
rect 58716 373866 58768 373872
rect 58624 370524 58676 370530
rect 58624 370466 58676 370472
rect 58624 349104 58676 349110
rect 58624 349046 58676 349052
rect 57980 291916 58032 291922
rect 57980 291858 58032 291864
rect 57886 273320 57942 273329
rect 57886 273255 57942 273264
rect 57796 263492 57848 263498
rect 57796 263434 57848 263440
rect 57702 188728 57758 188737
rect 57702 188663 57758 188672
rect 57716 187785 57744 188663
rect 57702 187776 57758 187785
rect 57702 187711 57758 187720
rect 57702 185464 57758 185473
rect 57702 185399 57758 185408
rect 57610 82512 57666 82521
rect 57610 82447 57666 82456
rect 57716 75585 57744 185399
rect 57900 163305 57928 273255
rect 57980 271176 58032 271182
rect 57980 271118 58032 271124
rect 57992 260914 58020 271118
rect 58636 264994 58664 349046
rect 58900 348696 58952 348702
rect 58900 348638 58952 348644
rect 58624 264988 58676 264994
rect 58624 264930 58676 264936
rect 58636 264897 58664 264930
rect 58622 264888 58678 264897
rect 58622 264823 58678 264832
rect 58912 263702 58940 348638
rect 59004 273057 59032 490554
rect 59084 463072 59136 463078
rect 59084 463014 59136 463020
rect 58990 273048 59046 273057
rect 58990 272983 59046 272992
rect 58900 263696 58952 263702
rect 58900 263638 58952 263644
rect 57980 260908 58032 260914
rect 57980 260850 58032 260856
rect 57980 260364 58032 260370
rect 57980 260306 58032 260312
rect 57992 259418 58020 260306
rect 57980 259412 58032 259418
rect 57980 259354 58032 259360
rect 57886 163296 57942 163305
rect 57886 163231 57942 163240
rect 57796 151768 57848 151774
rect 57796 151710 57848 151716
rect 57808 150521 57836 151710
rect 57794 150512 57850 150521
rect 57794 150447 57850 150456
rect 57796 81456 57848 81462
rect 57796 81398 57848 81404
rect 57702 75576 57758 75585
rect 57702 75511 57758 75520
rect 57426 73808 57482 73817
rect 57426 73743 57482 73752
rect 57060 43920 57112 43926
rect 57060 43862 57112 43868
rect 57244 42832 57296 42838
rect 57244 42774 57296 42780
rect 56968 39704 57020 39710
rect 56968 39646 57020 39652
rect 56416 39568 56468 39574
rect 56416 39510 56468 39516
rect 53656 39432 53708 39438
rect 53656 39374 53708 39380
rect 51908 39364 51960 39370
rect 51908 39306 51960 39312
rect 2780 31748 2832 31754
rect 2780 31690 2832 31696
rect 2792 31385 2820 31690
rect 2778 31376 2834 31385
rect 2778 31311 2834 31320
rect 2792 3534 2820 31311
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 57256 3466 57284 42774
rect 57808 41342 57836 81398
rect 57900 53417 57928 163231
rect 57992 131073 58020 259354
rect 58992 240100 59044 240106
rect 58992 240042 59044 240048
rect 58808 240032 58860 240038
rect 58808 239974 58860 239980
rect 58622 237416 58678 237425
rect 58622 237351 58678 237360
rect 58636 150686 58664 237351
rect 58820 229094 58848 239974
rect 58900 239556 58952 239562
rect 58900 239498 58952 239504
rect 58912 238649 58940 239498
rect 58898 238640 58954 238649
rect 58898 238575 58954 238584
rect 58912 237425 58940 238575
rect 58898 237416 58954 237425
rect 58898 237351 58954 237360
rect 58820 229066 58940 229094
rect 58624 150680 58676 150686
rect 58624 150622 58676 150628
rect 58624 150408 58676 150414
rect 58624 150350 58676 150356
rect 57978 131064 58034 131073
rect 57978 130999 58034 131008
rect 57886 53408 57942 53417
rect 57886 53343 57942 53352
rect 57900 44130 57928 53343
rect 57888 44124 57940 44130
rect 57888 44066 57940 44072
rect 57900 42838 57928 44066
rect 57888 42832 57940 42838
rect 57888 42774 57940 42780
rect 57796 41336 57848 41342
rect 57796 41278 57848 41284
rect 58636 41138 58664 150350
rect 58912 130694 58940 229066
rect 59004 151814 59032 240042
rect 59096 165617 59124 463014
rect 59176 459264 59228 459270
rect 59176 459206 59228 459212
rect 59082 165608 59138 165617
rect 59082 165543 59138 165552
rect 59188 153882 59216 459206
rect 59280 154086 59308 492594
rect 60108 492590 60136 495094
rect 60292 495023 60582 495051
rect 60844 495023 61042 495051
rect 61120 495023 61502 495051
rect 61978 495023 62068 495051
rect 60096 492584 60148 492590
rect 60096 492526 60148 492532
rect 60292 489914 60320 495023
rect 60740 490340 60792 490346
rect 60740 490282 60792 490288
rect 59372 489886 60320 489914
rect 59372 483546 59400 489886
rect 59820 489796 59872 489802
rect 59820 489738 59872 489744
rect 59728 486940 59780 486946
rect 59728 486882 59780 486888
rect 59636 484152 59688 484158
rect 59636 484094 59688 484100
rect 59360 483540 59412 483546
rect 59360 483482 59412 483488
rect 59360 407788 59412 407794
rect 59360 407730 59412 407736
rect 59372 346934 59400 407730
rect 59648 407522 59676 484094
rect 59636 407516 59688 407522
rect 59636 407458 59688 407464
rect 59740 373114 59768 486882
rect 59728 373108 59780 373114
rect 59728 373050 59780 373056
rect 59360 346928 59412 346934
rect 59360 346870 59412 346876
rect 59728 292256 59780 292262
rect 59728 292198 59780 292204
rect 59740 260846 59768 292198
rect 59832 262721 59860 489738
rect 60002 465896 60058 465905
rect 60002 465831 60058 465840
rect 59912 463684 59964 463690
rect 59912 463626 59964 463632
rect 59818 262712 59874 262721
rect 59818 262647 59874 262656
rect 59728 260840 59780 260846
rect 59728 260782 59780 260788
rect 59740 236026 59768 260782
rect 59728 236020 59780 236026
rect 59728 235962 59780 235968
rect 59360 154556 59412 154562
rect 59360 154498 59412 154504
rect 59268 154080 59320 154086
rect 59268 154022 59320 154028
rect 59176 153876 59228 153882
rect 59176 153818 59228 153824
rect 59372 153338 59400 154498
rect 59360 153332 59412 153338
rect 59360 153274 59412 153280
rect 59004 151786 59124 151814
rect 59096 130762 59124 151786
rect 59268 151224 59320 151230
rect 59268 151166 59320 151172
rect 59280 150414 59308 151166
rect 59268 150408 59320 150414
rect 59268 150350 59320 150356
rect 59084 130756 59136 130762
rect 59084 130698 59136 130704
rect 58900 130688 58952 130694
rect 58900 130630 58952 130636
rect 58990 130656 59046 130665
rect 58990 130591 59046 130600
rect 59004 44402 59032 130591
rect 58992 44396 59044 44402
rect 58992 44338 59044 44344
rect 58624 41132 58676 41138
rect 58624 41074 58676 41080
rect 59096 40866 59124 130698
rect 59268 130688 59320 130694
rect 59268 130630 59320 130636
rect 59176 130416 59228 130422
rect 59176 130358 59228 130364
rect 59084 40860 59136 40866
rect 59084 40802 59136 40808
rect 59188 39642 59216 130358
rect 59176 39636 59228 39642
rect 59176 39578 59228 39584
rect 59280 39506 59308 130630
rect 59372 81462 59400 153274
rect 59832 131102 59860 262647
rect 59924 154018 59952 463626
rect 59912 154012 59964 154018
rect 59912 153954 59964 153960
rect 60016 153950 60044 465831
rect 60752 458862 60780 490282
rect 60844 480962 60872 495023
rect 61120 490346 61148 495023
rect 61936 492584 61988 492590
rect 61936 492526 61988 492532
rect 61108 490340 61160 490346
rect 61108 490282 61160 490288
rect 61948 489190 61976 492526
rect 62040 492386 62068 495023
rect 62224 495023 62330 495051
rect 62806 495023 62896 495051
rect 62120 492584 62172 492590
rect 62120 492526 62172 492532
rect 62028 492380 62080 492386
rect 62028 492322 62080 492328
rect 61936 489184 61988 489190
rect 61936 489126 61988 489132
rect 60832 480956 60884 480962
rect 60832 480898 60884 480904
rect 62132 460086 62160 492526
rect 62224 461718 62252 495023
rect 62764 492380 62816 492386
rect 62764 492322 62816 492328
rect 62776 475386 62804 492322
rect 62868 492046 62896 495023
rect 62960 495023 63250 495051
rect 63512 495023 63710 495051
rect 63788 495023 64170 495051
rect 64248 495023 64538 495051
rect 62960 492590 62988 495023
rect 62948 492584 63000 492590
rect 62948 492526 63000 492532
rect 63040 492584 63092 492590
rect 63040 492526 63092 492532
rect 63052 492318 63080 492526
rect 63040 492312 63092 492318
rect 63040 492254 63092 492260
rect 62856 492040 62908 492046
rect 62856 491982 62908 491988
rect 62764 475380 62816 475386
rect 62764 475322 62816 475328
rect 62212 461712 62264 461718
rect 62212 461654 62264 461660
rect 63512 460222 63540 495023
rect 63788 492538 63816 495023
rect 63604 492510 63816 492538
rect 63604 460222 63632 492510
rect 64248 489914 64276 495023
rect 64880 492380 64932 492386
rect 64880 492322 64932 492328
rect 63696 489886 64276 489914
rect 63696 462806 63724 489886
rect 64892 465526 64920 492322
rect 64984 465594 65012 495037
rect 65076 495023 65458 495051
rect 65536 495023 65918 495051
rect 66272 495023 66378 495051
rect 66456 495023 66746 495051
rect 66824 495023 67206 495051
rect 67682 495023 67864 495051
rect 65076 465662 65104 495023
rect 65536 492386 65564 495023
rect 66272 492674 66300 495023
rect 66180 492646 66300 492674
rect 65524 492380 65576 492386
rect 65524 492322 65576 492328
rect 66180 492289 66208 492646
rect 66456 492538 66484 495023
rect 66272 492510 66484 492538
rect 66166 492280 66222 492289
rect 66166 492215 66222 492224
rect 65064 465656 65116 465662
rect 65064 465598 65116 465604
rect 64972 465588 65024 465594
rect 64972 465530 65024 465536
rect 64880 465520 64932 465526
rect 64880 465462 64932 465468
rect 63684 462800 63736 462806
rect 63684 462742 63736 462748
rect 63500 460216 63552 460222
rect 63500 460158 63552 460164
rect 63592 460216 63644 460222
rect 63592 460158 63644 460164
rect 66272 460154 66300 492510
rect 66824 489914 66852 495023
rect 67732 492448 67784 492454
rect 67732 492390 67784 492396
rect 67640 492380 67692 492386
rect 67640 492322 67692 492328
rect 66364 489886 66852 489914
rect 66364 468450 66392 489886
rect 66352 468444 66404 468450
rect 66352 468386 66404 468392
rect 67652 460426 67680 492322
rect 67640 460420 67692 460426
rect 67640 460362 67692 460368
rect 66260 460148 66312 460154
rect 66260 460090 66312 460096
rect 62120 460080 62172 460086
rect 67744 460057 67772 492390
rect 67836 469130 67864 495023
rect 67928 495023 68126 495051
rect 68204 495023 68494 495051
rect 68664 495023 68954 495051
rect 69032 495023 69414 495051
rect 69584 495023 69874 495051
rect 69952 495023 70334 495051
rect 70504 495023 70702 495051
rect 70872 495023 71162 495051
rect 71240 495023 71622 495051
rect 71884 495023 72082 495051
rect 72160 495023 72542 495051
rect 67928 492386 67956 495023
rect 68204 492454 68232 495023
rect 68192 492448 68244 492454
rect 68192 492390 68244 492396
rect 68284 492448 68336 492454
rect 68284 492390 68336 492396
rect 67916 492380 67968 492386
rect 67916 492322 67968 492328
rect 67824 469124 67876 469130
rect 67824 469066 67876 469072
rect 68296 466410 68324 492390
rect 68376 492380 68428 492386
rect 68376 492322 68428 492328
rect 68284 466404 68336 466410
rect 68284 466346 68336 466352
rect 68388 466342 68416 492322
rect 68664 491745 68692 495023
rect 68928 492312 68980 492318
rect 68926 492280 68928 492289
rect 68980 492280 68982 492289
rect 68926 492215 68982 492224
rect 68650 491736 68706 491745
rect 68650 491671 68706 491680
rect 68376 466336 68428 466342
rect 68376 466278 68428 466284
rect 69032 460873 69060 495023
rect 69112 492720 69164 492726
rect 69112 492662 69164 492668
rect 69018 460864 69074 460873
rect 69018 460799 69074 460808
rect 69124 460601 69152 492662
rect 69584 489914 69612 495023
rect 69952 492726 69980 495023
rect 69940 492720 69992 492726
rect 69940 492662 69992 492668
rect 70400 490748 70452 490754
rect 70400 490690 70452 490696
rect 69216 489886 69612 489914
rect 69216 463457 69244 489886
rect 69202 463448 69258 463457
rect 69202 463383 69258 463392
rect 69110 460592 69166 460601
rect 69110 460527 69166 460536
rect 70412 460494 70440 490690
rect 70504 463321 70532 495023
rect 70872 490754 70900 495023
rect 70860 490748 70912 490754
rect 70860 490690 70912 490696
rect 71240 489914 71268 495023
rect 71780 492448 71832 492454
rect 71780 492390 71832 492396
rect 70596 489886 71268 489914
rect 70596 469062 70624 489886
rect 70584 469056 70636 469062
rect 70584 468998 70636 469004
rect 70490 463312 70546 463321
rect 70490 463247 70546 463256
rect 71792 460737 71820 492390
rect 71778 460728 71834 460737
rect 71778 460663 71834 460672
rect 71884 460562 71912 495023
rect 72160 492454 72188 495023
rect 72896 492561 72924 495037
rect 73172 495023 73370 495051
rect 72882 492552 72938 492561
rect 72882 492487 72938 492496
rect 72148 492448 72200 492454
rect 71962 492416 72018 492425
rect 72148 492390 72200 492396
rect 72516 492448 72568 492454
rect 72516 492390 72568 492396
rect 71962 492351 72018 492360
rect 71976 491774 72004 492351
rect 71964 491768 72016 491774
rect 71964 491710 72016 491716
rect 72528 470594 72556 492390
rect 72436 470566 72556 470594
rect 72436 469198 72464 470566
rect 72424 469192 72476 469198
rect 72424 469134 72476 469140
rect 73172 461553 73200 495023
rect 73816 491706 73844 495037
rect 73804 491700 73856 491706
rect 73804 491642 73856 491648
rect 74276 491609 74304 495037
rect 74552 495023 74658 495051
rect 74736 495023 75118 495051
rect 75288 495023 75578 495051
rect 74552 491842 74580 495023
rect 74632 492720 74684 492726
rect 74632 492662 74684 492668
rect 74540 491836 74592 491842
rect 74540 491778 74592 491784
rect 74262 491600 74318 491609
rect 74262 491535 74318 491544
rect 73158 461544 73214 461553
rect 73158 461479 73214 461488
rect 71872 460556 71924 460562
rect 71872 460498 71924 460504
rect 70400 460488 70452 460494
rect 74644 460465 74672 492662
rect 70400 460430 70452 460436
rect 74630 460456 74686 460465
rect 74630 460391 74686 460400
rect 74736 460193 74764 495023
rect 75288 492726 75316 495023
rect 75276 492720 75328 492726
rect 75276 492662 75328 492668
rect 75920 492720 75972 492726
rect 75920 492662 75972 492668
rect 75932 460698 75960 492662
rect 76024 492153 76052 495037
rect 76208 495023 76498 495051
rect 76576 495023 76866 495051
rect 76010 492144 76066 492153
rect 76010 492079 76066 492088
rect 76208 489914 76236 495023
rect 76576 492726 76604 495023
rect 76564 492720 76616 492726
rect 76564 492662 76616 492668
rect 77312 492017 77340 495037
rect 77772 492425 77800 495037
rect 77864 495023 78246 495051
rect 77758 492416 77814 492425
rect 77758 492351 77814 492360
rect 77298 492008 77354 492017
rect 77298 491943 77354 491952
rect 77864 489914 77892 495023
rect 78692 492810 78720 495037
rect 78600 492782 78720 492810
rect 78784 495023 79074 495051
rect 79152 495023 79534 495051
rect 79704 495023 79994 495051
rect 80164 495023 80454 495051
rect 78600 492289 78628 492782
rect 78680 492720 78732 492726
rect 78680 492662 78732 492668
rect 78586 492280 78642 492289
rect 78586 492215 78642 492224
rect 76024 489886 76236 489914
rect 77312 489886 77892 489914
rect 75920 460692 75972 460698
rect 75920 460634 75972 460640
rect 76024 460329 76052 489886
rect 77312 460766 77340 489886
rect 78692 460834 78720 492662
rect 78680 460828 78732 460834
rect 78680 460770 78732 460776
rect 77300 460760 77352 460766
rect 77300 460702 77352 460708
rect 78784 460630 78812 495023
rect 79152 489914 79180 495023
rect 79704 492726 79732 495023
rect 79692 492720 79744 492726
rect 79692 492662 79744 492668
rect 80060 490408 80112 490414
rect 80060 490350 80112 490356
rect 78876 489886 79180 489914
rect 78876 460902 78904 489886
rect 78864 460896 78916 460902
rect 78864 460838 78916 460844
rect 78772 460624 78824 460630
rect 78772 460566 78824 460572
rect 76010 460320 76066 460329
rect 76010 460255 76066 460264
rect 74722 460184 74778 460193
rect 74722 460119 74778 460128
rect 62120 460022 62172 460028
rect 67730 460048 67786 460057
rect 67730 459983 67786 459992
rect 80072 459105 80100 490350
rect 80164 463185 80192 495023
rect 80808 491881 80836 495037
rect 80992 495023 81282 495051
rect 80794 491872 80850 491881
rect 80794 491807 80850 491816
rect 80992 490414 81020 495023
rect 81728 491910 81756 495037
rect 81912 495023 82202 495051
rect 82280 495023 82662 495051
rect 81716 491904 81768 491910
rect 81716 491846 81768 491852
rect 80980 490408 81032 490414
rect 80980 490350 81032 490356
rect 81532 490408 81584 490414
rect 81532 490350 81584 490356
rect 81544 465769 81572 490350
rect 81912 485774 81940 495023
rect 82280 490414 82308 495023
rect 82912 494964 82964 494970
rect 82912 494906 82964 494912
rect 82268 490408 82320 490414
rect 82268 490350 82320 490356
rect 82820 490408 82872 490414
rect 82820 490350 82872 490356
rect 81636 485746 81940 485774
rect 81530 465760 81586 465769
rect 81530 465695 81586 465704
rect 81636 463554 81664 485746
rect 82832 466274 82860 490350
rect 82820 466268 82872 466274
rect 82820 466210 82872 466216
rect 82924 466138 82952 494906
rect 83032 494850 83060 495037
rect 83200 495023 83490 495051
rect 83568 495023 83950 495051
rect 83200 494970 83228 495023
rect 83188 494964 83240 494970
rect 83188 494906 83240 494912
rect 83032 494822 83228 494850
rect 83200 485774 83228 494822
rect 83568 490414 83596 495023
rect 84396 492522 84424 495037
rect 84488 495023 84870 495051
rect 84948 495023 85238 495051
rect 85714 495023 85804 495051
rect 84384 492516 84436 492522
rect 84384 492458 84436 492464
rect 83556 490408 83608 490414
rect 83556 490350 83608 490356
rect 84292 490408 84344 490414
rect 84292 490350 84344 490356
rect 83016 485746 83228 485774
rect 83016 466206 83044 485746
rect 83004 466200 83056 466206
rect 83004 466142 83056 466148
rect 82912 466132 82964 466138
rect 82912 466074 82964 466080
rect 84304 466041 84332 490350
rect 84488 485774 84516 495023
rect 84948 490414 84976 495023
rect 85776 490482 85804 495023
rect 85868 495023 86158 495051
rect 86328 495023 86618 495051
rect 87094 495023 87184 495051
rect 85764 490476 85816 490482
rect 85764 490418 85816 490424
rect 84936 490408 84988 490414
rect 84936 490350 84988 490356
rect 85580 490408 85632 490414
rect 85580 490350 85632 490356
rect 84396 485746 84516 485774
rect 84396 466313 84424 485746
rect 84382 466304 84438 466313
rect 84382 466239 84438 466248
rect 84290 466032 84346 466041
rect 84290 465967 84346 465976
rect 81624 463548 81676 463554
rect 81624 463490 81676 463496
rect 80150 463176 80206 463185
rect 80150 463111 80206 463120
rect 85592 462874 85620 490350
rect 85868 490226 85896 495023
rect 85948 490476 86000 490482
rect 85948 490418 86000 490424
rect 85684 490198 85896 490226
rect 85684 463418 85712 490198
rect 85960 485774 85988 490418
rect 86328 490414 86356 495023
rect 87052 490476 87104 490482
rect 87052 490418 87104 490424
rect 86316 490408 86368 490414
rect 86316 490350 86368 490356
rect 86960 490408 87012 490414
rect 86960 490350 87012 490356
rect 85776 485746 85988 485774
rect 85776 466177 85804 485746
rect 86224 483540 86276 483546
rect 86224 483482 86276 483488
rect 85762 466168 85818 466177
rect 85762 466103 85818 466112
rect 85672 463412 85724 463418
rect 85672 463354 85724 463360
rect 85580 462868 85632 462874
rect 85580 462810 85632 462816
rect 86236 462330 86264 483482
rect 86972 463622 87000 490350
rect 86960 463616 87012 463622
rect 86960 463558 87012 463564
rect 87064 462942 87092 490418
rect 87156 463146 87184 495023
rect 87248 495023 87446 495051
rect 87616 495023 87906 495051
rect 88382 495023 88472 495051
rect 87248 490414 87276 495023
rect 87616 490482 87644 495023
rect 87604 490476 87656 490482
rect 87604 490418 87656 490424
rect 87236 490408 87288 490414
rect 87236 490350 87288 490356
rect 88444 463214 88472 495023
rect 88812 492590 88840 495037
rect 88904 495023 89194 495051
rect 89272 495023 89654 495051
rect 89824 495023 90114 495051
rect 88800 492584 88852 492590
rect 88800 492526 88852 492532
rect 88904 490362 88932 495023
rect 88536 490334 88932 490362
rect 88536 463282 88564 490334
rect 89272 485774 89300 495023
rect 88628 485746 89300 485774
rect 88628 463486 88656 485746
rect 88616 463480 88668 463486
rect 88616 463422 88668 463428
rect 89824 463350 89852 495023
rect 90560 493406 90588 495037
rect 90652 495023 91034 495051
rect 91112 495023 91402 495051
rect 91480 495023 91862 495051
rect 92032 495023 92322 495051
rect 92676 495023 92782 495051
rect 92952 495023 93242 495051
rect 93320 495023 93610 495051
rect 93872 495023 94070 495051
rect 94148 495023 94530 495051
rect 94608 495023 94990 495051
rect 90548 493400 90600 493406
rect 90548 493342 90600 493348
rect 90652 489914 90680 495023
rect 91112 492590 91140 495023
rect 91100 492584 91152 492590
rect 91480 492538 91508 495023
rect 91100 492526 91152 492532
rect 89916 489886 90680 489914
rect 91204 492510 91508 492538
rect 89812 463344 89864 463350
rect 89812 463286 89864 463292
rect 88524 463276 88576 463282
rect 88524 463218 88576 463224
rect 88432 463208 88484 463214
rect 88432 463150 88484 463156
rect 87144 463140 87196 463146
rect 87144 463082 87196 463088
rect 87052 462936 87104 462942
rect 87052 462878 87104 462884
rect 86224 462324 86276 462330
rect 86224 462266 86276 462272
rect 80058 459096 80114 459105
rect 80058 459031 80114 459040
rect 89916 458969 89944 489886
rect 91204 463690 91232 492510
rect 92032 489914 92060 495023
rect 92572 492584 92624 492590
rect 92572 492526 92624 492532
rect 92480 492516 92532 492522
rect 92480 492458 92532 492464
rect 91296 489886 92060 489914
rect 91192 463684 91244 463690
rect 91192 463626 91244 463632
rect 89902 458960 89958 458969
rect 89902 458895 89958 458904
rect 60740 458856 60792 458862
rect 91296 458833 91324 489886
rect 92492 459270 92520 492458
rect 92584 460358 92612 492526
rect 92676 465905 92704 495023
rect 92952 492522 92980 495023
rect 93320 492590 93348 495023
rect 93308 492584 93360 492590
rect 93308 492526 93360 492532
rect 92940 492516 92992 492522
rect 92940 492458 92992 492464
rect 92662 465896 92718 465905
rect 92662 465831 92718 465840
rect 93872 463049 93900 495023
rect 94148 492538 94176 495023
rect 93964 492510 94176 492538
rect 93858 463040 93914 463049
rect 93858 462975 93914 462984
rect 93964 462913 93992 492510
rect 94608 489914 94636 495023
rect 95344 491978 95372 495037
rect 95436 495023 95818 495051
rect 95332 491972 95384 491978
rect 95332 491914 95384 491920
rect 94056 489886 94636 489914
rect 94056 468994 94084 489886
rect 94044 468988 94096 468994
rect 94044 468930 94096 468936
rect 95436 463078 95464 495023
rect 96264 490618 96292 495037
rect 96252 490612 96304 490618
rect 96252 490554 96304 490560
rect 96724 489054 96752 495037
rect 96816 495023 97198 495051
rect 96712 489048 96764 489054
rect 96712 488990 96764 488996
rect 96816 488986 96844 495023
rect 97552 492114 97580 495037
rect 97540 492108 97592 492114
rect 97540 492050 97592 492056
rect 98012 489122 98040 495037
rect 98104 495023 98486 495051
rect 98656 495023 98946 495051
rect 98104 489870 98132 495023
rect 98656 489914 98684 495023
rect 99392 493338 99420 495037
rect 99484 495023 99774 495051
rect 99380 493332 99432 493338
rect 99380 493274 99432 493280
rect 98196 489886 98684 489914
rect 98092 489864 98144 489870
rect 98092 489806 98144 489812
rect 98000 489116 98052 489122
rect 98000 489058 98052 489064
rect 96804 488980 96856 488986
rect 96804 488922 96856 488928
rect 98196 465798 98224 489886
rect 98184 465792 98236 465798
rect 98184 465734 98236 465740
rect 99484 465730 99512 495023
rect 100220 492182 100248 495037
rect 100312 495023 100694 495051
rect 100772 495023 101154 495051
rect 101232 495023 101522 495051
rect 101600 495023 101982 495051
rect 100208 492176 100260 492182
rect 100208 492118 100260 492124
rect 100312 489914 100340 495023
rect 99576 489886 100340 489914
rect 99472 465724 99524 465730
rect 99472 465666 99524 465672
rect 95424 463072 95476 463078
rect 95424 463014 95476 463020
rect 93950 462904 94006 462913
rect 93950 462839 94006 462848
rect 92572 460352 92624 460358
rect 92572 460294 92624 460300
rect 92480 459264 92532 459270
rect 92480 459206 92532 459212
rect 99576 459202 99604 489886
rect 100772 463010 100800 495023
rect 101232 492538 101260 495023
rect 100864 492510 101260 492538
rect 100864 465934 100892 492510
rect 101600 489914 101628 495023
rect 102232 492516 102284 492522
rect 102232 492458 102284 492464
rect 100956 489886 101628 489914
rect 100956 466002 100984 489886
rect 102244 468790 102272 492458
rect 102428 492250 102456 495037
rect 102520 495023 102902 495051
rect 103072 495023 103362 495051
rect 103624 495023 103730 495051
rect 103808 495023 104190 495051
rect 102416 492244 102468 492250
rect 102416 492186 102468 492192
rect 102520 489914 102548 495023
rect 103072 492522 103100 495023
rect 103060 492516 103112 492522
rect 103060 492458 103112 492464
rect 102336 489886 102548 489914
rect 102232 468784 102284 468790
rect 102232 468726 102284 468732
rect 102336 466070 102364 489886
rect 103624 468858 103652 495023
rect 103808 489914 103836 495023
rect 104636 492386 104664 495037
rect 104912 495023 105110 495051
rect 105188 495023 105570 495051
rect 105648 495023 105938 495051
rect 106292 495023 106398 495051
rect 106476 495023 106858 495051
rect 106936 495023 107318 495051
rect 104624 492380 104676 492386
rect 104624 492322 104676 492328
rect 104912 492318 104940 495023
rect 105188 492504 105216 495023
rect 105004 492476 105216 492504
rect 104900 492312 104952 492318
rect 104900 492254 104952 492260
rect 103716 489886 103836 489914
rect 103612 468852 103664 468858
rect 103612 468794 103664 468800
rect 102324 466064 102376 466070
rect 102324 466006 102376 466012
rect 100944 465996 100996 466002
rect 100944 465938 100996 465944
rect 100852 465928 100904 465934
rect 100852 465870 100904 465876
rect 100760 463004 100812 463010
rect 100760 462946 100812 462952
rect 103716 460290 103744 489886
rect 105004 468926 105032 492476
rect 105648 489914 105676 495023
rect 106292 492454 106320 495023
rect 106372 492516 106424 492522
rect 106372 492458 106424 492464
rect 106280 492448 106332 492454
rect 106280 492390 106332 492396
rect 105096 489886 105676 489914
rect 104992 468920 105044 468926
rect 104992 468862 105044 468868
rect 105096 468586 105124 489886
rect 106384 468722 106412 492458
rect 106372 468716 106424 468722
rect 106372 468658 106424 468664
rect 106476 468654 106504 495023
rect 106936 492522 106964 495023
rect 106924 492516 106976 492522
rect 106924 492458 106976 492464
rect 107660 492516 107712 492522
rect 107660 492458 107712 492464
rect 106464 468648 106516 468654
rect 106464 468590 106516 468596
rect 105084 468580 105136 468586
rect 105084 468522 105136 468528
rect 107672 462913 107700 492458
rect 107764 463010 107792 495037
rect 107856 495023 108146 495051
rect 108224 495023 108606 495051
rect 107856 492522 107884 495023
rect 107844 492516 107896 492522
rect 107844 492458 107896 492464
rect 108224 489914 108252 495023
rect 107856 489886 108252 489914
rect 107856 465798 107884 489886
rect 107844 465792 107896 465798
rect 107844 465734 107896 465740
rect 109052 465730 109080 495037
rect 109542 495023 109816 495051
rect 109910 495023 110184 495051
rect 109788 493338 109816 495023
rect 109776 493332 109828 493338
rect 109776 493274 109828 493280
rect 110156 492114 110184 495023
rect 110144 492108 110196 492114
rect 110144 492050 110196 492056
rect 110340 491978 110368 495037
rect 110328 491972 110380 491978
rect 110328 491914 110380 491920
rect 110800 489530 110828 495037
rect 111260 489734 111288 495037
rect 111248 489728 111300 489734
rect 111248 489670 111300 489676
rect 111720 489598 111748 495037
rect 111892 490408 111944 490414
rect 111892 490350 111944 490356
rect 111708 489592 111760 489598
rect 111708 489534 111760 489540
rect 110788 489524 110840 489530
rect 110788 489466 110840 489472
rect 111904 467158 111932 490350
rect 112088 489666 112116 495037
rect 112272 495023 112562 495051
rect 112640 495023 113022 495051
rect 113376 495023 113482 495051
rect 112076 489660 112128 489666
rect 112076 489602 112128 489608
rect 112272 485774 112300 495023
rect 112640 490414 112668 495023
rect 112628 490408 112680 490414
rect 112628 490350 112680 490356
rect 111996 485746 112300 485774
rect 111892 467152 111944 467158
rect 111892 467094 111944 467100
rect 109040 465724 109092 465730
rect 109040 465666 109092 465672
rect 107752 463004 107804 463010
rect 107752 462946 107804 462952
rect 107658 462904 107714 462913
rect 107658 462839 107714 462848
rect 111996 461786 112024 485746
rect 113376 465866 113404 495023
rect 113928 486266 113956 495037
rect 114296 487830 114324 495037
rect 114572 495023 114770 495051
rect 114284 487824 114336 487830
rect 114284 487766 114336 487772
rect 113916 486260 113968 486266
rect 113916 486202 113968 486208
rect 114572 482322 114600 495023
rect 115216 489394 115244 495037
rect 115676 489569 115704 495037
rect 115662 489560 115718 489569
rect 115662 489495 115718 489504
rect 116044 489462 116072 495037
rect 116032 489456 116084 489462
rect 116032 489398 116084 489404
rect 115204 489388 115256 489394
rect 115204 489330 115256 489336
rect 116504 487082 116532 495037
rect 116964 487150 116992 495037
rect 116952 487144 117004 487150
rect 116952 487086 117004 487092
rect 116492 487076 116544 487082
rect 116492 487018 116544 487024
rect 117424 486878 117452 495037
rect 117412 486872 117464 486878
rect 117412 486814 117464 486820
rect 117884 486810 117912 495037
rect 117872 486804 117924 486810
rect 117872 486746 117924 486752
rect 118252 486742 118280 495037
rect 118742 495023 118832 495051
rect 118700 492516 118752 492522
rect 118700 492458 118752 492464
rect 118712 489802 118740 492458
rect 118700 489796 118752 489802
rect 118700 489738 118752 489744
rect 118240 486736 118292 486742
rect 118240 486678 118292 486684
rect 118804 486402 118832 495023
rect 118896 495023 119186 495051
rect 119264 495023 119646 495051
rect 120122 495023 120212 495051
rect 118792 486396 118844 486402
rect 118792 486338 118844 486344
rect 118896 486334 118924 495023
rect 119264 492522 119292 495023
rect 119252 492516 119304 492522
rect 119252 492458 119304 492464
rect 120080 492516 120132 492522
rect 120080 492458 120132 492464
rect 118884 486328 118936 486334
rect 118884 486270 118936 486276
rect 114560 482316 114612 482322
rect 114560 482258 114612 482264
rect 113364 465860 113416 465866
rect 113364 465802 113416 465808
rect 111984 461780 112036 461786
rect 111984 461722 112036 461728
rect 103704 460284 103756 460290
rect 103704 460226 103756 460232
rect 99564 459196 99616 459202
rect 99564 459138 99616 459144
rect 120092 459134 120120 492458
rect 120184 489297 120212 495023
rect 120276 495023 120474 495051
rect 120552 495023 120934 495051
rect 121104 495023 121394 495051
rect 121564 495023 121854 495051
rect 121932 495023 122222 495051
rect 122300 495023 122682 495051
rect 123036 495023 123142 495051
rect 123312 495023 123602 495051
rect 123680 495023 124062 495051
rect 124232 495023 124430 495051
rect 124600 495023 124890 495051
rect 124968 495023 125350 495051
rect 120276 489433 120304 495023
rect 120552 492522 120580 495023
rect 120540 492516 120592 492522
rect 120540 492458 120592 492464
rect 121104 489914 121132 495023
rect 121460 492244 121512 492250
rect 121460 492186 121512 492192
rect 120368 489886 121132 489914
rect 120368 489705 120396 489886
rect 120354 489696 120410 489705
rect 120354 489631 120410 489640
rect 120262 489424 120318 489433
rect 120262 489359 120318 489368
rect 120170 489288 120226 489297
rect 120170 489223 120226 489232
rect 121472 486985 121500 492186
rect 121564 487014 121592 495023
rect 121932 492250 121960 495023
rect 121920 492244 121972 492250
rect 121920 492186 121972 492192
rect 122300 489914 122328 495023
rect 122932 492516 122984 492522
rect 122932 492458 122984 492464
rect 122840 492448 122892 492454
rect 122840 492390 122892 492396
rect 121656 489886 122328 489914
rect 121552 487008 121604 487014
rect 121458 486976 121514 486985
rect 121552 486950 121604 486956
rect 121458 486911 121514 486920
rect 121656 486849 121684 489886
rect 121642 486840 121698 486849
rect 121642 486775 121698 486784
rect 122852 483993 122880 492390
rect 122944 484022 122972 492458
rect 123036 486713 123064 495023
rect 123312 492522 123340 495023
rect 123300 492516 123352 492522
rect 123300 492458 123352 492464
rect 123680 492454 123708 495023
rect 123668 492448 123720 492454
rect 123668 492390 123720 492396
rect 123022 486704 123078 486713
rect 123022 486639 123078 486648
rect 124232 484226 124260 495023
rect 124312 492516 124364 492522
rect 124312 492458 124364 492464
rect 124220 484220 124272 484226
rect 124220 484162 124272 484168
rect 124324 484090 124352 492458
rect 124600 489914 124628 495023
rect 124968 492522 124996 495023
rect 124956 492516 125008 492522
rect 124956 492458 125008 492464
rect 125692 492516 125744 492522
rect 125692 492458 125744 492464
rect 125600 492448 125652 492454
rect 125600 492390 125652 492396
rect 124416 489886 124628 489914
rect 124312 484084 124364 484090
rect 124312 484026 124364 484032
rect 122932 484016 122984 484022
rect 122838 483984 122894 483993
rect 122932 483958 122984 483964
rect 124416 483954 124444 489886
rect 122838 483919 122894 483928
rect 124404 483948 124456 483954
rect 124404 483890 124456 483896
rect 125612 460290 125640 492390
rect 125704 483857 125732 492458
rect 125796 489161 125824 495037
rect 125888 495023 126270 495051
rect 126348 495023 126638 495051
rect 125888 492522 125916 495023
rect 125876 492516 125928 492522
rect 125876 492458 125928 492464
rect 126348 492454 126376 495023
rect 126980 492516 127032 492522
rect 126980 492458 127032 492464
rect 126336 492448 126388 492454
rect 126336 492390 126388 492396
rect 125782 489152 125838 489161
rect 125782 489087 125838 489096
rect 125690 483848 125746 483857
rect 125690 483783 125746 483792
rect 126992 483721 127020 492458
rect 127084 486577 127112 495037
rect 127176 495023 127558 495051
rect 127728 495023 128018 495051
rect 127176 492522 127204 495023
rect 127164 492516 127216 492522
rect 127164 492458 127216 492464
rect 127728 489914 127756 495023
rect 128360 494964 128412 494970
rect 128360 494906 128412 494912
rect 127176 489886 127756 489914
rect 127070 486568 127126 486577
rect 127070 486503 127126 486512
rect 127176 486441 127204 489886
rect 127162 486432 127218 486441
rect 127162 486367 127218 486376
rect 126978 483712 127034 483721
rect 126978 483647 127034 483656
rect 128372 483614 128400 494906
rect 128464 492674 128492 495037
rect 128556 495023 128846 495051
rect 129016 495023 129306 495051
rect 129782 495023 129964 495051
rect 128556 494970 128584 495023
rect 128544 494964 128596 494970
rect 128544 494906 128596 494912
rect 128464 492646 128584 492674
rect 128556 492402 128584 492646
rect 128464 492374 128584 492402
rect 128464 484362 128492 492374
rect 129016 489914 129044 495023
rect 129936 492590 129964 495023
rect 130028 495023 130226 495051
rect 130304 495023 130594 495051
rect 130672 495023 131054 495051
rect 131316 495023 131514 495051
rect 131592 495023 131974 495051
rect 132144 495023 132434 495051
rect 132512 495023 132802 495051
rect 132880 495023 133262 495051
rect 133432 495023 133722 495051
rect 133892 495023 134182 495051
rect 134352 495023 134642 495051
rect 134720 495023 135010 495051
rect 135272 495023 135470 495051
rect 135640 495023 135930 495051
rect 136008 495023 136390 495051
rect 129924 492584 129976 492590
rect 129924 492526 129976 492532
rect 129740 492516 129792 492522
rect 129740 492458 129792 492464
rect 129648 492040 129700 492046
rect 129648 491982 129700 491988
rect 128556 489886 129044 489914
rect 128556 486538 128584 489886
rect 129660 487801 129688 491982
rect 129752 489258 129780 492458
rect 130028 492402 130056 495023
rect 130108 492584 130160 492590
rect 130108 492526 130160 492532
rect 129844 492374 130056 492402
rect 129740 489252 129792 489258
rect 129740 489194 129792 489200
rect 129646 487792 129702 487801
rect 129646 487727 129702 487736
rect 128544 486532 128596 486538
rect 128544 486474 128596 486480
rect 129844 486470 129872 492374
rect 130120 492266 130148 492526
rect 129936 492238 130148 492266
rect 129936 486674 129964 492238
rect 130304 489914 130332 495023
rect 130672 492522 130700 495023
rect 130660 492516 130712 492522
rect 130660 492458 130712 492464
rect 131120 492516 131172 492522
rect 131120 492458 131172 492464
rect 130028 489886 130332 489914
rect 130028 486946 130056 489886
rect 130016 486940 130068 486946
rect 130016 486882 130068 486888
rect 129924 486668 129976 486674
rect 129924 486610 129976 486616
rect 129832 486464 129884 486470
rect 129832 486406 129884 486412
rect 128452 484356 128504 484362
rect 128452 484298 128504 484304
rect 128360 483608 128412 483614
rect 128360 483550 128412 483556
rect 125600 460284 125652 460290
rect 125600 460226 125652 460232
rect 120080 459128 120132 459134
rect 120080 459070 120132 459076
rect 131132 459066 131160 492458
rect 131212 492448 131264 492454
rect 131212 492390 131264 492396
rect 131224 483750 131252 492390
rect 131316 486606 131344 495023
rect 131592 492522 131620 495023
rect 131580 492516 131632 492522
rect 131580 492458 131632 492464
rect 132144 492454 132172 495023
rect 132132 492448 132184 492454
rect 132132 492390 132184 492396
rect 132512 489326 132540 495023
rect 132880 492538 132908 495023
rect 132604 492510 132908 492538
rect 132500 489320 132552 489326
rect 132500 489262 132552 489268
rect 131304 486600 131356 486606
rect 131304 486542 131356 486548
rect 132604 483818 132632 492510
rect 133432 489914 133460 495023
rect 132696 489886 133460 489914
rect 132696 483886 132724 489886
rect 132684 483880 132736 483886
rect 132684 483822 132736 483828
rect 132592 483812 132644 483818
rect 132592 483754 132644 483760
rect 131212 483744 131264 483750
rect 131212 483686 131264 483692
rect 131120 459060 131172 459066
rect 131120 459002 131172 459008
rect 133892 458930 133920 495023
rect 133972 492516 134024 492522
rect 133972 492458 134024 492464
rect 133984 458998 134012 492458
rect 134352 489914 134380 495023
rect 134720 492522 134748 495023
rect 134708 492516 134760 492522
rect 134708 492458 134760 492464
rect 134076 489886 134380 489914
rect 134076 484294 134104 489886
rect 134064 484288 134116 484294
rect 134064 484230 134116 484236
rect 135272 458998 135300 495023
rect 135352 492516 135404 492522
rect 135352 492458 135404 492464
rect 135364 484158 135392 492458
rect 135640 489914 135668 495023
rect 136008 492522 136036 495023
rect 136640 494964 136692 494970
rect 136640 494906 136692 494912
rect 135996 492516 136048 492522
rect 135996 492458 136048 492464
rect 135456 489886 135668 489914
rect 135456 489326 135484 489886
rect 135444 489320 135496 489326
rect 135444 489262 135496 489268
rect 135352 484152 135404 484158
rect 135352 484094 135404 484100
rect 136652 459066 136680 494906
rect 136744 492674 136772 495037
rect 136928 495023 137218 495051
rect 137296 495023 137678 495051
rect 136928 494970 136956 495023
rect 136916 494964 136968 494970
rect 136916 494906 136968 494912
rect 136744 492646 136864 492674
rect 136836 492402 136864 492646
rect 136744 492374 136864 492402
rect 136744 489462 136772 492374
rect 137296 489914 137324 495023
rect 138020 492516 138072 492522
rect 138020 492458 138072 492464
rect 136836 489886 137324 489914
rect 136732 489456 136784 489462
rect 136732 489398 136784 489404
rect 136836 489258 136864 489886
rect 136824 489252 136876 489258
rect 136824 489194 136876 489200
rect 136640 459060 136692 459066
rect 136640 459002 136692 459008
rect 133972 458992 134024 458998
rect 133972 458934 134024 458940
rect 135260 458992 135312 458998
rect 135260 458934 135312 458940
rect 138032 458930 138060 492458
rect 138124 489394 138152 495037
rect 138216 495023 138598 495051
rect 138676 495023 138966 495051
rect 138216 489530 138244 495023
rect 138676 492522 138704 495023
rect 139412 492658 139440 495037
rect 139504 495023 139886 495051
rect 140056 495023 140346 495051
rect 139400 492652 139452 492658
rect 139400 492594 139452 492600
rect 138664 492516 138716 492522
rect 138664 492458 138716 492464
rect 139400 492516 139452 492522
rect 139400 492458 139452 492464
rect 138204 489524 138256 489530
rect 138204 489466 138256 489472
rect 138112 489388 138164 489394
rect 138112 489330 138164 489336
rect 139412 466138 139440 492458
rect 139400 466132 139452 466138
rect 139400 466074 139452 466080
rect 139504 465866 139532 495023
rect 139860 492652 139912 492658
rect 139860 492594 139912 492600
rect 139872 492046 139900 492594
rect 140056 492522 140084 495023
rect 140044 492516 140096 492522
rect 140044 492458 140096 492464
rect 139860 492040 139912 492046
rect 139860 491982 139912 491988
rect 140792 466206 140820 495037
rect 140884 495023 141174 495051
rect 141344 495023 141634 495051
rect 141712 495023 142094 495051
rect 142264 495023 142554 495051
rect 142632 495023 142922 495051
rect 143000 495023 143382 495051
rect 143644 495023 143842 495051
rect 143920 495023 144302 495051
rect 144472 495023 144762 495051
rect 140780 466200 140832 466206
rect 140780 466142 140832 466148
rect 140884 466070 140912 495023
rect 140964 492516 141016 492522
rect 140964 492458 141016 492464
rect 140872 466064 140924 466070
rect 140872 466006 140924 466012
rect 140976 466002 141004 492458
rect 141344 489914 141372 495023
rect 141712 492522 141740 495023
rect 141700 492516 141752 492522
rect 141700 492458 141752 492464
rect 142160 491292 142212 491298
rect 142160 491234 142212 491240
rect 141068 489886 141372 489914
rect 140964 465996 141016 466002
rect 140964 465938 141016 465944
rect 141068 465934 141096 489886
rect 141056 465928 141108 465934
rect 141056 465870 141108 465876
rect 139492 465860 139544 465866
rect 139492 465802 139544 465808
rect 142172 459134 142200 491234
rect 142264 463078 142292 495023
rect 142632 491298 142660 495023
rect 142620 491292 142672 491298
rect 142620 491234 142672 491240
rect 143000 489914 143028 495023
rect 143540 492516 143592 492522
rect 143540 492458 143592 492464
rect 142356 489886 143028 489914
rect 142356 463146 142384 489886
rect 143552 478145 143580 492458
rect 143644 483682 143672 495023
rect 143920 492522 143948 495023
rect 143908 492516 143960 492522
rect 143908 492458 143960 492464
rect 144472 489914 144500 495023
rect 145116 491881 145144 495037
rect 145208 495023 145590 495051
rect 145760 495023 146050 495051
rect 146526 495023 146616 495051
rect 145102 491872 145158 491881
rect 145102 491807 145158 491816
rect 145208 491722 145236 495023
rect 143736 489886 144500 489914
rect 144932 491694 145236 491722
rect 143736 486441 143764 489886
rect 143722 486432 143778 486441
rect 143722 486367 143778 486376
rect 143632 483676 143684 483682
rect 143632 483618 143684 483624
rect 143538 478136 143594 478145
rect 143538 478071 143594 478080
rect 144932 472569 144960 491694
rect 145760 489914 145788 495023
rect 146300 492516 146352 492522
rect 146300 492458 146352 492464
rect 145024 489886 145788 489914
rect 145024 483721 145052 489886
rect 145010 483712 145066 483721
rect 145010 483647 145066 483656
rect 146312 475425 146340 492458
rect 146588 492017 146616 495023
rect 146680 495023 146970 495051
rect 147048 495023 147338 495051
rect 146574 492008 146630 492017
rect 146574 491943 146630 491952
rect 146680 489914 146708 495023
rect 147048 492522 147076 495023
rect 147036 492516 147088 492522
rect 147036 492458 147088 492464
rect 147784 492289 147812 495037
rect 147876 495023 148258 495051
rect 148336 495023 148718 495051
rect 147770 492280 147826 492289
rect 147770 492215 147826 492224
rect 147876 492130 147904 495023
rect 146404 489886 146708 489914
rect 147692 492102 147904 492130
rect 146404 478174 146432 489886
rect 146392 478168 146444 478174
rect 146392 478110 146444 478116
rect 146298 475416 146354 475425
rect 146298 475351 146354 475360
rect 144918 472560 144974 472569
rect 144918 472495 144974 472504
rect 147692 465769 147720 492102
rect 148336 489914 148364 495023
rect 149164 492153 149192 495037
rect 149256 495023 149546 495051
rect 150022 495023 150296 495051
rect 149150 492144 149206 492153
rect 149150 492079 149206 492088
rect 149256 489914 149284 495023
rect 150268 492425 150296 495023
rect 150452 492658 150480 495037
rect 150544 495023 150926 495051
rect 151310 495023 151492 495051
rect 150440 492652 150492 492658
rect 150440 492594 150492 492600
rect 150440 492516 150492 492522
rect 150440 492458 150492 492464
rect 150254 492416 150310 492425
rect 150254 492351 150310 492360
rect 147784 489886 148364 489914
rect 149072 489886 149284 489914
rect 147784 486577 147812 489886
rect 147770 486568 147826 486577
rect 147770 486503 147826 486512
rect 149072 481030 149100 489886
rect 149060 481024 149112 481030
rect 149060 480966 149112 480972
rect 147678 465760 147734 465769
rect 147678 465695 147734 465704
rect 142344 463140 142396 463146
rect 142344 463082 142396 463088
rect 142252 463072 142304 463078
rect 142252 463014 142304 463020
rect 142160 459128 142212 459134
rect 142160 459070 142212 459076
rect 133880 458924 133932 458930
rect 133880 458866 133932 458872
rect 138020 458924 138072 458930
rect 138020 458866 138072 458872
rect 150452 458833 150480 492458
rect 150544 479505 150572 495023
rect 151464 492318 151492 495023
rect 151556 495023 151754 495051
rect 152230 495023 152320 495051
rect 151556 492522 151584 495023
rect 151544 492516 151596 492522
rect 151544 492458 151596 492464
rect 151452 492312 151504 492318
rect 151452 492254 151504 492260
rect 152292 492182 152320 495023
rect 152384 495023 152674 495051
rect 152280 492176 152332 492182
rect 152280 492118 152332 492124
rect 152384 489914 152412 495023
rect 153120 492454 153148 495037
rect 153518 495023 153792 495051
rect 153108 492448 153160 492454
rect 153108 492390 153160 492396
rect 153764 490521 153792 495023
rect 153948 491842 153976 495037
rect 154040 495023 154422 495051
rect 154898 495023 155264 495051
rect 153936 491836 153988 491842
rect 153936 491778 153988 491784
rect 153750 490512 153806 490521
rect 153750 490447 153806 490456
rect 154040 489914 154068 495023
rect 155236 492250 155264 495023
rect 155328 492590 155356 495037
rect 155420 495023 155710 495051
rect 155972 495023 156170 495051
rect 156646 495023 156736 495051
rect 155316 492584 155368 492590
rect 155316 492526 155368 492532
rect 155224 492244 155276 492250
rect 155224 492186 155276 492192
rect 155420 489914 155448 495023
rect 151832 489886 152412 489914
rect 153212 489886 154068 489914
rect 154592 489886 155448 489914
rect 150530 479496 150586 479505
rect 150530 479431 150586 479440
rect 151832 476785 151860 489886
rect 151818 476776 151874 476785
rect 151818 476711 151874 476720
rect 153212 475561 153240 489886
rect 153198 475552 153254 475561
rect 153198 475487 153254 475496
rect 154592 460329 154620 489886
rect 155972 468489 156000 495023
rect 156708 492658 156736 495023
rect 156800 495023 157090 495051
rect 156696 492652 156748 492658
rect 156696 492594 156748 492600
rect 156800 489914 156828 495023
rect 157340 492516 157392 492522
rect 157340 492458 157392 492464
rect 156064 489886 156828 489914
rect 156064 469849 156092 489886
rect 156050 469840 156106 469849
rect 156050 469775 156106 469784
rect 155958 468480 156014 468489
rect 155958 468415 156014 468424
rect 154578 460320 154634 460329
rect 154578 460255 154634 460264
rect 157352 460193 157380 492458
rect 157444 474065 157472 495037
rect 157934 495023 158024 495051
rect 157996 491910 158024 495023
rect 158088 495023 158378 495051
rect 158732 495023 158838 495051
rect 158916 495023 159298 495051
rect 159376 495023 159666 495051
rect 160142 495023 160232 495051
rect 158088 492522 158116 495023
rect 158076 492516 158128 492522
rect 158076 492458 158128 492464
rect 157984 491904 158036 491910
rect 157984 491846 158036 491852
rect 157430 474056 157486 474065
rect 157430 473991 157486 474000
rect 158732 463185 158760 495023
rect 158916 492538 158944 495023
rect 158824 492510 158944 492538
rect 158824 476814 158852 492510
rect 159376 489914 159404 495023
rect 160100 492516 160152 492522
rect 160100 492458 160152 492464
rect 158916 489886 159404 489914
rect 158916 487830 158944 489886
rect 158904 487824 158956 487830
rect 158904 487766 158956 487772
rect 158812 476808 158864 476814
rect 158812 476750 158864 476756
rect 160112 463282 160140 492458
rect 160204 464370 160232 495023
rect 160296 495023 160586 495051
rect 160664 495023 161046 495051
rect 161522 495023 161704 495051
rect 160296 465905 160324 495023
rect 160664 492522 160692 495023
rect 161572 492788 161624 492794
rect 161572 492730 161624 492736
rect 161480 492720 161532 492726
rect 161480 492662 161532 492668
rect 160652 492516 160704 492522
rect 160652 492458 160704 492464
rect 160836 492448 160888 492454
rect 160836 492390 160888 492396
rect 160848 492182 160876 492390
rect 160836 492176 160888 492182
rect 160836 492118 160888 492124
rect 160928 492176 160980 492182
rect 160928 492118 160980 492124
rect 160940 491842 160968 492118
rect 160928 491836 160980 491842
rect 160928 491778 160980 491784
rect 160282 465896 160338 465905
rect 160282 465831 160338 465840
rect 160192 464364 160244 464370
rect 160192 464306 160244 464312
rect 160100 463276 160152 463282
rect 160100 463218 160152 463224
rect 158718 463176 158774 463185
rect 158718 463111 158774 463120
rect 157338 460184 157394 460193
rect 157338 460119 157394 460128
rect 161492 459105 161520 492662
rect 161584 461553 161612 492730
rect 161676 474026 161704 495023
rect 161768 495023 161874 495051
rect 161952 495023 162334 495051
rect 162412 495023 162794 495051
rect 162964 495023 163254 495051
rect 163332 495023 163622 495051
rect 164098 495023 164188 495051
rect 161768 492726 161796 495023
rect 161952 492794 161980 495023
rect 161940 492788 161992 492794
rect 161940 492730 161992 492736
rect 161756 492720 161808 492726
rect 161756 492662 161808 492668
rect 162412 492538 162440 495023
rect 162860 492720 162912 492726
rect 162860 492662 162912 492668
rect 161768 492510 162440 492538
rect 161768 479534 161796 492510
rect 162124 492108 162176 492114
rect 162124 492050 162176 492056
rect 161756 479528 161808 479534
rect 161756 479470 161808 479476
rect 161664 474020 161716 474026
rect 161664 473962 161716 473968
rect 161570 461544 161626 461553
rect 161570 461479 161626 461488
rect 162136 460494 162164 492050
rect 162124 460488 162176 460494
rect 162124 460430 162176 460436
rect 161478 459096 161534 459105
rect 161478 459031 161534 459040
rect 162872 458969 162900 492662
rect 162964 467158 162992 495023
rect 163332 492726 163360 495023
rect 163320 492720 163372 492726
rect 163320 492662 163372 492668
rect 164160 492114 164188 495023
rect 164344 495023 164542 495051
rect 164712 495023 165002 495051
rect 165080 495023 165462 495051
rect 165632 495023 165830 495051
rect 166000 495023 166290 495051
rect 166766 495023 166948 495051
rect 164240 492720 164292 492726
rect 164240 492662 164292 492668
rect 164148 492108 164200 492114
rect 164148 492050 164200 492056
rect 162952 467152 163004 467158
rect 162952 467094 163004 467100
rect 164252 464438 164280 492662
rect 164344 469985 164372 495023
rect 164712 489914 164740 495023
rect 165080 492726 165108 495023
rect 165068 492720 165120 492726
rect 165068 492662 165120 492668
rect 164436 489886 164740 489914
rect 164436 471306 164464 489886
rect 164424 471300 164476 471306
rect 164424 471242 164476 471248
rect 164330 469976 164386 469985
rect 164330 469911 164386 469920
rect 164240 464432 164292 464438
rect 164240 464374 164292 464380
rect 165632 461786 165660 495023
rect 166000 489914 166028 495023
rect 166920 491774 166948 495023
rect 167000 492788 167052 492794
rect 167000 492730 167052 492736
rect 166908 491768 166960 491774
rect 166908 491710 166960 491716
rect 165724 489886 166028 489914
rect 165724 485110 165752 489886
rect 165712 485104 165764 485110
rect 165712 485046 165764 485052
rect 165620 461780 165672 461786
rect 165620 461722 165672 461728
rect 167012 460465 167040 492730
rect 167092 492720 167144 492726
rect 167092 492662 167144 492668
rect 166998 460456 167054 460465
rect 167104 460426 167132 492662
rect 167196 483682 167224 495037
rect 167288 495023 167670 495051
rect 167748 495023 168038 495051
rect 168392 495023 168498 495051
rect 168576 495023 168958 495051
rect 169128 495023 169418 495051
rect 169894 495023 169984 495051
rect 167288 492726 167316 495023
rect 167748 492794 167776 495023
rect 167736 492788 167788 492794
rect 167736 492730 167788 492736
rect 167276 492720 167328 492726
rect 167276 492662 167328 492668
rect 167184 483676 167236 483682
rect 167184 483618 167236 483624
rect 166998 460391 167054 460400
rect 167092 460420 167144 460426
rect 167092 460362 167144 460368
rect 168392 460358 168420 495023
rect 168472 492720 168524 492726
rect 168472 492662 168524 492668
rect 168484 463214 168512 492662
rect 168576 482322 168604 495023
rect 169128 492726 169156 495023
rect 169116 492720 169168 492726
rect 169116 492662 169168 492668
rect 169852 492720 169904 492726
rect 169852 492662 169904 492668
rect 169760 491836 169812 491842
rect 169760 491778 169812 491784
rect 168564 482316 168616 482322
rect 168564 482258 168616 482264
rect 169772 463321 169800 491778
rect 169864 466041 169892 492662
rect 169850 466032 169906 466041
rect 169850 465967 169906 465976
rect 169758 463312 169814 463321
rect 169758 463247 169814 463256
rect 168472 463208 168524 463214
rect 168472 463150 168524 463156
rect 169956 463049 169984 495023
rect 170048 495023 170246 495051
rect 170416 495023 170706 495051
rect 170048 491842 170076 495023
rect 170416 492726 170444 495023
rect 170404 492720 170456 492726
rect 170404 492662 170456 492668
rect 170036 491836 170088 491842
rect 170036 491778 170088 491784
rect 169942 463040 169998 463049
rect 169942 462975 169998 462984
rect 168380 460352 168432 460358
rect 168380 460294 168432 460300
rect 171152 459241 171180 495037
rect 171336 495023 171626 495051
rect 171704 495023 171994 495051
rect 172072 495023 172454 495051
rect 172532 495023 172914 495051
rect 172992 495023 173374 495051
rect 173544 495023 173834 495051
rect 173912 495023 174202 495051
rect 174280 495023 174662 495051
rect 174832 495023 175122 495051
rect 175384 495023 175582 495051
rect 175752 495023 176042 495051
rect 176120 495023 176410 495051
rect 171232 492720 171284 492726
rect 171232 492662 171284 492668
rect 171244 461854 171272 492662
rect 171232 461848 171284 461854
rect 171232 461790 171284 461796
rect 171336 461689 171364 495023
rect 171704 489914 171732 495023
rect 172072 492726 172100 495023
rect 172060 492720 172112 492726
rect 172060 492662 172112 492668
rect 171428 489886 171732 489914
rect 171428 489161 171456 489886
rect 171414 489152 171470 489161
rect 171414 489087 171470 489096
rect 171322 461680 171378 461689
rect 171322 461615 171378 461624
rect 172532 459377 172560 495023
rect 172612 492720 172664 492726
rect 172612 492662 172664 492668
rect 172624 460698 172652 492662
rect 172992 489914 173020 495023
rect 173544 492726 173572 495023
rect 173532 492720 173584 492726
rect 173532 492662 173584 492668
rect 172716 489886 173020 489914
rect 172716 467129 172744 489886
rect 172702 467120 172758 467129
rect 172702 467055 172758 467064
rect 172612 460692 172664 460698
rect 172612 460634 172664 460640
rect 172518 459368 172574 459377
rect 172518 459303 172574 459312
rect 173912 459270 173940 495023
rect 173992 492720 174044 492726
rect 173992 492662 174044 492668
rect 174004 466274 174032 492662
rect 174280 489914 174308 495023
rect 174832 492726 174860 495023
rect 174820 492720 174872 492726
rect 174820 492662 174872 492668
rect 175280 492720 175332 492726
rect 175280 492662 175332 492668
rect 174096 489886 174308 489914
rect 174096 468586 174124 489886
rect 174084 468580 174136 468586
rect 174084 468522 174136 468528
rect 173992 466268 174044 466274
rect 173992 466210 174044 466216
rect 175292 463418 175320 492662
rect 175384 467226 175412 495023
rect 175752 489914 175780 495023
rect 176120 492726 176148 495023
rect 176752 494964 176804 494970
rect 176752 494906 176804 494912
rect 176108 492720 176160 492726
rect 176108 492662 176160 492668
rect 176660 492720 176712 492726
rect 176660 492662 176712 492668
rect 175476 489886 175780 489914
rect 175476 467294 175504 489886
rect 175464 467288 175516 467294
rect 175464 467230 175516 467236
rect 175372 467220 175424 467226
rect 175372 467162 175424 467168
rect 176672 466342 176700 492662
rect 176764 469946 176792 494906
rect 176872 494850 176900 495037
rect 177040 495023 177330 495051
rect 177408 495023 177790 495051
rect 177040 494970 177068 495023
rect 177028 494964 177080 494970
rect 177028 494906 177080 494912
rect 176872 494822 177068 494850
rect 177040 489954 177068 494822
rect 177408 492726 177436 495023
rect 177396 492720 177448 492726
rect 177396 492662 177448 492668
rect 178040 492720 178092 492726
rect 178040 492662 178092 492668
rect 176872 489926 177068 489954
rect 176872 489914 176900 489926
rect 176856 489886 176900 489914
rect 176856 471374 176884 489886
rect 176844 471368 176896 471374
rect 176844 471310 176896 471316
rect 176752 469940 176804 469946
rect 176752 469882 176804 469888
rect 176660 466336 176712 466342
rect 176660 466278 176712 466284
rect 175280 463412 175332 463418
rect 175280 463354 175332 463360
rect 173900 459264 173952 459270
rect 171138 459232 171194 459241
rect 173900 459206 173952 459212
rect 178052 459202 178080 492662
rect 178144 472734 178172 495037
rect 178236 495023 178618 495051
rect 178696 495023 179078 495051
rect 178236 479602 178264 495023
rect 178696 492726 178724 495023
rect 178684 492720 178736 492726
rect 178684 492662 178736 492668
rect 179420 492720 179472 492726
rect 179420 492662 179472 492668
rect 178224 479596 178276 479602
rect 178224 479538 178276 479544
rect 178132 472728 178184 472734
rect 178132 472670 178184 472676
rect 178316 462324 178368 462330
rect 178316 462266 178368 462272
rect 178328 461417 178356 462266
rect 178314 461408 178370 461417
rect 178314 461343 178370 461352
rect 178328 461038 178356 461343
rect 178316 461032 178368 461038
rect 178316 460974 178368 460980
rect 179432 460562 179460 492662
rect 179524 460630 179552 495037
rect 179616 495023 179998 495051
rect 180076 495023 180366 495051
rect 179616 478281 179644 495023
rect 180076 492726 180104 495023
rect 180064 492720 180116 492726
rect 180064 492662 180116 492668
rect 180064 489184 180116 489190
rect 180064 489126 180116 489132
rect 179602 478272 179658 478281
rect 179602 478207 179658 478216
rect 180076 462330 180104 489126
rect 180064 462324 180116 462330
rect 180064 462266 180116 462272
rect 180076 462233 180104 462266
rect 180062 462224 180118 462233
rect 180062 462159 180118 462168
rect 179512 460624 179564 460630
rect 179512 460566 179564 460572
rect 179420 460556 179472 460562
rect 179420 460498 179472 460504
rect 180812 459338 180840 495037
rect 180996 495023 181286 495051
rect 181456 495023 181746 495051
rect 182222 495023 182312 495051
rect 180892 492720 180944 492726
rect 180892 492662 180944 492668
rect 180904 462942 180932 492662
rect 180996 463350 181024 495023
rect 181456 492726 181484 495023
rect 181444 492720 181496 492726
rect 181444 492662 181496 492668
rect 182180 492720 182232 492726
rect 182180 492662 182232 492668
rect 180984 463344 181036 463350
rect 180984 463286 181036 463292
rect 180892 462936 180944 462942
rect 180892 462878 180944 462884
rect 182192 461922 182220 492662
rect 182284 461990 182312 495023
rect 182376 495023 182574 495051
rect 182744 495023 183034 495051
rect 182376 465594 182404 495023
rect 182744 492726 182772 495023
rect 182732 492720 182784 492726
rect 182732 492662 182784 492668
rect 183480 491774 183508 495037
rect 183572 495023 183954 495051
rect 184032 495023 184322 495051
rect 184400 495023 184782 495051
rect 185044 495023 185242 495051
rect 185718 495023 185808 495051
rect 183468 491768 183520 491774
rect 183468 491710 183520 491716
rect 182364 465588 182416 465594
rect 182364 465530 182416 465536
rect 182272 461984 182324 461990
rect 182272 461926 182324 461932
rect 182180 461916 182232 461922
rect 182180 461858 182232 461864
rect 183572 460902 183600 495023
rect 184032 492538 184060 495023
rect 183664 492510 184060 492538
rect 183664 463457 183692 492510
rect 184400 489914 184428 495023
rect 184940 492720 184992 492726
rect 184940 492662 184992 492668
rect 183756 489886 184428 489914
rect 183756 463486 183784 489886
rect 184952 463554 184980 492662
rect 185044 472802 185072 495023
rect 185780 492561 185808 495023
rect 185872 495023 186162 495051
rect 186424 495023 186530 495051
rect 187006 495023 187096 495051
rect 185872 492726 185900 495023
rect 185860 492720 185912 492726
rect 185860 492662 185912 492668
rect 185766 492552 185822 492561
rect 185766 492487 185822 492496
rect 186320 490408 186372 490414
rect 186320 490350 186372 490356
rect 185032 472796 185084 472802
rect 185032 472738 185084 472744
rect 184940 463548 184992 463554
rect 184940 463490 184992 463496
rect 183744 463480 183796 463486
rect 183650 463448 183706 463457
rect 183744 463422 183796 463428
rect 183650 463383 183706 463392
rect 183560 460896 183612 460902
rect 183560 460838 183612 460844
rect 186332 459513 186360 490350
rect 186424 462194 186452 495023
rect 187068 491745 187096 495023
rect 187160 495023 187450 495051
rect 187804 495023 187910 495051
rect 188080 495023 188370 495051
rect 188448 495023 188738 495051
rect 187054 491736 187110 491745
rect 187054 491671 187110 491680
rect 187160 490414 187188 495023
rect 187148 490408 187200 490414
rect 187148 490350 187200 490356
rect 187700 490204 187752 490210
rect 187700 490146 187752 490152
rect 186412 462188 186464 462194
rect 186412 462130 186464 462136
rect 187712 460154 187740 490146
rect 187804 462874 187832 495023
rect 188080 485774 188108 495023
rect 188448 490210 188476 495023
rect 188436 490204 188488 490210
rect 188436 490146 188488 490152
rect 189080 486804 189132 486810
rect 189080 486746 189132 486752
rect 187896 485746 188108 485774
rect 187896 465662 187924 485746
rect 187884 465656 187936 465662
rect 187884 465598 187936 465604
rect 187792 462868 187844 462874
rect 187792 462810 187844 462816
rect 187700 460148 187752 460154
rect 187700 460090 187752 460096
rect 186318 459504 186374 459513
rect 186318 459439 186374 459448
rect 180800 459332 180852 459338
rect 180800 459274 180852 459280
rect 171138 459167 171194 459176
rect 178040 459196 178092 459202
rect 178040 459138 178092 459144
rect 162858 458960 162914 458969
rect 162858 458895 162914 458904
rect 60740 458798 60792 458804
rect 91282 458824 91338 458833
rect 91282 458759 91338 458768
rect 150438 458824 150494 458833
rect 189092 458794 189120 486746
rect 189184 459406 189212 495037
rect 189276 495023 189658 495051
rect 189736 495023 190118 495051
rect 189276 460766 189304 495023
rect 189736 486810 189764 495023
rect 190184 492176 190236 492182
rect 190184 492118 190236 492124
rect 190196 492046 190224 492118
rect 190092 492040 190144 492046
rect 190092 491982 190144 491988
rect 190184 492040 190236 492046
rect 190184 491982 190236 491988
rect 190104 491638 190132 491982
rect 190092 491632 190144 491638
rect 190092 491574 190144 491580
rect 189724 486804 189776 486810
rect 189724 486746 189776 486752
rect 190472 463622 190500 495037
rect 190564 495023 190946 495051
rect 191024 495023 191406 495051
rect 191882 495023 191972 495051
rect 190564 463690 190592 495023
rect 191024 485774 191052 495023
rect 191104 492312 191156 492318
rect 191104 492254 191156 492260
rect 191194 492280 191250 492289
rect 191116 491706 191144 492254
rect 191194 492215 191250 492224
rect 191104 491700 191156 491706
rect 191104 491642 191156 491648
rect 191208 491473 191236 492215
rect 191194 491464 191250 491473
rect 191194 491399 191250 491408
rect 191840 490612 191892 490618
rect 191840 490554 191892 490560
rect 190656 485746 191052 485774
rect 190656 466410 190684 485746
rect 190644 466404 190696 466410
rect 190644 466346 190696 466352
rect 190552 463684 190604 463690
rect 190552 463626 190604 463632
rect 190460 463616 190512 463622
rect 190460 463558 190512 463564
rect 190918 461000 190974 461009
rect 190918 460935 190920 460944
rect 190972 460935 190974 460944
rect 190920 460906 190972 460912
rect 189264 460760 189316 460766
rect 189264 460702 189316 460708
rect 191852 459542 191880 490554
rect 191944 462126 191972 495023
rect 192036 495023 192326 495051
rect 192404 495023 192694 495051
rect 192864 495023 193154 495051
rect 193324 495023 193614 495051
rect 193784 495023 194074 495051
rect 191932 462120 191984 462126
rect 191932 462062 191984 462068
rect 192036 462058 192064 495023
rect 192404 490618 192432 495023
rect 192484 491972 192536 491978
rect 192484 491914 192536 491920
rect 192392 490612 192444 490618
rect 192392 490554 192444 490560
rect 192116 490408 192168 490414
rect 192116 490350 192168 490356
rect 192128 465526 192156 490350
rect 192116 465520 192168 465526
rect 192116 465462 192168 465468
rect 192496 462262 192524 491914
rect 192864 490414 192892 495023
rect 192852 490408 192904 490414
rect 192852 490350 192904 490356
rect 193220 490408 193272 490414
rect 193220 490350 193272 490356
rect 192484 462256 192536 462262
rect 192484 462198 192536 462204
rect 192024 462052 192076 462058
rect 192024 461994 192076 462000
rect 193232 460086 193260 490350
rect 193324 462806 193352 495023
rect 193784 490414 193812 495023
rect 194520 491978 194548 495037
rect 194918 495023 195008 495051
rect 194980 492182 195008 495023
rect 195072 495023 195362 495051
rect 195440 495023 195822 495051
rect 196298 495023 196664 495051
rect 194968 492176 195020 492182
rect 194968 492118 195020 492124
rect 194508 491972 194560 491978
rect 194508 491914 194560 491920
rect 193864 491632 193916 491638
rect 193864 491574 193916 491580
rect 193772 490408 193824 490414
rect 193772 490350 193824 490356
rect 193312 462800 193364 462806
rect 193312 462742 193364 462748
rect 193876 460834 193904 491574
rect 194600 490408 194652 490414
rect 194600 490350 194652 490356
rect 193864 460828 193916 460834
rect 193864 460770 193916 460776
rect 193220 460080 193272 460086
rect 193220 460022 193272 460028
rect 191840 459536 191892 459542
rect 191840 459478 191892 459484
rect 194612 459474 194640 490350
rect 195072 485774 195100 495023
rect 195440 490414 195468 495023
rect 195428 490408 195480 490414
rect 195428 490350 195480 490356
rect 194704 485746 195100 485774
rect 194704 460018 194732 485746
rect 194692 460012 194744 460018
rect 194692 459954 194744 459960
rect 194600 459468 194652 459474
rect 194600 459410 194652 459416
rect 189172 459400 189224 459406
rect 189172 459342 189224 459348
rect 150438 458759 150494 458768
rect 189080 458788 189132 458794
rect 189080 458730 189132 458736
rect 105450 375048 105506 375057
rect 105450 374983 105506 374992
rect 60740 374944 60792 374950
rect 60740 374886 60792 374892
rect 60752 349110 60780 374886
rect 62120 374876 62172 374882
rect 62120 374818 62172 374824
rect 60740 349104 60792 349110
rect 60740 349046 60792 349052
rect 62132 348702 62160 374818
rect 105464 374066 105492 374983
rect 140962 374912 141018 374921
rect 140962 374847 141018 374856
rect 140976 374814 141004 374847
rect 140964 374808 141016 374814
rect 140964 374750 141016 374756
rect 163410 374640 163466 374649
rect 163410 374575 163466 374584
rect 165986 374640 166042 374649
rect 165986 374575 165988 374584
rect 163424 374542 163452 374575
rect 166040 374575 166042 374584
rect 179326 374640 179382 374649
rect 179326 374575 179382 374584
rect 165988 374546 166040 374552
rect 163412 374536 163464 374542
rect 143538 374504 143594 374513
rect 143538 374439 143594 374448
rect 153474 374504 153530 374513
rect 153474 374439 153530 374448
rect 158534 374504 158590 374513
rect 158534 374439 158536 374448
rect 143552 374134 143580 374439
rect 148966 374368 149022 374377
rect 153488 374338 153516 374439
rect 158588 374439 158590 374448
rect 160926 374504 160982 374513
rect 163412 374478 163464 374484
rect 160926 374439 160982 374448
rect 158536 374410 158588 374416
rect 160940 374406 160968 374439
rect 160928 374400 160980 374406
rect 160928 374342 160980 374348
rect 148966 374303 149022 374312
rect 153476 374332 153528 374338
rect 148980 374270 149008 374303
rect 153476 374274 153528 374280
rect 148968 374264 149020 374270
rect 146206 374232 146262 374241
rect 148968 374206 149020 374212
rect 146206 374167 146208 374176
rect 146260 374167 146262 374176
rect 146208 374138 146260 374144
rect 143540 374128 143592 374134
rect 143540 374070 143592 374076
rect 105452 374060 105504 374066
rect 105452 374002 105504 374008
rect 116124 373924 116176 373930
rect 116124 373866 116176 373872
rect 139216 373924 139268 373930
rect 139216 373866 139268 373872
rect 103520 373856 103572 373862
rect 98366 373824 98422 373833
rect 98366 373759 98422 373768
rect 103518 373824 103520 373833
rect 103572 373824 103574 373833
rect 103518 373759 103574 373768
rect 110418 373824 110474 373833
rect 110418 373759 110474 373768
rect 113548 373788 113600 373794
rect 95054 373688 95110 373697
rect 95054 373623 95110 373632
rect 96158 373688 96214 373697
rect 96158 373623 96214 373632
rect 90178 373416 90234 373425
rect 90178 373351 90234 373360
rect 90192 373318 90220 373351
rect 95068 373318 95096 373623
rect 96066 373416 96122 373425
rect 96172 373386 96200 373623
rect 98274 373552 98330 373561
rect 98274 373487 98330 373496
rect 98288 373454 98316 373487
rect 98380 373454 98408 373759
rect 110432 373590 110460 373759
rect 113548 373730 113600 373736
rect 113560 373697 113588 373730
rect 116136 373697 116164 373866
rect 136456 373856 136508 373862
rect 136456 373798 136508 373804
rect 131028 373788 131080 373794
rect 131028 373730 131080 373736
rect 118332 373720 118384 373726
rect 113546 373688 113602 373697
rect 113546 373623 113602 373632
rect 116122 373688 116178 373697
rect 116122 373623 116178 373632
rect 118330 373688 118332 373697
rect 128912 373720 128964 373726
rect 118384 373688 118386 373697
rect 118330 373623 118386 373632
rect 121366 373688 121422 373697
rect 121366 373623 121422 373632
rect 124126 373688 124182 373697
rect 124126 373623 124182 373632
rect 125690 373688 125746 373697
rect 125690 373623 125692 373632
rect 121380 373590 121408 373623
rect 110420 373584 110472 373590
rect 107842 373552 107898 373561
rect 110420 373526 110472 373532
rect 121368 373584 121420 373590
rect 121368 373526 121420 373532
rect 124140 373522 124168 373623
rect 125744 373623 125746 373632
rect 128910 373688 128912 373697
rect 131040 373697 131068 373730
rect 136468 373697 136496 373798
rect 139228 373697 139256 373866
rect 128964 373688 128966 373697
rect 128910 373623 128966 373632
rect 131026 373688 131082 373697
rect 131026 373623 131082 373632
rect 133694 373688 133750 373697
rect 133694 373623 133696 373632
rect 125692 373594 125744 373600
rect 133748 373623 133750 373632
rect 136454 373688 136510 373697
rect 136454 373623 136510 373632
rect 139214 373688 139270 373697
rect 139214 373623 139270 373632
rect 151726 373688 151782 373697
rect 151726 373623 151782 373632
rect 133696 373594 133748 373600
rect 107842 373487 107844 373496
rect 107896 373487 107898 373496
rect 124128 373516 124180 373522
rect 107844 373458 107896 373464
rect 124128 373458 124180 373464
rect 98276 373448 98328 373454
rect 98276 373390 98328 373396
rect 98368 373448 98420 373454
rect 98368 373390 98420 373396
rect 96066 373351 96068 373360
rect 96120 373351 96122 373360
rect 96160 373380 96212 373386
rect 96068 373322 96120 373328
rect 96160 373322 96212 373328
rect 90180 373312 90232 373318
rect 88338 373280 88394 373289
rect 90180 373254 90232 373260
rect 95056 373312 95108 373318
rect 95056 373254 95108 373260
rect 100850 373280 100906 373289
rect 88338 373215 88394 373224
rect 151740 373250 151768 373623
rect 156510 373552 156566 373561
rect 156510 373487 156566 373496
rect 100850 373215 100852 373224
rect 88352 373182 88380 373215
rect 100904 373215 100906 373224
rect 151728 373244 151780 373250
rect 100852 373186 100904 373192
rect 151728 373186 151780 373192
rect 156524 373182 156552 373487
rect 88340 373176 88392 373182
rect 156512 373176 156564 373182
rect 88340 373118 88392 373124
rect 92386 373144 92442 373153
rect 92386 373079 92442 373088
rect 93674 373144 93730 373153
rect 156512 373118 156564 373124
rect 93674 373079 93676 373088
rect 84750 372600 84806 372609
rect 84750 372535 84752 372544
rect 84804 372535 84806 372544
rect 86774 372600 86830 372609
rect 86774 372535 86830 372544
rect 88062 372600 88118 372609
rect 88062 372535 88118 372544
rect 89350 372600 89406 372609
rect 89350 372535 89406 372544
rect 90914 372600 90970 372609
rect 90914 372535 90970 372544
rect 91558 372600 91614 372609
rect 91558 372535 91614 372544
rect 84752 372506 84804 372512
rect 86788 372502 86816 372535
rect 86776 372496 86828 372502
rect 79506 372464 79562 372473
rect 79506 372399 79562 372408
rect 84566 372464 84622 372473
rect 86776 372438 86828 372444
rect 84566 372399 84622 372408
rect 78310 372328 78366 372337
rect 78310 372263 78366 372272
rect 76838 371784 76894 371793
rect 76838 371719 76894 371728
rect 77206 371784 77262 371793
rect 77206 371719 77262 371728
rect 76852 369578 76880 371719
rect 76840 369572 76892 369578
rect 76840 369514 76892 369520
rect 77220 369442 77248 371719
rect 78324 371482 78352 372263
rect 79520 372230 79548 372399
rect 79508 372224 79560 372230
rect 79508 372166 79560 372172
rect 78312 371476 78364 371482
rect 78312 371418 78364 371424
rect 79520 371346 79548 372166
rect 81438 372056 81494 372065
rect 81438 371991 81494 372000
rect 80060 371408 80112 371414
rect 80058 371376 80060 371385
rect 80112 371376 80114 371385
rect 79508 371340 79560 371346
rect 80058 371311 80114 371320
rect 79508 371282 79560 371288
rect 81452 371278 81480 371991
rect 83830 371512 83886 371521
rect 83830 371447 83886 371456
rect 81440 371272 81492 371278
rect 81440 371214 81492 371220
rect 77208 369436 77260 369442
rect 77208 369378 77260 369384
rect 83844 369102 83872 371447
rect 84580 371278 84608 372399
rect 88076 371686 88104 372535
rect 88064 371680 88116 371686
rect 88064 371622 88116 371628
rect 89364 371550 89392 372535
rect 90928 371618 90956 372535
rect 91572 372434 91600 372535
rect 91560 372428 91612 372434
rect 91560 372370 91612 372376
rect 92400 372366 92428 373079
rect 93728 373079 93730 373088
rect 93676 373050 93728 373056
rect 100024 372836 100076 372842
rect 100024 372778 100076 372784
rect 100036 372609 100064 372778
rect 93398 372600 93454 372609
rect 93398 372535 93454 372544
rect 100022 372600 100078 372609
rect 100022 372535 100078 372544
rect 104622 372600 104678 372609
rect 104622 372535 104678 372544
rect 112994 372600 113050 372609
rect 112994 372535 113050 372544
rect 114466 372600 114522 372609
rect 114466 372535 114522 372544
rect 92388 372360 92440 372366
rect 92388 372302 92440 372308
rect 93412 372298 93440 372535
rect 93400 372292 93452 372298
rect 93400 372234 93452 372240
rect 102046 371648 102102 371657
rect 90916 371612 90968 371618
rect 102046 371583 102102 371592
rect 90916 371554 90968 371560
rect 89352 371544 89404 371550
rect 89352 371486 89404 371492
rect 101678 371376 101734 371385
rect 101678 371311 101734 371320
rect 84568 371272 84620 371278
rect 84568 371214 84620 371220
rect 83832 369096 83884 369102
rect 83832 369038 83884 369044
rect 101692 368966 101720 371311
rect 102060 369170 102088 371583
rect 102782 371376 102838 371385
rect 102782 371311 102838 371320
rect 102048 369164 102100 369170
rect 102048 369106 102100 369112
rect 101680 368960 101732 368966
rect 101680 368902 101732 368908
rect 102796 368898 102824 371311
rect 104636 371074 104664 372535
rect 110142 372328 110198 372337
rect 110142 372263 110198 372272
rect 107014 371648 107070 371657
rect 107014 371583 107070 371592
rect 108854 371648 108910 371657
rect 108854 371583 108910 371592
rect 105634 371376 105690 371385
rect 105634 371311 105690 371320
rect 104624 371068 104676 371074
rect 104624 371010 104676 371016
rect 102784 368892 102836 368898
rect 102784 368834 102836 368840
rect 105648 368830 105676 371311
rect 106188 371272 106240 371278
rect 106188 371214 106240 371220
rect 106200 370394 106228 371214
rect 106188 370388 106240 370394
rect 106188 370330 106240 370336
rect 107028 369073 107056 371583
rect 108868 369374 108896 371583
rect 110156 370569 110184 372263
rect 113008 372026 113036 372535
rect 112996 372020 113048 372026
rect 112996 371962 113048 371968
rect 114480 371754 114508 372535
rect 114468 371748 114520 371754
rect 114468 371690 114520 371696
rect 111614 371648 111670 371657
rect 111614 371583 111670 371592
rect 110142 370560 110198 370569
rect 110142 370495 110198 370504
rect 108856 369368 108908 369374
rect 108856 369310 108908 369316
rect 111628 369306 111656 371583
rect 111616 369300 111668 369306
rect 111616 369242 111668 369248
rect 107014 369064 107070 369073
rect 107014 368999 107070 369008
rect 105636 368824 105688 368830
rect 105636 368766 105688 368772
rect 179340 351966 179368 374575
rect 182730 372464 182786 372473
rect 182730 372399 182786 372408
rect 182744 371822 182772 372399
rect 183282 371920 183338 371929
rect 183282 371855 183338 371864
rect 182732 371816 182784 371822
rect 182732 371758 182784 371764
rect 182744 371142 182772 371758
rect 183296 371210 183324 371855
rect 183284 371204 183336 371210
rect 183284 371146 183336 371152
rect 182732 371136 182784 371142
rect 182732 371078 182784 371084
rect 196636 370666 196664 495023
rect 196728 371006 196756 495037
rect 196820 495023 197110 495051
rect 196716 371000 196768 371006
rect 196716 370942 196768 370948
rect 196820 370734 196848 495023
rect 197572 494834 197600 495037
rect 197648 495023 198030 495051
rect 198108 495023 198490 495051
rect 197560 494828 197612 494834
rect 197560 494770 197612 494776
rect 197648 492538 197676 495023
rect 197464 492510 197676 492538
rect 196992 492176 197044 492182
rect 196992 492118 197044 492124
rect 196900 460284 196952 460290
rect 196900 460226 196952 460232
rect 196808 370728 196860 370734
rect 196808 370670 196860 370676
rect 196624 370660 196676 370666
rect 196624 370602 196676 370608
rect 179328 351960 179380 351966
rect 179326 351928 179328 351937
rect 179380 351928 179382 351937
rect 179326 351863 179382 351872
rect 191288 351212 191340 351218
rect 191288 351154 191340 351160
rect 179696 350600 179748 350606
rect 179694 350568 179696 350577
rect 191300 350577 191328 351154
rect 196636 350606 196664 350637
rect 196624 350600 196676 350606
rect 179748 350568 179750 350577
rect 179694 350503 179750 350512
rect 191286 350568 191342 350577
rect 191286 350503 191342 350512
rect 196622 350568 196624 350577
rect 196676 350568 196678 350577
rect 196622 350503 196678 350512
rect 62120 348696 62172 348702
rect 62120 348638 62172 348644
rect 110972 264920 111024 264926
rect 110970 264888 110972 264897
rect 111024 264888 111026 264897
rect 110970 264823 111026 264832
rect 125966 264888 126022 264897
rect 125966 264823 125968 264832
rect 126020 264823 126022 264832
rect 128358 264888 128414 264897
rect 128358 264823 128414 264832
rect 130934 264888 130990 264897
rect 130934 264823 130990 264832
rect 133418 264888 133474 264897
rect 133418 264823 133474 264832
rect 135902 264888 135958 264897
rect 135902 264823 135958 264832
rect 138478 264888 138534 264897
rect 138478 264823 138534 264832
rect 125968 264794 126020 264800
rect 128372 264722 128400 264823
rect 130948 264790 130976 264823
rect 130936 264784 130988 264790
rect 130936 264726 130988 264732
rect 128360 264716 128412 264722
rect 128360 264658 128412 264664
rect 133432 264654 133460 264823
rect 133420 264648 133472 264654
rect 133420 264590 133472 264596
rect 135916 264586 135944 264823
rect 135904 264580 135956 264586
rect 135904 264522 135956 264528
rect 138492 264518 138520 264823
rect 140870 264752 140926 264761
rect 140870 264687 140926 264696
rect 143538 264752 143594 264761
rect 143538 264687 143594 264696
rect 145930 264752 145986 264761
rect 145930 264687 145986 264696
rect 148506 264752 148562 264761
rect 148506 264687 148562 264696
rect 138480 264512 138532 264518
rect 138480 264454 138532 264460
rect 140884 264382 140912 264687
rect 143552 264450 143580 264687
rect 143540 264444 143592 264450
rect 143540 264386 143592 264392
rect 140872 264376 140924 264382
rect 140872 264318 140924 264324
rect 145944 264314 145972 264687
rect 145932 264308 145984 264314
rect 145932 264250 145984 264256
rect 148520 264246 148548 264687
rect 148508 264240 148560 264246
rect 60738 264208 60794 264217
rect 148508 264182 148560 264188
rect 60738 264143 60794 264152
rect 62212 264172 62264 264178
rect 60752 239970 60780 264143
rect 62212 264114 62264 264120
rect 62120 264104 62172 264110
rect 62120 264046 62172 264052
rect 62132 263634 62160 264046
rect 62224 263770 62252 264114
rect 62212 263764 62264 263770
rect 62212 263706 62264 263712
rect 89996 263764 90048 263770
rect 89996 263706 90048 263712
rect 62120 263628 62172 263634
rect 62120 263570 62172 263576
rect 60740 239964 60792 239970
rect 60740 239906 60792 239912
rect 60648 239624 60700 239630
rect 60648 239566 60700 239572
rect 60660 238610 60688 239566
rect 62132 239290 62160 263570
rect 62224 240038 62252 263706
rect 62304 263696 62356 263702
rect 62304 263638 62356 263644
rect 62316 240106 62344 263638
rect 90008 263537 90036 263706
rect 92388 263696 92440 263702
rect 92388 263638 92440 263644
rect 91284 263628 91336 263634
rect 91284 263570 91336 263576
rect 91296 263537 91324 263570
rect 92400 263537 92428 263638
rect 120908 263560 120960 263566
rect 80058 263528 80114 263537
rect 80058 263463 80114 263472
rect 88338 263528 88394 263537
rect 88338 263463 88394 263472
rect 89994 263528 90050 263537
rect 89994 263463 90050 263472
rect 90730 263528 90786 263537
rect 90730 263463 90786 263472
rect 91282 263528 91338 263537
rect 91282 263463 91338 263472
rect 92386 263528 92442 263537
rect 92386 263463 92442 263472
rect 93582 263528 93638 263537
rect 93582 263463 93638 263472
rect 96066 263528 96122 263537
rect 96066 263463 96122 263472
rect 98090 263528 98146 263537
rect 98090 263463 98146 263472
rect 101034 263528 101090 263537
rect 101034 263463 101090 263472
rect 103518 263528 103574 263537
rect 103518 263463 103574 263472
rect 105634 263528 105690 263537
rect 105634 263463 105690 263472
rect 108210 263528 108266 263537
rect 108210 263463 108266 263472
rect 109314 263528 109370 263537
rect 109314 263463 109370 263472
rect 113362 263528 113418 263537
rect 113362 263463 113418 263472
rect 115938 263528 115994 263537
rect 115938 263463 115994 263472
rect 116214 263528 116270 263537
rect 116214 263463 116270 263472
rect 118054 263528 118110 263537
rect 118054 263463 118110 263472
rect 120906 263528 120908 263537
rect 155960 263560 156012 263566
rect 120960 263528 120962 263537
rect 120906 263463 120962 263472
rect 123482 263528 123538 263537
rect 123482 263463 123484 263472
rect 66258 262848 66314 262857
rect 66258 262783 66314 262792
rect 78678 262848 78734 262857
rect 78678 262783 78734 262792
rect 64880 260024 64932 260030
rect 64880 259966 64932 259972
rect 64892 241602 64920 259966
rect 64880 241596 64932 241602
rect 64880 241538 64932 241544
rect 66076 241528 66128 241534
rect 66272 241482 66300 262783
rect 77298 262304 77354 262313
rect 77298 262239 77354 262248
rect 66128 241476 66300 241482
rect 66076 241470 66300 241476
rect 66088 241454 66300 241470
rect 66272 241126 66300 241454
rect 77312 241194 77340 262239
rect 78692 241330 78720 262783
rect 78680 241324 78732 241330
rect 78680 241266 78732 241272
rect 80072 241262 80100 263463
rect 81438 263256 81494 263265
rect 81438 263191 81494 263200
rect 84750 263256 84806 263265
rect 84750 263191 84806 263200
rect 80150 262848 80206 262857
rect 80150 262783 80206 262792
rect 80164 260409 80192 262783
rect 80150 260400 80206 260409
rect 80150 260335 80206 260344
rect 81452 241398 81480 263191
rect 82082 263120 82138 263129
rect 82082 263055 82138 263064
rect 81440 241392 81492 241398
rect 81440 241334 81492 241340
rect 80060 241256 80112 241262
rect 80060 241198 80112 241204
rect 77300 241188 77352 241194
rect 77300 241130 77352 241136
rect 66260 241120 66312 241126
rect 66260 241062 66312 241068
rect 67548 240780 67600 240786
rect 67548 240722 67600 240728
rect 62304 240100 62356 240106
rect 62304 240042 62356 240048
rect 62212 240032 62264 240038
rect 62212 239974 62264 239980
rect 67560 239834 67588 240722
rect 67548 239828 67600 239834
rect 67548 239770 67600 239776
rect 82096 239766 82124 263055
rect 84198 262984 84254 262993
rect 84198 262919 84254 262928
rect 84212 260710 84240 262919
rect 84200 260704 84252 260710
rect 84200 260646 84252 260652
rect 84764 260642 84792 263191
rect 87602 262984 87658 262993
rect 87602 262919 87658 262928
rect 85946 262576 86002 262585
rect 85946 262511 86002 262520
rect 84752 260636 84804 260642
rect 84752 260578 84804 260584
rect 85960 260098 85988 262511
rect 87616 260574 87644 262919
rect 88352 262682 88380 263463
rect 88614 262984 88670 262993
rect 88614 262919 88670 262928
rect 88340 262676 88392 262682
rect 88340 262618 88392 262624
rect 87604 260568 87656 260574
rect 87604 260510 87656 260516
rect 88628 260506 88656 262919
rect 90744 262750 90772 263463
rect 93596 262818 93624 263463
rect 96080 262886 96108 263463
rect 96526 263256 96582 263265
rect 96582 263214 96660 263242
rect 96526 263191 96582 263200
rect 96068 262880 96120 262886
rect 96068 262822 96120 262828
rect 93584 262812 93636 262818
rect 93584 262754 93636 262760
rect 90732 262744 90784 262750
rect 90732 262686 90784 262692
rect 96528 262676 96580 262682
rect 96528 262618 96580 262624
rect 89720 262404 89772 262410
rect 89720 262346 89772 262352
rect 88616 260500 88668 260506
rect 88616 260442 88668 260448
rect 89732 260438 89760 262346
rect 89720 260432 89772 260438
rect 89720 260374 89772 260380
rect 96540 260273 96568 262618
rect 96526 260264 96582 260273
rect 96526 260199 96582 260208
rect 85948 260092 86000 260098
rect 85948 260034 86000 260040
rect 96632 241126 96660 263214
rect 98104 262954 98132 263463
rect 99470 263256 99526 263265
rect 99470 263191 99526 263200
rect 98092 262948 98144 262954
rect 98092 262890 98144 262896
rect 97906 262304 97962 262313
rect 99286 262304 99342 262313
rect 97962 262262 98040 262290
rect 97906 262239 97962 262248
rect 96620 241120 96672 241126
rect 96620 241062 96672 241068
rect 98012 240786 98040 262262
rect 99342 262262 99420 262290
rect 99286 262239 99342 262248
rect 99392 241466 99420 262262
rect 99484 260302 99512 263191
rect 101048 263022 101076 263463
rect 103532 263090 103560 263463
rect 105648 263158 105676 263463
rect 108224 263226 108252 263463
rect 108212 263220 108264 263226
rect 108212 263162 108264 263168
rect 105636 263152 105688 263158
rect 105636 263094 105688 263100
rect 103520 263084 103572 263090
rect 103520 263026 103572 263032
rect 101036 263016 101088 263022
rect 100758 262984 100814 262993
rect 101036 262958 101088 262964
rect 100758 262919 100814 262928
rect 100024 262472 100076 262478
rect 100024 262414 100076 262420
rect 99472 260296 99524 260302
rect 99472 260238 99524 260244
rect 99380 241460 99432 241466
rect 99380 241402 99432 241408
rect 98000 240780 98052 240786
rect 98000 240722 98052 240728
rect 82084 239760 82136 239766
rect 82084 239702 82136 239708
rect 100036 239698 100064 262414
rect 100772 260778 100800 262919
rect 101770 262712 101826 262721
rect 101770 262647 101772 262656
rect 101824 262647 101826 262656
rect 102322 262712 102378 262721
rect 102322 262647 102378 262656
rect 105082 262712 105138 262721
rect 105082 262647 105138 262656
rect 108026 262712 108082 262721
rect 108026 262647 108082 262656
rect 101772 262618 101824 262624
rect 100760 260772 100812 260778
rect 100760 260714 100812 260720
rect 102336 260370 102364 262647
rect 102324 260364 102376 260370
rect 102324 260306 102376 260312
rect 105096 260234 105124 262647
rect 107566 262440 107622 262449
rect 107622 262398 107792 262426
rect 107566 262375 107622 262384
rect 107566 262304 107622 262313
rect 107622 262262 107700 262290
rect 107566 262239 107622 262248
rect 105084 260228 105136 260234
rect 105084 260170 105136 260176
rect 100024 239692 100076 239698
rect 100024 239634 100076 239640
rect 107672 239630 107700 262262
rect 107660 239624 107712 239630
rect 107660 239566 107712 239572
rect 107764 239562 107792 262398
rect 108040 260166 108068 262647
rect 109328 262410 109356 263463
rect 113376 263294 113404 263463
rect 115952 263430 115980 263463
rect 115940 263424 115992 263430
rect 114374 263392 114430 263401
rect 115940 263366 115992 263372
rect 114374 263327 114430 263336
rect 113364 263288 113416 263294
rect 113364 263230 113416 263236
rect 114388 262886 114416 263327
rect 114376 262880 114428 262886
rect 114376 262822 114428 262828
rect 114650 262576 114706 262585
rect 114650 262511 114706 262520
rect 109316 262404 109368 262410
rect 109316 262346 109368 262352
rect 110418 262304 110474 262313
rect 110418 262239 110474 262248
rect 113178 262304 113234 262313
rect 113178 262239 113234 262248
rect 108028 260160 108080 260166
rect 108028 260102 108080 260108
rect 107752 239556 107804 239562
rect 107752 239498 107804 239504
rect 110432 239494 110460 262239
rect 110420 239488 110472 239494
rect 110420 239430 110472 239436
rect 113192 239426 113220 262239
rect 114664 260137 114692 262511
rect 116228 262478 116256 263463
rect 118068 263362 118096 263463
rect 123536 263463 123538 263472
rect 150990 263528 151046 263537
rect 150990 263463 151046 263472
rect 155958 263528 155960 263537
rect 156012 263528 156014 263537
rect 155958 263463 156014 263472
rect 158534 263528 158590 263537
rect 158534 263463 158536 263472
rect 123484 263434 123536 263440
rect 151004 263430 151032 263463
rect 158588 263463 158590 263472
rect 161110 263528 161166 263537
rect 161110 263463 161166 263472
rect 163502 263528 163558 263537
rect 163502 263463 163558 263472
rect 166078 263528 166134 263537
rect 166078 263463 166134 263472
rect 158536 263434 158588 263440
rect 150992 263424 151044 263430
rect 150992 263366 151044 263372
rect 161124 263362 161152 263463
rect 118056 263356 118108 263362
rect 118056 263298 118108 263304
rect 161112 263356 161164 263362
rect 161112 263298 161164 263304
rect 163516 263226 163544 263463
rect 166092 263294 166120 263463
rect 166080 263288 166132 263294
rect 166080 263230 166132 263236
rect 163504 263220 163556 263226
rect 163504 263162 163556 263168
rect 183376 263016 183428 263022
rect 118698 262984 118754 262993
rect 183376 262958 183428 262964
rect 118698 262919 118754 262928
rect 116216 262472 116268 262478
rect 116216 262414 116268 262420
rect 118712 260846 118740 262919
rect 183388 262313 183416 262958
rect 183468 262948 183520 262954
rect 183468 262890 183520 262896
rect 183480 262449 183508 262890
rect 183466 262440 183522 262449
rect 183466 262375 183522 262384
rect 183374 262304 183430 262313
rect 183374 262239 183430 262248
rect 118700 260840 118752 260846
rect 118700 260782 118752 260788
rect 114650 260128 114706 260137
rect 114650 260063 114706 260072
rect 180156 241052 180208 241058
rect 180156 240994 180208 241000
rect 179328 240916 179380 240922
rect 179328 240858 179380 240864
rect 179340 240281 179368 240858
rect 180168 240281 180196 240994
rect 183388 240990 183416 262239
rect 183376 240984 183428 240990
rect 183376 240926 183428 240932
rect 183480 240854 183508 262375
rect 196636 241058 196664 350503
rect 196912 262886 196940 460226
rect 197004 370598 197032 492118
rect 197360 491904 197412 491910
rect 197360 491846 197412 491852
rect 197372 491609 197400 491846
rect 197358 491600 197414 491609
rect 197358 491535 197414 491544
rect 197084 466132 197136 466138
rect 197084 466074 197136 466080
rect 197096 374270 197124 466074
rect 197084 374264 197136 374270
rect 197084 374206 197136 374212
rect 197464 370870 197492 492510
rect 198108 492402 198136 495023
rect 198860 494850 198888 495037
rect 199120 495023 199318 495051
rect 199488 495023 199778 495051
rect 200254 495023 200344 495051
rect 198280 494828 198332 494834
rect 198860 494822 199056 494850
rect 198280 494770 198332 494776
rect 197556 492374 198136 492402
rect 197556 371142 197584 492374
rect 197636 492040 197688 492046
rect 197636 491982 197688 491988
rect 197648 491745 197676 491982
rect 198096 491836 198148 491842
rect 198096 491778 198148 491784
rect 197634 491736 197690 491745
rect 197634 491671 197690 491680
rect 197728 491700 197780 491706
rect 197728 491642 197780 491648
rect 197740 491337 197768 491642
rect 197726 491328 197782 491337
rect 197726 491263 197782 491272
rect 197820 466200 197872 466206
rect 197820 466142 197872 466148
rect 197636 463004 197688 463010
rect 197636 462946 197688 462952
rect 197544 371136 197596 371142
rect 197544 371078 197596 371084
rect 197452 370864 197504 370870
rect 197452 370806 197504 370812
rect 196992 370592 197044 370598
rect 196992 370534 197044 370540
rect 197648 263430 197676 462946
rect 197728 460488 197780 460494
rect 197728 460430 197780 460436
rect 197636 263424 197688 263430
rect 197636 263366 197688 263372
rect 197740 263226 197768 460430
rect 197832 373250 197860 466142
rect 198004 459128 198056 459134
rect 198004 459070 198056 459076
rect 197912 458992 197964 458998
rect 197912 458934 197964 458940
rect 197924 373590 197952 458934
rect 198016 374542 198044 459070
rect 198004 374536 198056 374542
rect 198004 374478 198056 374484
rect 197912 373584 197964 373590
rect 197912 373526 197964 373532
rect 197820 373244 197872 373250
rect 197820 373186 197872 373192
rect 198004 273964 198056 273970
rect 198004 273906 198056 273912
rect 197728 263220 197780 263226
rect 197728 263162 197780 263168
rect 196900 262880 196952 262886
rect 196900 262822 196952 262828
rect 196912 258074 196940 262822
rect 196820 258046 196940 258074
rect 196716 242140 196768 242146
rect 196716 242082 196768 242088
rect 196624 241052 196676 241058
rect 196624 240994 196676 241000
rect 183468 240848 183520 240854
rect 183468 240790 183520 240796
rect 179326 240272 179382 240281
rect 179326 240207 179382 240216
rect 180154 240272 180210 240281
rect 180154 240207 180210 240216
rect 190918 240272 190974 240281
rect 190918 240207 190920 240216
rect 190972 240207 190974 240216
rect 190920 240178 190972 240184
rect 113180 239420 113232 239426
rect 113180 239362 113232 239368
rect 62120 239284 62172 239290
rect 62120 239226 62172 239232
rect 60648 238604 60700 238610
rect 60648 238546 60700 238552
rect 96066 154728 96122 154737
rect 96066 154663 96122 154672
rect 113362 154728 113418 154737
rect 113362 154663 113418 154672
rect 163318 154728 163374 154737
rect 163318 154663 163320 154672
rect 96080 154494 96108 154663
rect 96068 154488 96120 154494
rect 96068 154430 96120 154436
rect 98460 154420 98512 154426
rect 98460 154362 98512 154368
rect 98472 154193 98500 154362
rect 101036 154352 101088 154358
rect 101036 154294 101088 154300
rect 101048 154193 101076 154294
rect 105820 154284 105872 154290
rect 105820 154226 105872 154232
rect 105832 154193 105860 154226
rect 98458 154184 98514 154193
rect 98458 154119 98514 154128
rect 101034 154184 101090 154193
rect 101034 154119 101090 154128
rect 105818 154184 105874 154193
rect 105818 154119 105874 154128
rect 108210 154184 108266 154193
rect 113376 154154 113404 154663
rect 163372 154663 163374 154672
rect 165894 154728 165950 154737
rect 165894 154663 165950 154672
rect 163320 154634 163372 154640
rect 165908 154630 165936 154663
rect 165896 154624 165948 154630
rect 165896 154566 165948 154572
rect 138386 154320 138442 154329
rect 138386 154255 138442 154264
rect 138400 154222 138428 154255
rect 138388 154216 138440 154222
rect 138388 154158 138440 154164
rect 143538 154184 143594 154193
rect 108210 154119 108212 154128
rect 108264 154119 108266 154128
rect 113364 154148 113416 154154
rect 108212 154090 108264 154096
rect 113364 154090 113416 154096
rect 114468 154148 114520 154154
rect 143538 154119 143594 154128
rect 114468 154090 114520 154096
rect 60004 153944 60056 153950
rect 60004 153886 60056 153892
rect 111156 153400 111208 153406
rect 111156 153342 111208 153348
rect 111168 153105 111196 153342
rect 114480 153218 114508 154090
rect 143552 154086 143580 154119
rect 143540 154080 143592 154086
rect 143540 154022 143592 154028
rect 145930 154048 145986 154057
rect 145930 153983 145932 153992
rect 145984 153983 145986 153992
rect 150898 154048 150954 154057
rect 150898 153983 150954 153992
rect 145932 153954 145984 153960
rect 150912 153950 150940 153983
rect 150900 153944 150952 153950
rect 150900 153886 150952 153892
rect 153290 153912 153346 153921
rect 153290 153847 153292 153856
rect 153344 153847 153346 153856
rect 153292 153818 153344 153824
rect 118700 153332 118752 153338
rect 118700 153274 118752 153280
rect 114744 153264 114796 153270
rect 114480 153190 114692 153218
rect 114744 153206 114796 153212
rect 75918 153096 75974 153105
rect 75918 153031 75974 153040
rect 77298 153096 77354 153105
rect 77298 153031 77354 153040
rect 78678 153096 78734 153105
rect 78678 153031 78734 153040
rect 81438 153096 81494 153105
rect 81438 153031 81494 153040
rect 82818 153096 82874 153105
rect 82818 153031 82874 153040
rect 84198 153096 84254 153105
rect 84198 153031 84254 153040
rect 85578 153096 85634 153105
rect 85578 153031 85634 153040
rect 86958 153096 87014 153105
rect 86958 153031 87014 153040
rect 88430 153096 88486 153105
rect 88430 153031 88486 153040
rect 89810 153096 89866 153105
rect 89810 153031 89866 153040
rect 91098 153096 91154 153105
rect 91098 153031 91154 153040
rect 92478 153096 92534 153105
rect 92478 153031 92534 153040
rect 93858 153096 93914 153105
rect 93858 153031 93914 153040
rect 95238 153096 95294 153105
rect 95238 153031 95294 153040
rect 96618 153096 96674 153105
rect 96618 153031 96674 153040
rect 97998 153096 98054 153105
rect 97998 153031 98054 153040
rect 99378 153096 99434 153105
rect 99378 153031 99434 153040
rect 100850 153096 100906 153105
rect 100850 153031 100906 153040
rect 102138 153096 102194 153105
rect 102138 153031 102194 153040
rect 103610 153096 103666 153105
rect 103610 153031 103666 153040
rect 106370 153096 106426 153105
rect 106370 153031 106426 153040
rect 109038 153096 109094 153105
rect 109038 153031 109094 153040
rect 110418 153096 110474 153105
rect 110418 153031 110474 153040
rect 111154 153096 111210 153105
rect 111154 153031 111210 153040
rect 111798 153096 111854 153105
rect 111798 153031 111854 153040
rect 114558 153096 114614 153105
rect 114558 153031 114614 153040
rect 60004 151360 60056 151366
rect 60004 151302 60056 151308
rect 60016 150686 60044 151302
rect 60004 150680 60056 150686
rect 60004 150622 60056 150628
rect 59912 133340 59964 133346
rect 59912 133282 59964 133288
rect 59820 131096 59872 131102
rect 59820 131038 59872 131044
rect 59360 81456 59412 81462
rect 59360 81398 59412 81404
rect 59832 43994 59860 131038
rect 59820 43988 59872 43994
rect 59820 43930 59872 43936
rect 59924 42294 59952 133282
rect 59912 42288 59964 42294
rect 59912 42230 59964 42236
rect 60016 41070 60044 150622
rect 75932 130218 75960 153031
rect 76010 152552 76066 152561
rect 76010 152487 76066 152496
rect 76024 130286 76052 152487
rect 77312 130354 77340 153031
rect 78692 133482 78720 153031
rect 80058 152008 80114 152017
rect 80058 151943 80114 151952
rect 80072 133550 80100 151943
rect 80060 133544 80112 133550
rect 80060 133486 80112 133492
rect 78680 133476 78732 133482
rect 78680 133418 78732 133424
rect 81452 133414 81480 153031
rect 81440 133408 81492 133414
rect 81440 133350 81492 133356
rect 82832 130626 82860 153031
rect 84212 130898 84240 153031
rect 84290 152008 84346 152017
rect 84290 151943 84346 151952
rect 84200 130892 84252 130898
rect 84200 130834 84252 130840
rect 82820 130620 82872 130626
rect 82820 130562 82872 130568
rect 84304 130558 84332 151943
rect 85592 130830 85620 153031
rect 85580 130824 85632 130830
rect 85580 130766 85632 130772
rect 84292 130552 84344 130558
rect 84292 130494 84344 130500
rect 86972 130490 87000 153031
rect 88338 152416 88394 152425
rect 88338 152351 88394 152360
rect 88352 152318 88380 152351
rect 88340 152312 88392 152318
rect 88340 152254 88392 152260
rect 88444 130966 88472 153031
rect 88890 152824 88946 152833
rect 88890 152759 88946 152768
rect 88904 152561 88932 152759
rect 88890 152552 88946 152561
rect 88890 152487 88946 152496
rect 89718 152416 89774 152425
rect 89718 152351 89720 152360
rect 89772 152351 89774 152360
rect 89720 152322 89772 152328
rect 88432 130960 88484 130966
rect 88432 130902 88484 130908
rect 89824 130694 89852 153031
rect 91112 131034 91140 153031
rect 91190 152824 91246 152833
rect 91190 152759 91246 152768
rect 91100 131028 91152 131034
rect 91100 130970 91152 130976
rect 91204 130762 91232 152759
rect 91192 130756 91244 130762
rect 91192 130698 91244 130704
rect 89812 130688 89864 130694
rect 89812 130630 89864 130636
rect 86960 130484 87012 130490
rect 86960 130426 87012 130432
rect 92492 130422 92520 153031
rect 93872 131102 93900 153031
rect 93860 131096 93912 131102
rect 93860 131038 93912 131044
rect 95252 130529 95280 153031
rect 96632 151434 96660 153031
rect 97264 152380 97316 152386
rect 97264 152322 97316 152328
rect 96620 151428 96672 151434
rect 96620 151370 96672 151376
rect 97276 130665 97304 152322
rect 98012 151638 98040 153031
rect 98644 151904 98696 151910
rect 98644 151846 98696 151852
rect 98000 151632 98052 151638
rect 98000 151574 98052 151580
rect 98656 133113 98684 151846
rect 98642 133104 98698 133113
rect 98642 133039 98698 133048
rect 97262 130656 97318 130665
rect 97262 130591 97318 130600
rect 95238 130520 95294 130529
rect 95238 130455 95294 130464
rect 92480 130416 92532 130422
rect 99392 130393 99420 153031
rect 100758 152824 100814 152833
rect 100758 152759 100814 152768
rect 100772 152386 100800 152759
rect 100760 152380 100812 152386
rect 100760 152322 100812 152328
rect 100864 151298 100892 153031
rect 100852 151292 100904 151298
rect 100852 151234 100904 151240
rect 102152 131073 102180 153031
rect 103518 152824 103574 152833
rect 103518 152759 103574 152768
rect 103532 152454 103560 152759
rect 103520 152448 103572 152454
rect 103520 152390 103572 152396
rect 103624 133822 103652 153031
rect 106278 152824 106334 152833
rect 106278 152759 106334 152768
rect 104898 152144 104954 152153
rect 104898 152079 104954 152088
rect 104912 151910 104940 152079
rect 104900 151904 104952 151910
rect 104900 151846 104952 151852
rect 106292 151230 106320 152759
rect 106384 151366 106412 153031
rect 106372 151360 106424 151366
rect 106372 151302 106424 151308
rect 106280 151224 106332 151230
rect 106280 151166 106332 151172
rect 103612 133816 103664 133822
rect 103612 133758 103664 133764
rect 109052 133346 109080 153031
rect 109130 152824 109186 152833
rect 109130 152759 109186 152768
rect 109144 151162 109172 152759
rect 110432 151706 110460 153031
rect 110420 151700 110472 151706
rect 110420 151642 110472 151648
rect 109132 151156 109184 151162
rect 109132 151098 109184 151104
rect 111812 151094 111840 153031
rect 113178 152824 113234 152833
rect 113178 152759 113234 152768
rect 113192 152590 113220 152759
rect 113180 152584 113232 152590
rect 113180 152526 113232 152532
rect 111800 151088 111852 151094
rect 111800 151030 111852 151036
rect 109040 133340 109092 133346
rect 109040 133282 109092 133288
rect 114572 133278 114600 153031
rect 114560 133272 114612 133278
rect 114560 133214 114612 133220
rect 114664 133210 114692 153190
rect 114756 153105 114784 153206
rect 118712 153105 118740 153274
rect 155960 153196 156012 153202
rect 155960 153138 156012 153144
rect 135260 153128 135312 153134
rect 114742 153096 114798 153105
rect 114742 153031 114798 153040
rect 117318 153096 117374 153105
rect 117318 153031 117374 153040
rect 117502 153096 117558 153105
rect 117502 153031 117558 153040
rect 118698 153096 118754 153105
rect 118698 153031 118754 153040
rect 125598 153096 125654 153105
rect 125598 153031 125654 153040
rect 128358 153096 128414 153105
rect 128358 153031 128414 153040
rect 129738 153096 129794 153105
rect 129738 153031 129794 153040
rect 132774 153096 132830 153105
rect 132774 153031 132776 153040
rect 115938 152552 115994 152561
rect 115938 152487 115940 152496
rect 115992 152487 115994 152496
rect 115940 152458 115992 152464
rect 117332 133890 117360 153031
rect 117410 152824 117466 152833
rect 117410 152759 117466 152768
rect 117424 151774 117452 152759
rect 117516 152658 117544 153031
rect 125612 152862 125640 153031
rect 128372 152930 128400 153031
rect 129752 152998 129780 153031
rect 132828 153031 132830 153040
rect 135258 153096 135260 153105
rect 155972 153105 156000 153138
rect 135312 153096 135314 153105
rect 135258 153031 135314 153040
rect 155958 153096 156014 153105
rect 155958 153031 156014 153040
rect 132776 153002 132828 153008
rect 129740 152992 129792 152998
rect 129740 152934 129792 152940
rect 128360 152924 128412 152930
rect 128360 152866 128412 152872
rect 125600 152856 125652 152862
rect 120078 152824 120134 152833
rect 120078 152759 120134 152768
rect 122838 152824 122894 152833
rect 125600 152798 125652 152804
rect 183466 152824 183522 152833
rect 122838 152759 122840 152768
rect 120092 152726 120120 152759
rect 122892 152759 122894 152768
rect 183466 152759 183522 152768
rect 122840 152730 122892 152736
rect 120080 152720 120132 152726
rect 120080 152662 120132 152668
rect 183480 152658 183508 152759
rect 117504 152652 117556 152658
rect 117504 152594 117556 152600
rect 183468 152652 183520 152658
rect 183468 152594 183520 152600
rect 183466 152552 183522 152561
rect 183466 152487 183468 152496
rect 183520 152487 183522 152496
rect 183468 152458 183520 152464
rect 117412 151768 117464 151774
rect 117412 151710 117464 151716
rect 117320 133884 117372 133890
rect 117320 133826 117372 133832
rect 114652 133204 114704 133210
rect 114652 133146 114704 133152
rect 179052 131096 179104 131102
rect 102138 131064 102194 131073
rect 179052 131038 179104 131044
rect 102138 130999 102194 131008
rect 92480 130358 92532 130364
rect 99378 130384 99434 130393
rect 77300 130348 77352 130354
rect 99378 130319 99434 130328
rect 77300 130290 77352 130296
rect 76012 130280 76064 130286
rect 76012 130222 76064 130228
rect 75920 130212 75972 130218
rect 75920 130154 75972 130160
rect 179064 129849 179092 131038
rect 179788 131028 179840 131034
rect 179788 130970 179840 130976
rect 179800 129849 179828 130970
rect 183480 130490 183508 152458
rect 191748 131164 191800 131170
rect 191748 131106 191800 131112
rect 183468 130484 183520 130490
rect 183468 130426 183520 130432
rect 191760 130393 191788 131106
rect 196636 131034 196664 240994
rect 196728 240922 196756 242082
rect 196716 240916 196768 240922
rect 196716 240858 196768 240864
rect 196728 131102 196756 240858
rect 196820 154154 196848 258046
rect 198016 240242 198044 273906
rect 198004 240236 198056 240242
rect 198004 240178 198056 240184
rect 198016 163538 198044 240178
rect 198004 163532 198056 163538
rect 198004 163474 198056 163480
rect 196808 154148 196860 154154
rect 196808 154090 196860 154096
rect 197360 153264 197412 153270
rect 197360 153206 197412 153212
rect 197372 152658 197400 153206
rect 197360 152652 197412 152658
rect 197360 152594 197412 152600
rect 196716 131096 196768 131102
rect 196716 131038 196768 131044
rect 196624 131028 196676 131034
rect 196624 130970 196676 130976
rect 191746 130384 191802 130393
rect 191746 130319 191802 130328
rect 179050 129840 179106 129849
rect 179050 129775 179106 129784
rect 179786 129840 179842 129849
rect 179786 129775 179842 129784
rect 77114 44840 77170 44849
rect 77114 44775 77170 44784
rect 83094 44840 83150 44849
rect 83094 44775 83150 44784
rect 84198 44840 84254 44849
rect 84198 44775 84254 44784
rect 94502 44840 94558 44849
rect 94502 44775 94558 44784
rect 96986 44840 97042 44849
rect 96986 44775 97042 44784
rect 98090 44840 98146 44849
rect 98090 44775 98146 44784
rect 77128 44538 77156 44775
rect 77116 44532 77168 44538
rect 77116 44474 77168 44480
rect 83108 44470 83136 44775
rect 83096 44464 83148 44470
rect 83096 44406 83148 44412
rect 84212 44062 84240 44775
rect 84200 44056 84252 44062
rect 84200 43998 84252 44004
rect 94516 43994 94544 44775
rect 94504 43988 94556 43994
rect 94504 43930 94556 43936
rect 97000 43926 97028 44775
rect 96988 43920 97040 43926
rect 96988 43862 97040 43868
rect 98104 43858 98132 44775
rect 100758 44704 100814 44713
rect 100758 44639 100814 44648
rect 101770 44704 101826 44713
rect 101770 44639 101826 44648
rect 102782 44704 102838 44713
rect 102782 44639 102838 44648
rect 103886 44704 103942 44713
rect 103886 44639 103942 44648
rect 143538 44704 143594 44713
rect 143538 44639 143594 44648
rect 145930 44704 145986 44713
rect 145930 44639 145986 44648
rect 100772 44334 100800 44639
rect 101784 44402 101812 44639
rect 101772 44396 101824 44402
rect 101772 44338 101824 44344
rect 100760 44328 100812 44334
rect 100760 44270 100812 44276
rect 98092 43852 98144 43858
rect 98092 43794 98144 43800
rect 102796 43790 102824 44639
rect 102784 43784 102836 43790
rect 102784 43726 102836 43732
rect 103900 43722 103928 44639
rect 113270 44568 113326 44577
rect 113270 44503 113326 44512
rect 103888 43716 103940 43722
rect 103888 43658 103940 43664
rect 113284 43654 113312 44503
rect 143552 44266 143580 44639
rect 143540 44260 143592 44266
rect 143540 44202 143592 44208
rect 145944 44198 145972 44639
rect 145932 44192 145984 44198
rect 145932 44134 145984 44140
rect 158442 44160 158498 44169
rect 158442 44095 158498 44104
rect 160834 44160 160890 44169
rect 160834 44095 160890 44104
rect 115938 43752 115994 43761
rect 115938 43687 115994 43696
rect 113272 43648 113324 43654
rect 113272 43590 113324 43596
rect 115952 43586 115980 43687
rect 115940 43580 115992 43586
rect 115940 43522 115992 43528
rect 158456 43518 158484 44095
rect 158444 43512 158496 43518
rect 158444 43454 158496 43460
rect 160848 43450 160876 44095
rect 160836 43444 160888 43450
rect 160836 43386 160888 43392
rect 85394 43208 85450 43217
rect 85394 43143 85450 43152
rect 92386 43208 92442 43217
rect 92386 43143 92442 43152
rect 95882 43208 95938 43217
rect 95882 43143 95938 43152
rect 128358 43208 128414 43217
rect 128358 43143 128414 43152
rect 76010 42800 76066 42809
rect 76010 42735 76066 42744
rect 78218 42800 78274 42809
rect 78218 42735 78274 42744
rect 80426 42800 80482 42809
rect 80426 42735 80482 42744
rect 76024 42090 76052 42735
rect 76012 42084 76064 42090
rect 76012 42026 76064 42032
rect 60004 41064 60056 41070
rect 60004 41006 60056 41012
rect 78232 40730 78260 42735
rect 78770 41848 78826 41857
rect 78770 41783 78826 41792
rect 78220 40724 78272 40730
rect 78220 40666 78272 40672
rect 59268 39500 59320 39506
rect 59268 39442 59320 39448
rect 78784 39370 78812 41783
rect 80440 40662 80468 42735
rect 81806 41848 81862 41857
rect 81806 41783 81862 41792
rect 80428 40656 80480 40662
rect 80428 40598 80480 40604
rect 81820 39438 81848 41783
rect 85408 41002 85436 43143
rect 86498 42800 86554 42809
rect 86498 42735 86554 42744
rect 87602 42800 87658 42809
rect 87602 42735 87658 42744
rect 88338 42800 88394 42809
rect 88338 42735 88394 42744
rect 88614 42800 88670 42809
rect 88614 42735 88670 42744
rect 90730 42800 90786 42809
rect 90730 42735 90786 42744
rect 91282 42800 91338 42809
rect 91282 42735 91338 42744
rect 85396 40996 85448 41002
rect 85396 40938 85448 40944
rect 86512 40934 86540 42735
rect 86500 40928 86552 40934
rect 86500 40870 86552 40876
rect 87616 40798 87644 42735
rect 88352 42158 88380 42735
rect 88340 42152 88392 42158
rect 88340 42094 88392 42100
rect 87604 40792 87656 40798
rect 87604 40734 87656 40740
rect 88628 39574 88656 42735
rect 89994 41848 90050 41857
rect 89994 41783 90050 41792
rect 88616 39568 88668 39574
rect 88616 39510 88668 39516
rect 90008 39506 90036 41783
rect 90744 39778 90772 42735
rect 90732 39772 90784 39778
rect 90732 39714 90784 39720
rect 91296 39710 91324 42735
rect 92400 40866 92428 43143
rect 93306 42800 93362 42809
rect 93306 42735 93362 42744
rect 93674 42800 93730 42809
rect 93674 42735 93730 42744
rect 92388 40860 92440 40866
rect 92388 40802 92440 40808
rect 91284 39704 91336 39710
rect 91284 39646 91336 39652
rect 93320 39642 93348 42735
rect 93688 41206 93716 42735
rect 95896 42226 95924 43143
rect 96250 42800 96306 42809
rect 96250 42735 96306 42744
rect 106370 42800 106426 42809
rect 106370 42735 106426 42744
rect 107014 42800 107070 42809
rect 107014 42735 107070 42744
rect 108578 42800 108634 42809
rect 108578 42735 108634 42744
rect 111890 42800 111946 42809
rect 111890 42735 111946 42744
rect 113178 42800 113234 42809
rect 113178 42735 113234 42744
rect 114190 42800 114246 42809
rect 114190 42735 114246 42744
rect 115754 42800 115810 42809
rect 115754 42735 115810 42744
rect 116306 42800 116362 42809
rect 116306 42735 116362 42744
rect 118238 42800 118294 42809
rect 118238 42735 118294 42744
rect 119066 42800 119122 42809
rect 119066 42735 119122 42744
rect 96264 42362 96292 42735
rect 96252 42356 96304 42362
rect 96252 42298 96304 42304
rect 95884 42220 95936 42226
rect 95884 42162 95936 42168
rect 93676 41200 93728 41206
rect 93676 41142 93728 41148
rect 106384 41070 106412 42735
rect 107028 41138 107056 42735
rect 108592 42294 108620 42735
rect 108580 42288 108632 42294
rect 108580 42230 108632 42236
rect 109314 42256 109370 42265
rect 109314 42191 109370 42200
rect 111154 42256 111210 42265
rect 111154 42191 111210 42200
rect 107016 41132 107068 41138
rect 107016 41074 107068 41080
rect 106372 41064 106424 41070
rect 106372 41006 106424 41012
rect 109328 39846 109356 42191
rect 111168 39914 111196 42191
rect 111904 39982 111932 42735
rect 113192 42430 113220 42735
rect 113180 42424 113232 42430
rect 113180 42366 113232 42372
rect 114204 41274 114232 42735
rect 115768 41410 115796 42735
rect 115756 41404 115808 41410
rect 115756 41346 115808 41352
rect 114192 41268 114244 41274
rect 114192 41210 114244 41216
rect 116320 40050 116348 42735
rect 118252 42498 118280 42735
rect 118240 42492 118292 42498
rect 118240 42434 118292 42440
rect 119080 41342 119108 42735
rect 128372 42566 128400 43143
rect 133418 42800 133474 42809
rect 133418 42735 133474 42744
rect 135902 42800 135958 42809
rect 135902 42735 135958 42744
rect 155958 42800 156014 42809
rect 155958 42735 155960 42744
rect 133432 42634 133460 42735
rect 135916 42702 135944 42735
rect 156012 42735 156014 42744
rect 183466 42800 183522 42809
rect 183466 42735 183468 42744
rect 155960 42706 156012 42712
rect 183520 42735 183522 42744
rect 183468 42706 183520 42712
rect 197372 42702 197400 152594
rect 198016 131170 198044 163474
rect 198108 154086 198136 491778
rect 198188 491768 198240 491774
rect 198188 491710 198240 491716
rect 198200 264625 198228 491710
rect 198292 370802 198320 494770
rect 199028 491366 199056 494822
rect 199016 491360 199068 491366
rect 199016 491302 199068 491308
rect 199120 491178 199148 495023
rect 198752 491150 199148 491178
rect 198646 375320 198702 375329
rect 198646 375255 198702 375264
rect 198280 370796 198332 370802
rect 198280 370738 198332 370744
rect 198186 264616 198242 264625
rect 198186 264551 198242 264560
rect 198096 154080 198148 154086
rect 198096 154022 198148 154028
rect 198004 131164 198056 131170
rect 198004 131106 198056 131112
rect 197452 130484 197504 130490
rect 197452 130426 197504 130432
rect 197464 42770 197492 130426
rect 198016 130422 198044 131106
rect 198004 130416 198056 130422
rect 198004 130358 198056 130364
rect 198660 43518 198688 375255
rect 198752 370530 198780 491150
rect 199488 489914 199516 495023
rect 200316 492046 200344 495023
rect 200408 495023 200698 495051
rect 200776 495023 201066 495051
rect 200304 492040 200356 492046
rect 200210 492008 200266 492017
rect 200304 491982 200356 491988
rect 200210 491943 200266 491952
rect 200224 491745 200252 491943
rect 200210 491736 200266 491745
rect 200210 491671 200266 491680
rect 200408 489914 200436 495023
rect 200672 492244 200724 492250
rect 200672 492186 200724 492192
rect 200684 492153 200712 492186
rect 200670 492144 200726 492153
rect 200670 492079 200726 492088
rect 200776 489914 200804 495023
rect 200856 492380 200908 492386
rect 200856 492322 200908 492328
rect 200868 492289 200896 492322
rect 200854 492280 200910 492289
rect 200854 492215 200910 492224
rect 198844 489886 199516 489914
rect 200224 489886 200436 489914
rect 200684 489886 200804 489914
rect 198844 371210 198872 489886
rect 198924 489456 198976 489462
rect 198924 489398 198976 489404
rect 198936 373726 198964 489398
rect 199200 480956 199252 480962
rect 199200 480898 199252 480904
rect 199108 463140 199160 463146
rect 199108 463082 199160 463088
rect 199016 460216 199068 460222
rect 199016 460158 199068 460164
rect 199028 458386 199056 460158
rect 199016 458380 199068 458386
rect 199016 458322 199068 458328
rect 199028 454753 199056 458322
rect 199014 454744 199070 454753
rect 199014 454679 199070 454688
rect 198924 373720 198976 373726
rect 198924 373662 198976 373668
rect 198832 371204 198884 371210
rect 198832 371146 198884 371152
rect 198740 370524 198792 370530
rect 198740 370466 198792 370472
rect 199028 345014 199056 454679
rect 199120 374610 199148 463082
rect 199212 394641 199240 480898
rect 199384 475380 199436 475386
rect 199384 475322 199436 475328
rect 199292 459060 199344 459066
rect 199292 459002 199344 459008
rect 199198 394632 199254 394641
rect 199198 394567 199254 394576
rect 199108 374604 199160 374610
rect 199108 374546 199160 374552
rect 199304 373794 199332 459002
rect 199396 391377 199424 475322
rect 199568 462324 199620 462330
rect 199568 462266 199620 462272
rect 199580 461718 199608 462266
rect 199476 461712 199528 461718
rect 199476 461654 199528 461660
rect 199568 461712 199620 461718
rect 199568 461654 199620 461660
rect 199382 391368 199438 391377
rect 199382 391303 199438 391312
rect 199292 373788 199344 373794
rect 199292 373730 199344 373736
rect 199396 367810 199424 391303
rect 199488 389881 199516 461654
rect 199580 461417 199608 461654
rect 199566 461408 199622 461417
rect 199566 461343 199622 461352
rect 199568 458856 199620 458862
rect 199568 458798 199620 458804
rect 199580 392737 199608 458798
rect 199750 394632 199806 394641
rect 199750 394567 199806 394576
rect 199566 392728 199622 392737
rect 199566 392663 199622 392672
rect 199474 389872 199530 389881
rect 199474 389807 199530 389816
rect 199488 389201 199516 389807
rect 199474 389192 199530 389201
rect 199474 389127 199530 389136
rect 199384 367804 199436 367810
rect 199384 367746 199436 367752
rect 199396 367690 199424 367746
rect 199396 367662 199516 367690
rect 199382 366344 199438 366353
rect 199382 366279 199438 366288
rect 198844 344986 199056 345014
rect 198844 344185 198872 344986
rect 198830 344176 198886 344185
rect 198830 344111 198886 344120
rect 198738 284336 198794 284345
rect 198738 284271 198794 284280
rect 198752 175001 198780 284271
rect 198844 234025 198872 344111
rect 199396 287054 199424 366279
rect 199028 287026 199424 287054
rect 198922 280120 198978 280129
rect 198922 280055 198978 280064
rect 198830 234016 198886 234025
rect 198830 233951 198886 233960
rect 198738 174992 198794 175001
rect 198738 174927 198794 174936
rect 198936 171134 198964 280055
rect 199028 278633 199056 287026
rect 199290 282704 199346 282713
rect 199290 282639 199346 282648
rect 199106 281344 199162 281353
rect 199106 281279 199162 281288
rect 199014 278624 199070 278633
rect 199014 278559 199070 278568
rect 198844 171106 198964 171134
rect 198844 169833 198872 171106
rect 198830 169824 198886 169833
rect 198830 169759 198886 169768
rect 198738 168464 198794 168473
rect 198738 168399 198794 168408
rect 198752 59265 198780 168399
rect 198844 60489 198872 169759
rect 199028 168473 199056 278559
rect 199120 171329 199148 281279
rect 199198 234016 199254 234025
rect 199198 233951 199254 233960
rect 199106 171320 199162 171329
rect 199106 171255 199162 171264
rect 199014 168464 199070 168473
rect 199014 168399 199070 168408
rect 199120 61985 199148 171255
rect 199212 124137 199240 233951
rect 199304 172689 199332 282639
rect 199488 281353 199516 367662
rect 199580 359514 199608 392663
rect 199658 389192 199714 389201
rect 199658 389127 199714 389136
rect 199568 359508 199620 359514
rect 199568 359450 199620 359456
rect 199672 356726 199700 389127
rect 199764 383654 199792 394567
rect 199764 383626 199884 383654
rect 199856 363662 199884 383626
rect 200224 369714 200252 489886
rect 200304 489524 200356 489530
rect 200304 489466 200356 489472
rect 200316 373930 200344 489466
rect 200396 489388 200448 489394
rect 200396 489330 200448 489336
rect 200304 373924 200356 373930
rect 200304 373866 200356 373872
rect 200408 373862 200436 489330
rect 200488 466064 200540 466070
rect 200488 466006 200540 466012
rect 200500 374338 200528 466006
rect 200580 461032 200632 461038
rect 200580 460974 200632 460980
rect 200592 374649 200620 460974
rect 200578 374640 200634 374649
rect 200578 374575 200634 374584
rect 200488 374332 200540 374338
rect 200488 374274 200540 374280
rect 200396 373856 200448 373862
rect 200396 373798 200448 373804
rect 200684 369782 200712 489886
rect 200856 467288 200908 467294
rect 200856 467230 200908 467236
rect 200764 463276 200816 463282
rect 200764 463218 200816 463224
rect 200672 369776 200724 369782
rect 200672 369718 200724 369724
rect 200212 369708 200264 369714
rect 200212 369650 200264 369656
rect 199844 363656 199896 363662
rect 199844 363598 199896 363604
rect 199752 359508 199804 359514
rect 199752 359450 199804 359456
rect 199660 356720 199712 356726
rect 199660 356662 199712 356668
rect 199474 281344 199530 281353
rect 199474 281279 199530 281288
rect 199672 280129 199700 356662
rect 199764 282713 199792 359450
rect 199856 284345 199884 363598
rect 199842 284336 199898 284345
rect 199842 284271 199898 284280
rect 199750 282704 199806 282713
rect 199750 282639 199806 282648
rect 199658 280120 199714 280129
rect 199658 280055 199714 280064
rect 200120 240984 200172 240990
rect 200120 240926 200172 240932
rect 199382 174992 199438 175001
rect 199382 174927 199438 174936
rect 199290 172680 199346 172689
rect 199290 172615 199346 172624
rect 199198 124128 199254 124137
rect 199198 124063 199254 124072
rect 199304 63345 199332 172615
rect 199396 64705 199424 174927
rect 200132 152522 200160 240926
rect 200776 152726 200804 463218
rect 200868 263158 200896 467230
rect 200948 465588 201000 465594
rect 200948 465530 201000 465536
rect 200960 264246 200988 465530
rect 201040 458788 201092 458794
rect 201040 458730 201092 458736
rect 201052 369238 201080 458730
rect 201512 374746 201540 495037
rect 201696 495023 201986 495051
rect 202064 495023 202446 495051
rect 201592 492516 201644 492522
rect 201592 492458 201644 492464
rect 201500 374740 201552 374746
rect 201500 374682 201552 374688
rect 201604 374066 201632 492458
rect 201696 374678 201724 495023
rect 202064 492522 202092 495023
rect 202052 492516 202104 492522
rect 202052 492458 202104 492464
rect 201776 492312 201828 492318
rect 201774 492280 201776 492289
rect 201828 492280 201830 492289
rect 201774 492215 201830 492224
rect 202144 492108 202196 492114
rect 202144 492050 202196 492056
rect 202788 492108 202840 492114
rect 202788 492050 202840 492056
rect 201776 465996 201828 466002
rect 201776 465938 201828 465944
rect 201684 374672 201736 374678
rect 201684 374614 201736 374620
rect 201788 374474 201816 465938
rect 201868 458924 201920 458930
rect 201868 458866 201920 458872
rect 201880 374814 201908 458866
rect 201868 374808 201920 374814
rect 201868 374750 201920 374756
rect 201776 374468 201828 374474
rect 201776 374410 201828 374416
rect 201592 374060 201644 374066
rect 201592 374002 201644 374008
rect 201592 371272 201644 371278
rect 201592 371214 201644 371220
rect 201040 369232 201092 369238
rect 201040 369174 201092 369180
rect 201500 351960 201552 351966
rect 201500 351902 201552 351908
rect 200948 264240 201000 264246
rect 200948 264182 201000 264188
rect 200856 263152 200908 263158
rect 200856 263094 200908 263100
rect 201512 242146 201540 351902
rect 201604 263022 201632 371214
rect 201592 263016 201644 263022
rect 201592 262958 201644 262964
rect 201500 242140 201552 242146
rect 201500 242082 201552 242088
rect 201500 240848 201552 240854
rect 201500 240790 201552 240796
rect 201512 153270 201540 240790
rect 202156 154222 202184 492050
rect 202420 491360 202472 491366
rect 202420 491302 202472 491308
rect 202236 467220 202288 467226
rect 202236 467162 202288 467168
rect 202248 262886 202276 467162
rect 202328 460896 202380 460902
rect 202328 460838 202380 460844
rect 202340 264489 202368 460838
rect 202432 370938 202460 491302
rect 202800 372298 202828 492050
rect 202788 372292 202840 372298
rect 202788 372234 202840 372240
rect 202800 372094 202828 372234
rect 202788 372088 202840 372094
rect 202788 372030 202840 372036
rect 202420 370932 202472 370938
rect 202420 370874 202472 370880
rect 202892 369850 202920 495037
rect 203076 495023 203274 495051
rect 203352 495023 203734 495051
rect 203904 495023 204194 495051
rect 204272 495023 204654 495051
rect 204732 495023 205022 495051
rect 205192 495023 205482 495051
rect 205652 495023 205942 495051
rect 202972 492516 203024 492522
rect 202972 492458 203024 492464
rect 202984 373994 203012 492458
rect 203076 374814 203104 495023
rect 203352 489914 203380 495023
rect 203904 492522 203932 495023
rect 203892 492516 203944 492522
rect 203892 492458 203944 492464
rect 204168 491428 204220 491434
rect 204168 491370 204220 491376
rect 203168 489886 203380 489914
rect 203168 462330 203196 489886
rect 203248 489320 203300 489326
rect 203248 489262 203300 489268
rect 203156 462324 203208 462330
rect 203156 462266 203208 462272
rect 203064 374808 203116 374814
rect 203064 374750 203116 374756
rect 202984 373966 203104 373994
rect 203076 373289 203104 373966
rect 203260 373522 203288 489262
rect 203616 476808 203668 476814
rect 203616 476750 203668 476756
rect 203340 465928 203392 465934
rect 203340 465870 203392 465876
rect 203248 373516 203300 373522
rect 203248 373458 203300 373464
rect 203062 373280 203118 373289
rect 203062 373215 203118 373224
rect 202972 371816 203024 371822
rect 202972 371758 203024 371764
rect 202880 369844 202932 369850
rect 202880 369786 202932 369792
rect 202880 351212 202932 351218
rect 202880 351154 202932 351160
rect 202892 274650 202920 351154
rect 202880 274644 202932 274650
rect 202880 274586 202932 274592
rect 202892 273970 202920 274586
rect 202880 273964 202932 273970
rect 202880 273906 202932 273912
rect 202326 264480 202382 264489
rect 202326 264415 202382 264424
rect 202984 262954 203012 371758
rect 203076 369578 203104 373215
rect 203352 373182 203380 465870
rect 203524 460012 203576 460018
rect 203524 459954 203576 459960
rect 203340 373176 203392 373182
rect 203340 373118 203392 373124
rect 203536 369646 203564 459954
rect 203524 369640 203576 369646
rect 203524 369582 203576 369588
rect 203064 369572 203116 369578
rect 203064 369514 203116 369520
rect 203064 351960 203116 351966
rect 203064 351902 203116 351908
rect 203076 351218 203104 351902
rect 203064 351212 203116 351218
rect 203064 351154 203116 351160
rect 202972 262948 203024 262954
rect 202972 262890 203024 262896
rect 202236 262880 202288 262886
rect 202236 262822 202288 262828
rect 203628 164218 203656 476750
rect 203708 462936 203760 462942
rect 203708 462878 203760 462884
rect 203720 264314 203748 462878
rect 203800 460148 203852 460154
rect 203800 460090 203852 460096
rect 203812 276010 203840 460090
rect 204180 372366 204208 491370
rect 204272 372774 204300 495023
rect 204732 492504 204760 495023
rect 204364 492476 204760 492504
rect 204364 489190 204392 492476
rect 205192 489914 205220 495023
rect 204456 489886 205220 489914
rect 204352 489184 204404 489190
rect 204352 489126 204404 489132
rect 204352 465792 204404 465798
rect 204352 465734 204404 465740
rect 204260 372768 204312 372774
rect 204260 372710 204312 372716
rect 204168 372360 204220 372366
rect 204168 372302 204220 372308
rect 204180 371958 204208 372302
rect 204168 371952 204220 371958
rect 204168 371894 204220 371900
rect 204168 371816 204220 371822
rect 204168 371758 204220 371764
rect 204180 371346 204208 371758
rect 204168 371340 204220 371346
rect 204168 371282 204220 371288
rect 204272 369442 204300 372710
rect 204260 369436 204312 369442
rect 204260 369378 204312 369384
rect 203800 276004 203852 276010
rect 203800 275946 203852 275952
rect 203708 264308 203760 264314
rect 203708 264250 203760 264256
rect 204364 263566 204392 465734
rect 204456 405006 204484 489886
rect 205652 482390 205680 495023
rect 206388 492386 206416 495037
rect 206480 495023 206862 495051
rect 205732 492380 205784 492386
rect 205732 492322 205784 492328
rect 206376 492380 206428 492386
rect 206376 492322 206428 492328
rect 205744 492153 205772 492322
rect 205730 492144 205786 492153
rect 205730 492079 205786 492088
rect 206480 489914 206508 495023
rect 207232 494834 207260 495037
rect 207308 495023 207690 495051
rect 207768 495023 208150 495051
rect 207220 494828 207272 494834
rect 207220 494770 207272 494776
rect 207112 493332 207164 493338
rect 207112 493274 207164 493280
rect 205744 489886 206508 489914
rect 205640 482384 205692 482390
rect 205640 482326 205692 482332
rect 205088 472728 205140 472734
rect 205088 472670 205140 472676
rect 204902 465896 204958 465905
rect 204536 465860 204588 465866
rect 204902 465831 204958 465840
rect 204536 465802 204588 465808
rect 204444 405000 204496 405006
rect 204444 404942 204496 404948
rect 204548 374202 204576 465802
rect 204536 374196 204588 374202
rect 204536 374138 204588 374144
rect 204352 263560 204404 263566
rect 204352 263502 204404 263508
rect 203616 164212 203668 164218
rect 203616 164154 203668 164160
rect 202144 154216 202196 154222
rect 202144 154158 202196 154164
rect 201500 153264 201552 153270
rect 201500 153206 201552 153212
rect 200764 152720 200816 152726
rect 200764 152662 200816 152668
rect 204916 152590 204944 465831
rect 204996 460420 205048 460426
rect 204996 460362 205048 460368
rect 205008 154154 205036 460362
rect 205100 263430 205128 472670
rect 205640 465724 205692 465730
rect 205640 465666 205692 465672
rect 205364 465520 205416 465526
rect 205364 465462 205416 465468
rect 205180 462868 205232 462874
rect 205180 462810 205232 462816
rect 205088 263424 205140 263430
rect 205088 263366 205140 263372
rect 205192 262138 205220 462810
rect 205272 462188 205324 462194
rect 205272 462130 205324 462136
rect 205284 262721 205312 462130
rect 205376 369510 205404 465462
rect 205364 369504 205416 369510
rect 205364 369446 205416 369452
rect 205652 263498 205680 465666
rect 205744 409154 205772 489886
rect 205824 489252 205876 489258
rect 205824 489194 205876 489200
rect 205732 409148 205784 409154
rect 205732 409090 205784 409096
rect 205836 373658 205864 489194
rect 206560 471368 206612 471374
rect 206560 471310 206612 471316
rect 206284 462324 206336 462330
rect 206284 462266 206336 462272
rect 206296 385014 206324 462266
rect 206376 460352 206428 460358
rect 206376 460294 206428 460300
rect 206284 385008 206336 385014
rect 206284 384950 206336 384956
rect 206284 382288 206336 382294
rect 206284 382230 206336 382236
rect 205824 373652 205876 373658
rect 205824 373594 205876 373600
rect 206296 351966 206324 382230
rect 206284 351960 206336 351966
rect 206284 351902 206336 351908
rect 205640 263492 205692 263498
rect 205640 263434 205692 263440
rect 205270 262712 205326 262721
rect 205270 262647 205326 262656
rect 205180 262132 205232 262138
rect 205180 262074 205232 262080
rect 204996 154148 205048 154154
rect 204996 154090 205048 154096
rect 206388 154018 206416 460294
rect 206466 459096 206522 459105
rect 206466 459031 206522 459040
rect 206480 154290 206508 459031
rect 206572 263090 206600 471310
rect 206652 465656 206704 465662
rect 206652 465598 206704 465604
rect 206560 263084 206612 263090
rect 206560 263026 206612 263032
rect 206664 262206 206692 465598
rect 206836 462800 206888 462806
rect 206836 462742 206888 462748
rect 206744 459264 206796 459270
rect 206744 459206 206796 459212
rect 206756 273222 206784 459206
rect 206848 370462 206876 462742
rect 207020 462392 207072 462398
rect 207020 462334 207072 462340
rect 207032 461650 207060 462334
rect 207020 461644 207072 461650
rect 207020 461586 207072 461592
rect 207020 460964 207072 460970
rect 207020 460906 207072 460912
rect 207032 383654 207060 460906
rect 207020 383648 207072 383654
rect 207020 383590 207072 383596
rect 207032 382294 207060 383590
rect 207020 382288 207072 382294
rect 207020 382230 207072 382236
rect 206836 370456 206888 370462
rect 206836 370398 206888 370404
rect 206744 273216 206796 273222
rect 206744 273158 206796 273164
rect 207124 263362 207152 493274
rect 207204 491700 207256 491706
rect 207204 491642 207256 491648
rect 207216 372706 207244 491642
rect 207308 462398 207336 495023
rect 207388 494828 207440 494834
rect 207388 494770 207440 494776
rect 207296 462392 207348 462398
rect 207296 462334 207348 462340
rect 207400 458250 207428 494770
rect 207768 491706 207796 495023
rect 208492 492516 208544 492522
rect 208492 492458 208544 492464
rect 208400 492448 208452 492454
rect 208400 492390 208452 492396
rect 207756 491700 207808 491706
rect 207756 491642 207808 491648
rect 207848 466268 207900 466274
rect 207848 466210 207900 466216
rect 207662 466032 207718 466041
rect 207662 465967 207718 465976
rect 207480 463072 207532 463078
rect 207480 463014 207532 463020
rect 207388 458244 207440 458250
rect 207388 458186 207440 458192
rect 207492 374406 207520 463014
rect 207480 374400 207532 374406
rect 207480 374342 207532 374348
rect 207204 372700 207256 372706
rect 207204 372642 207256 372648
rect 207216 369102 207244 372642
rect 207204 369096 207256 369102
rect 207204 369038 207256 369044
rect 207112 263356 207164 263362
rect 207112 263298 207164 263304
rect 206652 262200 206704 262206
rect 206652 262142 206704 262148
rect 206468 154284 206520 154290
rect 206468 154226 206520 154232
rect 206376 154012 206428 154018
rect 206376 153954 206428 153960
rect 207676 152833 207704 465967
rect 207756 460692 207808 460698
rect 207756 460634 207808 460640
rect 207768 165578 207796 460634
rect 207860 264722 207888 466210
rect 207940 463412 207992 463418
rect 207940 463354 207992 463360
rect 207848 264716 207900 264722
rect 207848 264658 207900 264664
rect 207952 262818 207980 463354
rect 208032 459536 208084 459542
rect 208032 459478 208084 459484
rect 208044 370326 208072 459478
rect 208124 458244 208176 458250
rect 208124 458186 208176 458192
rect 208136 410582 208164 458186
rect 208124 410576 208176 410582
rect 208124 410518 208176 410524
rect 208122 373416 208178 373425
rect 208122 373351 208178 373360
rect 208032 370320 208084 370326
rect 208032 370262 208084 370268
rect 208136 369374 208164 373351
rect 208412 372502 208440 492390
rect 208504 372570 208532 492458
rect 208492 372564 208544 372570
rect 208492 372506 208544 372512
rect 208400 372496 208452 372502
rect 208400 372438 208452 372444
rect 208596 370258 208624 495037
rect 208688 495023 209070 495051
rect 209148 495023 209438 495051
rect 209792 495023 209898 495051
rect 209976 495023 210358 495051
rect 210528 495023 210818 495051
rect 211202 495023 211384 495051
rect 208688 492522 208716 495023
rect 208676 492516 208728 492522
rect 208676 492458 208728 492464
rect 209148 492454 209176 495023
rect 209136 492448 209188 492454
rect 209136 492390 209188 492396
rect 209228 492380 209280 492386
rect 209228 492322 209280 492328
rect 209044 485104 209096 485110
rect 209044 485046 209096 485052
rect 208860 460080 208912 460086
rect 208860 460022 208912 460028
rect 208584 370252 208636 370258
rect 208584 370194 208636 370200
rect 208872 369374 208900 460022
rect 208952 374876 209004 374882
rect 208952 374818 209004 374824
rect 208124 369368 208176 369374
rect 208124 369310 208176 369316
rect 208860 369368 208912 369374
rect 208860 369310 208912 369316
rect 208136 354674 208164 369310
rect 208964 369306 208992 374818
rect 208952 369300 209004 369306
rect 208952 369242 209004 369248
rect 208044 354646 208164 354674
rect 208044 264790 208072 354646
rect 208032 264784 208084 264790
rect 208032 264726 208084 264732
rect 207940 262812 207992 262818
rect 207940 262754 207992 262760
rect 208964 261526 208992 369242
rect 208952 261520 209004 261526
rect 208952 261462 209004 261468
rect 207756 165572 207808 165578
rect 207756 165514 207808 165520
rect 209056 153134 209084 485046
rect 209240 467158 209268 492322
rect 209136 467152 209188 467158
rect 209136 467094 209188 467100
rect 209228 467152 209280 467158
rect 209228 467094 209280 467100
rect 209044 153128 209096 153134
rect 209044 153070 209096 153076
rect 207662 152824 207718 152833
rect 209148 152794 209176 467094
rect 209320 466336 209372 466342
rect 209320 466278 209372 466284
rect 209226 463312 209282 463321
rect 209226 463247 209282 463256
rect 209240 153882 209268 463247
rect 209332 263226 209360 466278
rect 209412 461984 209464 461990
rect 209412 461926 209464 461932
rect 209424 264382 209452 461926
rect 209504 459400 209556 459406
rect 209504 459342 209556 459348
rect 209516 383586 209544 459342
rect 209504 383580 209556 383586
rect 209504 383522 209556 383528
rect 209792 373522 209820 495023
rect 209872 492516 209924 492522
rect 209872 492458 209924 492464
rect 209780 373516 209832 373522
rect 209780 373458 209832 373464
rect 209686 372600 209742 372609
rect 209686 372535 209742 372544
rect 209502 372056 209558 372065
rect 209502 371991 209558 372000
rect 209412 264376 209464 264382
rect 209412 264318 209464 264324
rect 209320 263220 209372 263226
rect 209320 263162 209372 263168
rect 209516 240786 209544 371991
rect 209594 371240 209650 371249
rect 209594 371175 209650 371184
rect 209504 240780 209556 240786
rect 209504 240722 209556 240728
rect 209228 153876 209280 153882
rect 209228 153818 209280 153824
rect 207662 152759 207718 152768
rect 209136 152788 209188 152794
rect 209136 152730 209188 152736
rect 204904 152584 204956 152590
rect 204904 152526 204956 152532
rect 200120 152516 200172 152522
rect 200120 152458 200172 152464
rect 199382 64696 199438 64705
rect 199382 64631 199438 64640
rect 199290 63336 199346 63345
rect 199290 63271 199346 63280
rect 199106 61976 199162 61985
rect 199106 61911 199162 61920
rect 198830 60480 198886 60489
rect 198830 60415 198886 60424
rect 198738 59256 198794 59265
rect 198738 59191 198794 59200
rect 198648 43512 198700 43518
rect 198648 43454 198700 43460
rect 209608 42770 209636 371175
rect 197452 42764 197504 42770
rect 197452 42706 197504 42712
rect 209596 42764 209648 42770
rect 209596 42706 209648 42712
rect 135904 42696 135956 42702
rect 183192 42696 183244 42702
rect 135904 42638 135956 42644
rect 183190 42664 183192 42673
rect 197360 42696 197412 42702
rect 183244 42664 183246 42673
rect 133420 42628 133472 42634
rect 197360 42638 197412 42644
rect 183190 42599 183246 42608
rect 133420 42570 133472 42576
rect 128360 42560 128412 42566
rect 128360 42502 128412 42508
rect 165802 42528 165858 42537
rect 165802 42463 165858 42472
rect 119068 41336 119120 41342
rect 119068 41278 119120 41284
rect 116308 40044 116360 40050
rect 116308 39986 116360 39992
rect 111892 39976 111944 39982
rect 165816 39953 165844 42463
rect 209700 42362 209728 372535
rect 209884 371618 209912 492458
rect 209872 371612 209924 371618
rect 209872 371554 209924 371560
rect 209976 371550 210004 495023
rect 210528 492522 210556 495023
rect 211160 492584 211212 492590
rect 211160 492526 211212 492532
rect 210516 492516 210568 492522
rect 210516 492458 210568 492464
rect 211172 491609 211200 492526
rect 211158 491600 211214 491609
rect 211158 491535 211214 491544
rect 210424 482316 210476 482322
rect 210424 482258 210476 482264
rect 210056 462256 210108 462262
rect 210056 462198 210108 462204
rect 209964 371544 210016 371550
rect 209964 371486 210016 371492
rect 210068 263294 210096 462198
rect 210240 460760 210292 460766
rect 210240 460702 210292 460708
rect 210252 369034 210280 460702
rect 210332 372496 210384 372502
rect 210332 372438 210384 372444
rect 210344 372026 210372 372438
rect 210332 372020 210384 372026
rect 210332 371962 210384 371968
rect 210240 369028 210292 369034
rect 210240 368970 210292 368976
rect 210056 263288 210108 263294
rect 210056 263230 210108 263236
rect 210344 262682 210372 371962
rect 210332 262676 210384 262682
rect 210332 262618 210384 262624
rect 210436 153202 210464 482258
rect 210608 479596 210660 479602
rect 210608 479538 210660 479544
rect 210516 463208 210568 463214
rect 210516 463150 210568 463156
rect 210528 153950 210556 463150
rect 210620 263294 210648 479538
rect 210700 472796 210752 472802
rect 210700 472738 210752 472744
rect 210712 263566 210740 472738
rect 210792 459332 210844 459338
rect 210792 459274 210844 459280
rect 210804 264450 210832 459274
rect 211068 373516 211120 373522
rect 211068 373458 211120 373464
rect 210976 372564 211028 372570
rect 210976 372506 211028 372512
rect 210988 372298 211016 372506
rect 210976 372292 211028 372298
rect 210976 372234 211028 372240
rect 210884 371408 210936 371414
rect 210884 371350 210936 371356
rect 210792 264444 210844 264450
rect 210792 264386 210844 264392
rect 210700 263560 210752 263566
rect 210700 263502 210752 263508
rect 210608 263288 210660 263294
rect 210608 263230 210660 263236
rect 210896 240990 210924 371350
rect 210988 241466 211016 372234
rect 211080 371686 211108 373458
rect 211356 372230 211384 495023
rect 211632 491434 211660 495037
rect 212092 492114 212120 495037
rect 212080 492108 212132 492114
rect 212080 492050 212132 492056
rect 212448 491972 212500 491978
rect 212448 491914 212500 491920
rect 211620 491428 211672 491434
rect 211620 491370 211672 491376
rect 211804 481024 211856 481030
rect 211804 480966 211856 480972
rect 211436 461916 211488 461922
rect 211436 461858 211488 461864
rect 211344 372224 211396 372230
rect 211344 372166 211396 372172
rect 211068 371680 211120 371686
rect 211068 371622 211120 371628
rect 211066 369200 211122 369209
rect 211066 369135 211122 369144
rect 210976 241460 211028 241466
rect 210976 241402 211028 241408
rect 210884 240984 210936 240990
rect 210884 240926 210936 240932
rect 210792 240780 210844 240786
rect 210792 240722 210844 240728
rect 210516 153944 210568 153950
rect 210516 153886 210568 153892
rect 210424 153196 210476 153202
rect 210424 153138 210476 153144
rect 210804 133686 210832 240722
rect 210792 133680 210844 133686
rect 210792 133622 210844 133628
rect 210896 130529 210924 240926
rect 210882 130520 210938 130529
rect 210882 130455 210938 130464
rect 211080 42566 211108 369135
rect 211448 264353 211476 461858
rect 211528 459468 211580 459474
rect 211528 459410 211580 459416
rect 211540 369578 211568 459410
rect 211618 372192 211674 372201
rect 211618 372127 211674 372136
rect 211528 369572 211580 369578
rect 211528 369514 211580 369520
rect 211434 264344 211490 264353
rect 211434 264279 211490 264288
rect 211632 263702 211660 372127
rect 211710 370560 211766 370569
rect 211710 370495 211766 370504
rect 211620 263696 211672 263702
rect 211620 263638 211672 263644
rect 211724 262070 211752 370495
rect 211712 262064 211764 262070
rect 211712 262006 211764 262012
rect 211068 42560 211120 42566
rect 211068 42502 211120 42508
rect 209688 42356 209740 42362
rect 209688 42298 209740 42304
rect 211816 42226 211844 480966
rect 211896 478168 211948 478174
rect 211896 478110 211948 478116
rect 211804 42220 211856 42226
rect 211804 42162 211856 42168
rect 211908 42090 211936 478110
rect 211988 471300 212040 471306
rect 211988 471242 212040 471248
rect 212000 152998 212028 471242
rect 212172 469940 212224 469946
rect 212172 469882 212224 469888
rect 212080 461848 212132 461854
rect 212080 461790 212132 461796
rect 211988 152992 212040 152998
rect 211988 152934 212040 152940
rect 212092 151774 212120 461790
rect 212184 262954 212212 469882
rect 212264 463480 212316 463486
rect 212264 463422 212316 463428
rect 212276 263498 212304 463422
rect 212460 370394 212488 491914
rect 212552 373318 212580 495037
rect 212644 495023 213026 495051
rect 213104 495023 213394 495051
rect 213472 495023 213854 495051
rect 213932 495023 214314 495051
rect 214392 495023 214774 495051
rect 214852 495023 215234 495051
rect 215404 495023 215602 495051
rect 215680 495023 216062 495051
rect 216232 495023 216522 495051
rect 216998 495023 217272 495051
rect 212644 373386 212672 495023
rect 212816 492652 212868 492658
rect 212816 492594 212868 492600
rect 212828 492561 212856 492594
rect 212814 492552 212870 492561
rect 212724 492516 212776 492522
rect 212814 492487 212870 492496
rect 212724 492458 212776 492464
rect 212736 373454 212764 492458
rect 213104 489914 213132 495023
rect 213472 492522 213500 495023
rect 213460 492516 213512 492522
rect 213460 492458 213512 492464
rect 212828 489886 213132 489914
rect 212828 380610 212856 489886
rect 213184 474020 213236 474026
rect 213184 473962 213236 473968
rect 212908 466404 212960 466410
rect 212908 466346 212960 466352
rect 212920 380730 212948 466346
rect 213000 460828 213052 460834
rect 213000 460770 213052 460776
rect 213012 383654 213040 460770
rect 213012 383626 213132 383654
rect 212908 380724 212960 380730
rect 212908 380666 212960 380672
rect 212828 380582 213040 380610
rect 212908 380520 212960 380526
rect 212908 380462 212960 380468
rect 212814 373688 212870 373697
rect 212814 373623 212870 373632
rect 212724 373448 212776 373454
rect 212724 373390 212776 373396
rect 212632 373380 212684 373386
rect 212632 373322 212684 373328
rect 212540 373312 212592 373318
rect 212540 373254 212592 373260
rect 212644 373182 212672 373322
rect 212632 373176 212684 373182
rect 212632 373118 212684 373124
rect 212736 373114 212764 373390
rect 212724 373108 212776 373114
rect 212724 373050 212776 373056
rect 212828 373046 212856 373623
rect 212816 373040 212868 373046
rect 212816 372982 212868 372988
rect 212724 372564 212776 372570
rect 212724 372506 212776 372512
rect 212736 371754 212764 372506
rect 212724 371748 212776 371754
rect 212724 371690 212776 371696
rect 212448 370388 212500 370394
rect 212448 370330 212500 370336
rect 212446 369200 212502 369209
rect 212446 369135 212502 369144
rect 212356 263628 212408 263634
rect 212356 263570 212408 263576
rect 212264 263492 212316 263498
rect 212264 263434 212316 263440
rect 212172 262948 212224 262954
rect 212172 262890 212224 262896
rect 212264 151836 212316 151842
rect 212264 151778 212316 151784
rect 212080 151768 212132 151774
rect 212080 151710 212132 151716
rect 211896 42084 211948 42090
rect 211896 42026 211948 42032
rect 212276 41138 212304 151778
rect 212368 133890 212396 263570
rect 212356 133884 212408 133890
rect 212356 133826 212408 133832
rect 212264 41132 212316 41138
rect 212264 41074 212316 41080
rect 111892 39918 111944 39924
rect 165802 39944 165858 39953
rect 111156 39908 111208 39914
rect 165802 39879 165858 39888
rect 111156 39850 111208 39856
rect 109316 39840 109368 39846
rect 109316 39782 109368 39788
rect 93308 39636 93360 39642
rect 93308 39578 93360 39584
rect 89996 39500 90048 39506
rect 89996 39442 90048 39448
rect 81808 39432 81860 39438
rect 81808 39374 81860 39380
rect 78772 39364 78824 39370
rect 78772 39306 78824 39312
rect 212368 39302 212396 133826
rect 212460 43722 212488 369135
rect 212736 364334 212764 371690
rect 212920 369442 212948 380462
rect 213012 373697 213040 380582
rect 213104 374134 213132 383626
rect 213092 374128 213144 374134
rect 213092 374070 213144 374076
rect 212998 373688 213054 373697
rect 212998 373623 213054 373632
rect 213090 373280 213146 373289
rect 213090 373215 213146 373224
rect 212908 369436 212960 369442
rect 212908 369378 212960 369384
rect 212736 364306 213040 364334
rect 213012 264178 213040 364306
rect 213000 264172 213052 264178
rect 213000 264114 213052 264120
rect 213012 263634 213040 264114
rect 213000 263628 213052 263634
rect 213000 263570 213052 263576
rect 212908 262064 212960 262070
rect 212908 262006 212960 262012
rect 212920 261594 212948 262006
rect 212908 261588 212960 261594
rect 212908 261530 212960 261536
rect 212816 261520 212868 261526
rect 212816 261462 212868 261468
rect 212828 149734 212856 261462
rect 212816 149728 212868 149734
rect 212816 149670 212868 149676
rect 212920 129674 212948 261530
rect 213104 260778 213132 373215
rect 213092 260772 213144 260778
rect 213092 260714 213144 260720
rect 213000 241324 213052 241330
rect 213000 241266 213052 241272
rect 213012 130558 213040 241266
rect 213196 152522 213224 473962
rect 213276 463548 213328 463554
rect 213276 463490 213328 463496
rect 213288 263265 213316 463490
rect 213458 459504 213514 459513
rect 213458 459439 213514 459448
rect 213368 372428 213420 372434
rect 213368 372370 213420 372376
rect 213380 371754 213408 372370
rect 213368 371748 213420 371754
rect 213368 371690 213420 371696
rect 213274 263256 213330 263265
rect 213274 263191 213330 263200
rect 213276 262676 213328 262682
rect 213276 262618 213328 262624
rect 213288 262274 213316 262618
rect 213276 262268 213328 262274
rect 213276 262210 213328 262216
rect 213184 152516 213236 152522
rect 213184 152458 213236 152464
rect 213288 151094 213316 262210
rect 213380 240922 213408 371690
rect 213472 263401 213500 459439
rect 213552 374468 213604 374474
rect 213552 374410 213604 374416
rect 213564 370258 213592 374410
rect 213826 373824 213882 373833
rect 213826 373759 213882 373768
rect 213644 373040 213696 373046
rect 213644 372982 213696 372988
rect 213552 370252 213604 370258
rect 213552 370194 213604 370200
rect 213458 263392 213514 263401
rect 213458 263327 213514 263336
rect 213564 260846 213592 370194
rect 213552 260840 213604 260846
rect 213552 260782 213604 260788
rect 213564 258074 213592 260782
rect 213472 258046 213592 258074
rect 213368 240916 213420 240922
rect 213368 240858 213420 240864
rect 213276 151088 213328 151094
rect 213276 151030 213328 151036
rect 213368 133884 213420 133890
rect 213368 133826 213420 133832
rect 213000 130552 213052 130558
rect 213000 130494 213052 130500
rect 212908 129668 212960 129674
rect 212908 129610 212960 129616
rect 212448 43716 212500 43722
rect 212448 43658 212500 43664
rect 213380 40730 213408 133826
rect 213472 129742 213500 258046
rect 213552 240576 213604 240582
rect 213552 240518 213604 240524
rect 213564 133890 213592 240518
rect 213656 240038 213684 372982
rect 213734 369200 213790 369209
rect 213734 369135 213790 369144
rect 213644 240032 213696 240038
rect 213644 239974 213696 239980
rect 213552 133884 213604 133890
rect 213552 133826 213604 133832
rect 213644 133476 213696 133482
rect 213644 133418 213696 133424
rect 213552 131164 213604 131170
rect 213552 131106 213604 131112
rect 213460 129736 213512 129742
rect 213460 129678 213512 129684
rect 213368 40724 213420 40730
rect 213368 40666 213420 40672
rect 213564 39370 213592 131106
rect 213656 40050 213684 133418
rect 213748 43654 213776 369135
rect 213736 43648 213788 43654
rect 213736 43590 213788 43596
rect 213840 42498 213868 373759
rect 213932 372842 213960 495023
rect 214392 492538 214420 495023
rect 214024 492510 214420 492538
rect 214024 372978 214052 492510
rect 214852 489914 214880 495023
rect 215300 492516 215352 492522
rect 215300 492458 215352 492464
rect 214116 489886 214880 489914
rect 214012 372972 214064 372978
rect 214012 372914 214064 372920
rect 213920 372836 213972 372842
rect 213920 372778 213972 372784
rect 213918 372464 213974 372473
rect 213918 372399 213974 372408
rect 213932 371793 213960 372399
rect 213918 371784 213974 371793
rect 213918 371719 213974 371728
rect 214024 368966 214052 372914
rect 214116 372638 214144 489886
rect 214656 468580 214708 468586
rect 214656 468522 214708 468528
rect 214564 464364 214616 464370
rect 214564 464306 214616 464312
rect 214380 463684 214432 463690
rect 214380 463626 214432 463632
rect 214288 459672 214340 459678
rect 214288 459614 214340 459620
rect 214104 372632 214156 372638
rect 214104 372574 214156 372580
rect 214116 369170 214144 372574
rect 214300 372473 214328 459614
rect 214286 372464 214342 372473
rect 214286 372399 214342 372408
rect 214104 369164 214156 369170
rect 214104 369106 214156 369112
rect 214392 369102 214420 463626
rect 214472 369164 214524 369170
rect 214472 369106 214524 369112
rect 214380 369096 214432 369102
rect 214380 369038 214432 369044
rect 214012 368960 214064 368966
rect 214012 368902 214064 368908
rect 214380 265396 214432 265402
rect 214380 265338 214432 265344
rect 214288 263696 214340 263702
rect 214288 263638 214340 263644
rect 214300 258074 214328 263638
rect 214392 260846 214420 265338
rect 214380 260840 214432 260846
rect 214380 260782 214432 260788
rect 214300 258046 214420 258074
rect 214288 241460 214340 241466
rect 214288 241402 214340 241408
rect 214300 240854 214328 241402
rect 214288 240848 214340 240854
rect 214288 240790 214340 240796
rect 214196 150476 214248 150482
rect 214196 150418 214248 150424
rect 214208 43790 214236 150418
rect 214300 130490 214328 240790
rect 214392 131073 214420 258046
rect 214484 238746 214512 369106
rect 214472 238740 214524 238746
rect 214472 238682 214524 238688
rect 214576 152454 214604 464306
rect 214668 265266 214696 468522
rect 214748 460624 214800 460630
rect 214748 460566 214800 460572
rect 214656 265260 214708 265266
rect 214656 265202 214708 265208
rect 214656 264784 214708 264790
rect 214656 264726 214708 264732
rect 214668 264110 214696 264726
rect 214656 264104 214708 264110
rect 214656 264046 214708 264052
rect 214760 263362 214788 460566
rect 214840 460556 214892 460562
rect 214840 460498 214892 460504
rect 214852 264586 214880 460498
rect 215312 373726 215340 492458
rect 215300 373720 215352 373726
rect 215300 373662 215352 373668
rect 215300 373584 215352 373590
rect 215300 373526 215352 373532
rect 214932 373516 214984 373522
rect 214932 373458 214984 373464
rect 214840 264580 214892 264586
rect 214840 264522 214892 264528
rect 214748 263356 214800 263362
rect 214748 263298 214800 263304
rect 214840 260840 214892 260846
rect 214840 260782 214892 260788
rect 214748 260772 214800 260778
rect 214748 260714 214800 260720
rect 214760 260166 214788 260714
rect 214748 260160 214800 260166
rect 214748 260102 214800 260108
rect 214656 241460 214708 241466
rect 214656 241402 214708 241408
rect 214564 152448 214616 152454
rect 214564 152390 214616 152396
rect 214668 133822 214696 241402
rect 214760 150414 214788 260102
rect 214748 150408 214800 150414
rect 214748 150350 214800 150356
rect 214656 133816 214708 133822
rect 214656 133758 214708 133764
rect 214668 133482 214696 133758
rect 214656 133476 214708 133482
rect 214656 133418 214708 133424
rect 214852 132494 214880 260782
rect 214944 241330 214972 373458
rect 215024 373448 215076 373454
rect 215024 373390 215076 373396
rect 215036 372706 215064 373390
rect 215208 372836 215260 372842
rect 215208 372778 215260 372784
rect 215024 372700 215076 372706
rect 215024 372642 215076 372648
rect 215036 265402 215064 372642
rect 215114 369200 215170 369209
rect 215114 369135 215170 369144
rect 215024 265396 215076 265402
rect 215024 265338 215076 265344
rect 215024 265260 215076 265266
rect 215024 265202 215076 265208
rect 215036 262750 215064 265202
rect 215024 262744 215076 262750
rect 215024 262686 215076 262692
rect 214932 241324 214984 241330
rect 214932 241266 214984 241272
rect 214932 240100 214984 240106
rect 214932 240042 214984 240048
rect 214944 151434 214972 240042
rect 214932 151428 214984 151434
rect 214932 151370 214984 151376
rect 214944 150482 214972 151370
rect 214932 150476 214984 150482
rect 214932 150418 214984 150424
rect 214932 149728 214984 149734
rect 214932 149670 214984 149676
rect 214484 132466 214880 132494
rect 214378 131064 214434 131073
rect 214378 130999 214434 131008
rect 214288 130484 214340 130490
rect 214288 130426 214340 130432
rect 214196 43784 214248 43790
rect 214196 43726 214248 43732
rect 213828 42492 213880 42498
rect 213828 42434 213880 42440
rect 214392 41274 214420 130999
rect 214484 130626 214512 132466
rect 214656 130688 214708 130694
rect 214656 130630 214708 130636
rect 214472 130620 214524 130626
rect 214472 130562 214524 130568
rect 214484 44470 214512 130562
rect 214668 130490 214696 130630
rect 214838 130520 214894 130529
rect 214656 130484 214708 130490
rect 214838 130455 214894 130464
rect 214656 130426 214708 130432
rect 214564 130416 214616 130422
rect 214564 130358 214616 130364
rect 214576 53174 214604 130358
rect 214564 53168 214616 53174
rect 214564 53110 214616 53116
rect 214472 44464 214524 44470
rect 214472 44406 214524 44412
rect 214380 41268 214432 41274
rect 214380 41210 214432 41216
rect 214668 40798 214696 130426
rect 214656 40792 214708 40798
rect 214656 40734 214708 40740
rect 213644 40044 213696 40050
rect 213644 39986 213696 39992
rect 214852 39982 214880 130455
rect 214944 41206 214972 149670
rect 215024 133680 215076 133686
rect 215024 133622 215076 133628
rect 215036 133278 215064 133622
rect 215024 133272 215076 133278
rect 215024 133214 215076 133220
rect 214932 41200 214984 41206
rect 214932 41142 214984 41148
rect 215036 40662 215064 133214
rect 215128 42430 215156 369135
rect 215220 238678 215248 372778
rect 215312 372774 215340 373526
rect 215300 372768 215352 372774
rect 215300 372710 215352 372716
rect 215404 372706 215432 495023
rect 215680 489914 215708 495023
rect 216232 492522 216260 495023
rect 216220 492516 216272 492522
rect 216220 492458 216272 492464
rect 217244 492425 217272 495023
rect 217336 495023 217442 495051
rect 217230 492416 217286 492425
rect 217230 492351 217286 492360
rect 217336 489914 217364 495023
rect 217796 492561 217824 495037
rect 218164 495023 218270 495051
rect 218348 495023 218730 495051
rect 218808 495023 219190 495051
rect 217782 492552 217838 492561
rect 217782 492487 217838 492496
rect 218060 492516 218112 492522
rect 218060 492458 218112 492464
rect 217416 492040 217468 492046
rect 217416 491982 217468 491988
rect 215496 489886 215708 489914
rect 216692 489886 217364 489914
rect 215496 374270 215524 489886
rect 215944 483676 215996 483682
rect 215944 483618 215996 483624
rect 215852 462120 215904 462126
rect 215852 462062 215904 462068
rect 215484 374264 215536 374270
rect 215484 374206 215536 374212
rect 215392 372700 215444 372706
rect 215392 372642 215444 372648
rect 215300 372156 215352 372162
rect 215300 372098 215352 372104
rect 215312 371822 215340 372098
rect 215300 371816 215352 371822
rect 215300 371758 215352 371764
rect 215496 371074 215524 374206
rect 215576 373720 215628 373726
rect 215576 373662 215628 373668
rect 215484 371068 215536 371074
rect 215484 371010 215536 371016
rect 215496 369918 215524 371010
rect 215484 369912 215536 369918
rect 215484 369854 215536 369860
rect 215300 368960 215352 368966
rect 215300 368902 215352 368908
rect 215312 240106 215340 368902
rect 215588 368830 215616 373662
rect 215864 369170 215892 462062
rect 215852 369164 215904 369170
rect 215852 369106 215904 369112
rect 215576 368824 215628 368830
rect 215576 368766 215628 368772
rect 215758 262984 215814 262993
rect 215758 262919 215814 262928
rect 215300 240100 215352 240106
rect 215300 240042 215352 240048
rect 215312 239766 215340 240042
rect 215668 240032 215720 240038
rect 215668 239974 215720 239980
rect 215300 239760 215352 239766
rect 215300 239702 215352 239708
rect 215680 239562 215708 239974
rect 215668 239556 215720 239562
rect 215668 239498 215720 239504
rect 215208 238672 215260 238678
rect 215208 238614 215260 238620
rect 215680 130422 215708 239498
rect 215668 130416 215720 130422
rect 215668 130358 215720 130364
rect 215772 130354 215800 262919
rect 215956 153066 215984 483618
rect 216036 479528 216088 479534
rect 216036 479470 216088 479476
rect 215944 153060 215996 153066
rect 215944 153002 215996 153008
rect 216048 152658 216076 479470
rect 216128 464432 216180 464438
rect 216128 464374 216180 464380
rect 216140 152930 216168 464374
rect 216220 463344 216272 463350
rect 216220 463286 216272 463292
rect 216232 264518 216260 463286
rect 216312 459604 216364 459610
rect 216312 459546 216364 459552
rect 216324 372337 216352 459546
rect 216692 385098 216720 489886
rect 217324 489184 217376 489190
rect 217324 489126 217376 489132
rect 216770 410952 216826 410961
rect 216770 410887 216826 410896
rect 216784 410582 216812 410887
rect 216772 410576 216824 410582
rect 216772 410518 216824 410524
rect 216772 409148 216824 409154
rect 216772 409090 216824 409096
rect 216784 408785 216812 409090
rect 216770 408776 216826 408785
rect 216770 408711 216826 408720
rect 216600 385070 216720 385098
rect 216600 384826 216628 385070
rect 216680 385008 216732 385014
rect 216678 384976 216680 384985
rect 216732 384976 216734 384985
rect 216678 384911 216734 384920
rect 216600 384798 216720 384826
rect 216692 383738 216720 384798
rect 216600 383710 216720 383738
rect 216600 383194 216628 383710
rect 216680 383648 216732 383654
rect 216680 383590 216732 383596
rect 216692 383353 216720 383590
rect 216678 383344 216734 383353
rect 216678 383279 216734 383288
rect 216600 383166 216720 383194
rect 216496 373584 216548 373590
rect 216496 373526 216548 373532
rect 216404 372700 216456 372706
rect 216404 372642 216456 372648
rect 216310 372328 216366 372337
rect 216310 372263 216366 372272
rect 216312 371816 216364 371822
rect 216312 371758 216364 371764
rect 216220 264512 216272 264518
rect 216220 264454 216272 264460
rect 216324 240582 216352 371758
rect 216416 368898 216444 372642
rect 216404 368892 216456 368898
rect 216404 368834 216456 368840
rect 216312 240576 216364 240582
rect 216312 240518 216364 240524
rect 216312 240440 216364 240446
rect 216312 240382 216364 240388
rect 216220 239420 216272 239426
rect 216220 239362 216272 239368
rect 216232 238746 216260 239362
rect 216220 238740 216272 238746
rect 216220 238682 216272 238688
rect 216128 152924 216180 152930
rect 216128 152866 216180 152872
rect 216036 152652 216088 152658
rect 216036 152594 216088 152600
rect 216232 151366 216260 238682
rect 216220 151360 216272 151366
rect 216220 151302 216272 151308
rect 216128 150476 216180 150482
rect 216128 150418 216180 150424
rect 216036 131096 216088 131102
rect 216036 131038 216088 131044
rect 215944 130484 215996 130490
rect 215944 130426 215996 130432
rect 215850 130384 215906 130393
rect 215760 130348 215812 130354
rect 215850 130319 215906 130328
rect 215760 130290 215812 130296
rect 215208 53168 215260 53174
rect 215208 53110 215260 53116
rect 215220 44130 215248 53110
rect 215772 44538 215800 130290
rect 215864 129674 215892 130319
rect 215956 129742 215984 130426
rect 215944 129736 215996 129742
rect 215944 129678 215996 129684
rect 215852 129668 215904 129674
rect 215852 129610 215904 129616
rect 215864 127634 215892 129610
rect 215852 127628 215904 127634
rect 215852 127570 215904 127576
rect 215956 127514 215984 129678
rect 215864 127486 215984 127514
rect 215760 44532 215812 44538
rect 215760 44474 215812 44480
rect 215208 44124 215260 44130
rect 215208 44066 215260 44072
rect 215864 44062 215892 127486
rect 215944 127424 215996 127430
rect 215944 127366 215996 127372
rect 215852 44056 215904 44062
rect 215852 43998 215904 44004
rect 215116 42424 215168 42430
rect 215116 42366 215168 42372
rect 215024 40656 215076 40662
rect 215024 40598 215076 40604
rect 214840 39976 214892 39982
rect 214840 39918 214892 39924
rect 215956 39846 215984 127366
rect 216048 40866 216076 131038
rect 216140 44198 216168 150418
rect 216128 44192 216180 44198
rect 216128 44134 216180 44140
rect 216232 43858 216260 151302
rect 216324 130762 216352 240382
rect 216416 239970 216444 368834
rect 216508 262993 216536 373526
rect 216692 372745 216720 383166
rect 216784 375358 216812 408711
rect 217230 407824 217286 407833
rect 217230 407759 217286 407768
rect 216864 405000 216916 405006
rect 216862 404968 216864 404977
rect 216916 404968 216918 404977
rect 216862 404903 216918 404912
rect 216772 375352 216824 375358
rect 216772 375294 216824 375300
rect 216784 375086 216812 375294
rect 216772 375080 216824 375086
rect 216772 375022 216824 375028
rect 216876 373969 216904 404903
rect 217048 383580 217100 383586
rect 217048 383522 217100 383528
rect 217060 383081 217088 383522
rect 217046 383072 217102 383081
rect 217046 383007 217102 383016
rect 217046 375320 217102 375329
rect 217046 375255 217102 375264
rect 217060 375057 217088 375255
rect 217046 375048 217102 375057
rect 217244 375018 217272 407759
rect 217336 404297 217364 489126
rect 217322 404288 217378 404297
rect 217322 404223 217378 404232
rect 217046 374983 217102 374992
rect 217232 375012 217284 375018
rect 216862 373960 216918 373969
rect 216862 373895 216918 373904
rect 216678 372736 216734 372745
rect 216678 372671 216734 372680
rect 216586 369880 216642 369889
rect 216586 369815 216642 369824
rect 216494 262984 216550 262993
rect 216494 262919 216550 262928
rect 216404 239964 216456 239970
rect 216404 239906 216456 239912
rect 216416 151502 216444 239906
rect 216404 151496 216456 151502
rect 216404 151438 216456 151444
rect 216416 150482 216444 151438
rect 216496 151088 216548 151094
rect 216496 151030 216548 151036
rect 216404 150476 216456 150482
rect 216404 150418 216456 150424
rect 216508 142154 216536 151030
rect 216416 142126 216536 142154
rect 216312 130756 216364 130762
rect 216312 130698 216364 130704
rect 216220 43852 216272 43858
rect 216220 43794 216272 43800
rect 216036 40860 216088 40866
rect 216036 40802 216088 40808
rect 215944 39840 215996 39846
rect 215944 39782 215996 39788
rect 216324 39506 216352 130698
rect 216416 39914 216444 142126
rect 216496 133204 216548 133210
rect 216496 133146 216548 133152
rect 216508 41342 216536 133146
rect 216600 42634 216628 369815
rect 216772 349240 216824 349246
rect 216772 349182 216824 349188
rect 216678 298072 216734 298081
rect 216678 298007 216734 298016
rect 216692 277394 216720 298007
rect 216784 287054 216812 349182
rect 216876 294953 216904 373895
rect 216956 372904 217008 372910
rect 216956 372846 217008 372852
rect 216968 296041 216996 372846
rect 216954 296032 217010 296041
rect 216954 295967 217010 295976
rect 216968 295361 216996 295967
rect 216954 295352 217010 295361
rect 216954 295287 217010 295296
rect 216862 294944 216918 294953
rect 216862 294879 216918 294888
rect 216876 294001 216904 294879
rect 216862 293992 216918 294001
rect 216862 293927 216918 293936
rect 217060 293185 217088 374983
rect 217232 374954 217284 374960
rect 217244 373994 217272 374954
rect 217244 373966 217364 373994
rect 217232 369912 217284 369918
rect 217232 369854 217284 369860
rect 217138 301880 217194 301889
rect 217138 301815 217194 301824
rect 217046 293176 217102 293185
rect 217046 293111 217102 293120
rect 216784 287026 216904 287054
rect 216692 277366 216812 277394
rect 216680 276004 216732 276010
rect 216680 275946 216732 275952
rect 216692 274961 216720 275946
rect 216678 274952 216734 274961
rect 216678 274887 216734 274896
rect 216680 274644 216732 274650
rect 216680 274586 216732 274592
rect 216692 273329 216720 274586
rect 216678 273320 216734 273329
rect 216678 273255 216734 273264
rect 216680 273216 216732 273222
rect 216680 273158 216732 273164
rect 216692 273057 216720 273158
rect 216678 273048 216734 273057
rect 216678 272983 216734 272992
rect 216784 272626 216812 277366
rect 216692 272598 216812 272626
rect 216692 187785 216720 272598
rect 216876 258074 216904 287026
rect 216784 258046 216904 258074
rect 216784 241466 216812 258046
rect 216772 241460 216824 241466
rect 216772 241402 216824 241408
rect 217048 239624 217100 239630
rect 217048 239566 217100 239572
rect 216770 193216 216826 193225
rect 216770 193151 216826 193160
rect 216784 191865 216812 193151
rect 216770 191856 216826 191865
rect 216770 191791 216826 191800
rect 216678 187776 216734 187785
rect 216678 187711 216734 187720
rect 216680 165572 216732 165578
rect 216680 165514 216732 165520
rect 216692 165073 216720 165514
rect 216678 165064 216734 165073
rect 216678 164999 216734 165008
rect 216680 163532 216732 163538
rect 216680 163474 216732 163480
rect 216692 163441 216720 163474
rect 216678 163432 216734 163441
rect 216678 163367 216734 163376
rect 216784 81977 216812 191791
rect 216862 191720 216918 191729
rect 216862 191655 216918 191664
rect 216770 81968 216826 81977
rect 216770 81903 216826 81912
rect 216876 81025 216904 191655
rect 216954 185056 217010 185065
rect 216954 184991 217010 185000
rect 216862 81016 216918 81025
rect 216862 80951 216918 80960
rect 216968 75041 216996 184991
rect 217060 171134 217088 239566
rect 217152 193225 217180 301815
rect 217244 264654 217272 369854
rect 217336 298081 217364 373966
rect 217428 371074 217456 491982
rect 217600 482384 217652 482390
rect 217600 482326 217652 482332
rect 217508 463616 217560 463622
rect 217508 463558 217560 463564
rect 217416 371068 217468 371074
rect 217416 371010 217468 371016
rect 217520 368966 217548 463558
rect 217612 406065 217640 482326
rect 217784 467152 217836 467158
rect 217784 467094 217836 467100
rect 217692 462392 217744 462398
rect 217692 462334 217744 462340
rect 217704 412570 217732 462334
rect 217796 422294 217824 467094
rect 217796 422266 218008 422294
rect 217704 412542 217916 412570
rect 217888 411913 217916 412542
rect 217874 411904 217930 411913
rect 217874 411839 217930 411848
rect 217690 410952 217746 410961
rect 217690 410887 217746 410896
rect 217598 406056 217654 406065
rect 217598 405991 217654 406000
rect 217612 373998 217640 405991
rect 217600 373992 217652 373998
rect 217600 373934 217652 373940
rect 217612 372910 217640 373934
rect 217600 372904 217652 372910
rect 217600 372846 217652 372852
rect 217508 368960 217560 368966
rect 217508 368902 217560 368908
rect 217704 300937 217732 410887
rect 217784 375352 217836 375358
rect 217784 375294 217836 375300
rect 217690 300928 217746 300937
rect 217690 300863 217746 300872
rect 217322 298072 217378 298081
rect 217322 298007 217378 298016
rect 217506 295352 217562 295361
rect 217506 295287 217562 295296
rect 217414 293992 217470 294001
rect 217414 293927 217470 293936
rect 217232 264648 217284 264654
rect 217232 264590 217284 264596
rect 217232 239828 217284 239834
rect 217232 239770 217284 239776
rect 217138 193216 217194 193225
rect 217138 193151 217194 193160
rect 217060 171106 217180 171134
rect 217048 164212 217100 164218
rect 217048 164154 217100 164160
rect 217060 163169 217088 164154
rect 217046 163160 217102 163169
rect 217046 163095 217102 163104
rect 217152 151230 217180 171106
rect 217140 151224 217192 151230
rect 217140 151166 217192 151172
rect 216954 75032 217010 75041
rect 216954 74967 217010 74976
rect 216678 53272 216734 53281
rect 216678 53207 216734 53216
rect 216692 53174 216720 53207
rect 216680 53168 216732 53174
rect 216680 53110 216732 53116
rect 217152 44266 217180 151166
rect 217244 130218 217272 239770
rect 217428 185065 217456 293927
rect 217520 186017 217548 295287
rect 217600 240304 217652 240310
rect 217600 240246 217652 240252
rect 217506 186008 217562 186017
rect 217506 185943 217562 185952
rect 217414 185056 217470 185065
rect 217414 184991 217470 185000
rect 217414 183288 217470 183297
rect 217414 183223 217470 183232
rect 217232 130212 217284 130218
rect 217232 130154 217284 130160
rect 217244 44402 217272 130154
rect 217428 73273 217456 183223
rect 217520 76129 217548 185943
rect 217612 130898 217640 240246
rect 217704 191729 217732 300863
rect 217796 298761 217824 375294
rect 217888 301889 217916 411839
rect 217980 407833 218008 422266
rect 217966 407824 218022 407833
rect 217966 407759 218022 407768
rect 217966 404288 218022 404297
rect 217966 404223 218022 404232
rect 217980 403209 218008 404223
rect 217966 403200 218022 403209
rect 217966 403135 218022 403144
rect 217980 375329 218008 403135
rect 217966 375320 218022 375329
rect 217966 375255 218022 375264
rect 217968 373176 218020 373182
rect 217968 373118 218020 373124
rect 217874 301880 217930 301889
rect 217874 301815 217930 301824
rect 217782 298752 217838 298761
rect 217782 298687 217838 298696
rect 217690 191720 217746 191729
rect 217690 191655 217746 191664
rect 217704 191049 217732 191655
rect 217690 191040 217746 191049
rect 217690 190975 217746 190984
rect 217796 188737 217824 298687
rect 217874 293176 217930 293185
rect 217874 293111 217930 293120
rect 217782 188728 217838 188737
rect 217782 188663 217838 188672
rect 217600 130892 217652 130898
rect 217600 130834 217652 130840
rect 217506 76120 217562 76129
rect 217506 76055 217562 76064
rect 217414 73264 217470 73273
rect 217414 73199 217470 73208
rect 217232 44396 217284 44402
rect 217232 44338 217284 44344
rect 217140 44260 217192 44266
rect 217140 44202 217192 44208
rect 216588 42628 216640 42634
rect 216588 42570 216640 42576
rect 216496 41336 216548 41342
rect 216496 41278 216548 41284
rect 216404 39908 216456 39914
rect 216404 39850 216456 39856
rect 217612 39574 217640 130834
rect 217796 78849 217824 188663
rect 217888 183297 217916 293111
rect 217980 239834 218008 373118
rect 218072 372502 218100 492458
rect 218164 372881 218192 495023
rect 218348 492538 218376 495023
rect 218256 492510 218376 492538
rect 218808 492522 218836 495023
rect 219544 492794 219572 495037
rect 219636 495023 220018 495051
rect 220096 495023 220478 495051
rect 220954 495023 221044 495051
rect 219532 492788 219584 492794
rect 219532 492730 219584 492736
rect 219636 492674 219664 495023
rect 219452 492646 219664 492674
rect 218796 492516 218848 492522
rect 218256 374882 218284 492510
rect 218796 492458 218848 492464
rect 218336 492176 218388 492182
rect 218336 492118 218388 492124
rect 218244 374876 218296 374882
rect 218244 374818 218296 374824
rect 218256 374202 218284 374818
rect 218244 374196 218296 374202
rect 218244 374138 218296 374144
rect 218150 372872 218206 372881
rect 218150 372807 218206 372816
rect 218060 372496 218112 372502
rect 218060 372438 218112 372444
rect 218348 350441 218376 492118
rect 218796 487824 218848 487830
rect 218796 487766 218848 487772
rect 218702 465760 218758 465769
rect 218702 465695 218758 465704
rect 218428 462052 218480 462058
rect 218428 461994 218480 462000
rect 218440 369306 218468 461994
rect 218518 371104 218574 371113
rect 218518 371039 218574 371048
rect 218428 369300 218480 369306
rect 218428 369242 218480 369248
rect 218334 350432 218390 350441
rect 218334 350367 218390 350376
rect 218532 264790 218560 371039
rect 218610 369064 218666 369073
rect 218610 368999 218666 369008
rect 218624 264858 218652 368999
rect 218612 264852 218664 264858
rect 218612 264794 218664 264800
rect 218520 264784 218572 264790
rect 218520 264726 218572 264732
rect 218426 263664 218482 263673
rect 218426 263599 218482 263608
rect 218336 240712 218388 240718
rect 218336 240654 218388 240660
rect 217968 239828 218020 239834
rect 217968 239770 218020 239776
rect 217980 239358 218008 239770
rect 217968 239352 218020 239358
rect 217968 239294 218020 239300
rect 217966 187776 218022 187785
rect 217966 187711 218022 187720
rect 217874 183288 217930 183297
rect 217874 183223 217930 183232
rect 217782 78840 217838 78849
rect 217782 78775 217838 78784
rect 217980 77897 218008 187711
rect 218242 153096 218298 153105
rect 218242 153031 218298 153040
rect 217966 77888 218022 77897
rect 217966 77823 218022 77832
rect 218256 42702 218284 153031
rect 218348 130966 218376 240654
rect 218336 130960 218388 130966
rect 218336 130902 218388 130908
rect 218244 42696 218296 42702
rect 218244 42638 218296 42644
rect 218440 42294 218468 263599
rect 218612 240032 218664 240038
rect 218612 239974 218664 239980
rect 218520 239488 218572 239494
rect 218520 239430 218572 239436
rect 218532 238678 218560 239430
rect 218520 238672 218572 238678
rect 218520 238614 218572 238620
rect 218532 151026 218560 238614
rect 218624 151570 218652 239974
rect 218612 151564 218664 151570
rect 218612 151506 218664 151512
rect 218520 151020 218572 151026
rect 218520 150962 218572 150968
rect 218520 130416 218572 130422
rect 218520 130358 218572 130364
rect 218532 44334 218560 130358
rect 218612 130280 218664 130286
rect 218612 130222 218664 130228
rect 218624 44606 218652 130222
rect 218612 44600 218664 44606
rect 218612 44542 218664 44548
rect 218520 44328 218572 44334
rect 218520 44270 218572 44276
rect 218428 42288 218480 42294
rect 218428 42230 218480 42236
rect 218716 42158 218744 465695
rect 218808 152386 218836 487766
rect 218888 461780 218940 461786
rect 218888 461722 218940 461728
rect 218900 152862 218928 461722
rect 218980 459196 219032 459202
rect 218980 459138 219032 459144
rect 218992 263022 219020 459138
rect 219452 374354 219480 492646
rect 219532 492584 219584 492590
rect 220096 492538 220124 495023
rect 221016 492794 221044 495023
rect 221108 495023 221398 495051
rect 221476 495023 221766 495051
rect 222242 495023 222608 495051
rect 221004 492788 221056 492794
rect 221004 492730 221056 492736
rect 221108 492538 221136 495023
rect 221188 492788 221240 492794
rect 221188 492730 221240 492736
rect 219532 492526 219584 492532
rect 219360 374326 219480 374354
rect 219256 373720 219308 373726
rect 219256 373662 219308 373668
rect 219360 373674 219388 374326
rect 219438 374096 219494 374105
rect 219438 374031 219494 374040
rect 219452 373794 219480 374031
rect 219440 373788 219492 373794
rect 219440 373730 219492 373736
rect 219164 373244 219216 373250
rect 219164 373186 219216 373192
rect 219072 373108 219124 373114
rect 219072 373050 219124 373056
rect 218980 263016 219032 263022
rect 218980 262958 219032 262964
rect 218980 240916 219032 240922
rect 218980 240858 219032 240864
rect 218888 152856 218940 152862
rect 218888 152798 218940 152804
rect 218796 152380 218848 152386
rect 218796 152322 218848 152328
rect 218888 151020 218940 151026
rect 218888 150962 218940 150968
rect 218796 130960 218848 130966
rect 218796 130902 218848 130908
rect 218704 42152 218756 42158
rect 218704 42094 218756 42100
rect 218808 41002 218836 130902
rect 218900 43994 218928 150962
rect 218992 131102 219020 240858
rect 219084 239630 219112 373050
rect 219176 264926 219204 373186
rect 219268 372774 219296 373662
rect 219360 373646 219480 373674
rect 219348 373312 219400 373318
rect 219348 373254 219400 373260
rect 219360 372881 219388 373254
rect 219346 372872 219402 372881
rect 219346 372807 219402 372816
rect 219256 372768 219308 372774
rect 219256 372710 219308 372716
rect 219164 264920 219216 264926
rect 219164 264862 219216 264868
rect 219268 240038 219296 372710
rect 219452 372570 219480 373646
rect 219440 372564 219492 372570
rect 219440 372506 219492 372512
rect 219544 372201 219572 492526
rect 219636 492510 220124 492538
rect 220832 492510 221136 492538
rect 219636 374134 219664 492510
rect 219992 492380 220044 492386
rect 219992 492322 220044 492328
rect 219624 374128 219676 374134
rect 219624 374070 219676 374076
rect 219624 373788 219676 373794
rect 219624 373730 219676 373736
rect 219530 372192 219586 372201
rect 219530 372127 219586 372136
rect 219532 371952 219584 371958
rect 219532 371894 219584 371900
rect 219544 364334 219572 371894
rect 219636 369073 219664 373730
rect 219900 372224 219952 372230
rect 219900 372166 219952 372172
rect 219808 371884 219860 371890
rect 219808 371826 219860 371832
rect 219716 371544 219768 371550
rect 219716 371486 219768 371492
rect 219622 369064 219678 369073
rect 219622 368999 219678 369008
rect 219544 364306 219664 364334
rect 219348 350532 219400 350538
rect 219348 350474 219400 350480
rect 219360 240718 219388 350474
rect 219532 241392 219584 241398
rect 219532 241334 219584 241340
rect 219348 240712 219400 240718
rect 219348 240654 219400 240660
rect 219348 240236 219400 240242
rect 219348 240178 219400 240184
rect 219256 240032 219308 240038
rect 219256 239974 219308 239980
rect 219164 239828 219216 239834
rect 219164 239770 219216 239776
rect 219072 239624 219124 239630
rect 219072 239566 219124 239572
rect 219176 151162 219204 239770
rect 219256 151564 219308 151570
rect 219256 151506 219308 151512
rect 219164 151156 219216 151162
rect 219164 151098 219216 151104
rect 218980 131096 219032 131102
rect 218980 131038 219032 131044
rect 218980 130824 219032 130830
rect 218980 130766 219032 130772
rect 218992 45554 219020 130766
rect 219072 130552 219124 130558
rect 219072 130494 219124 130500
rect 219084 55214 219112 130494
rect 219268 55214 219296 151506
rect 219360 130830 219388 240178
rect 219440 151836 219492 151842
rect 219440 151778 219492 151784
rect 219452 151706 219480 151778
rect 219440 151700 219492 151706
rect 219440 151642 219492 151648
rect 219544 131034 219572 241334
rect 219636 241262 219664 364306
rect 219624 241256 219676 241262
rect 219624 241198 219676 241204
rect 219728 240446 219756 371486
rect 219820 241126 219848 371826
rect 219912 241194 219940 372166
rect 219900 241188 219952 241194
rect 219900 241130 219952 241136
rect 219808 241120 219860 241126
rect 219808 241062 219860 241068
rect 219716 240440 219768 240446
rect 219716 240382 219768 240388
rect 219900 240100 219952 240106
rect 219900 240042 219952 240048
rect 219808 239896 219860 239902
rect 219808 239838 219860 239844
rect 219624 239692 219676 239698
rect 219624 239634 219676 239640
rect 219636 151298 219664 239634
rect 219820 151706 219848 239838
rect 219808 151700 219860 151706
rect 219808 151642 219860 151648
rect 219912 151638 219940 240042
rect 219900 151632 219952 151638
rect 219900 151574 219952 151580
rect 219624 151292 219676 151298
rect 219624 151234 219676 151240
rect 219532 131028 219584 131034
rect 219532 130970 219584 130976
rect 219348 130824 219400 130830
rect 219348 130766 219400 130772
rect 219544 129810 219572 130970
rect 219532 129804 219584 129810
rect 219532 129746 219584 129752
rect 219084 55186 219204 55214
rect 219268 55186 219388 55214
rect 218992 45526 219112 45554
rect 218978 44840 219034 44849
rect 218978 44775 219034 44784
rect 218888 43988 218940 43994
rect 218888 43930 218940 43936
rect 218992 43450 219020 44775
rect 218980 43444 219032 43450
rect 218980 43386 219032 43392
rect 218796 40996 218848 41002
rect 218796 40938 218848 40944
rect 219084 40934 219112 45526
rect 219072 40928 219124 40934
rect 219072 40870 219124 40876
rect 217600 39568 217652 39574
rect 217600 39510 217652 39516
rect 216312 39500 216364 39506
rect 216312 39442 216364 39448
rect 219176 39438 219204 55186
rect 219254 44840 219310 44849
rect 219254 44775 219310 44784
rect 219268 43586 219296 44775
rect 219256 43580 219308 43586
rect 219256 43522 219308 43528
rect 219360 41070 219388 55186
rect 219636 43926 219664 151234
rect 219808 151156 219860 151162
rect 219808 151098 219860 151104
rect 219716 129804 219768 129810
rect 219716 129746 219768 129752
rect 219624 43920 219676 43926
rect 219624 43862 219676 43868
rect 219348 41064 219400 41070
rect 219348 41006 219400 41012
rect 219728 39642 219756 129746
rect 219820 39778 219848 151098
rect 219808 39772 219860 39778
rect 219808 39714 219860 39720
rect 219912 39710 219940 151574
rect 220004 41410 220032 492322
rect 220832 459610 220860 492510
rect 220912 492448 220964 492454
rect 220912 492390 220964 492396
rect 220924 459678 220952 492390
rect 221200 489914 221228 492730
rect 221476 492454 221504 495023
rect 221464 492448 221516 492454
rect 221464 492390 221516 492396
rect 222580 490618 222608 495023
rect 222672 492386 222700 495037
rect 223162 495023 223528 495051
rect 223622 495023 223712 495051
rect 222660 492380 222712 492386
rect 222660 492322 222712 492328
rect 223500 491978 223528 495023
rect 223580 492516 223632 492522
rect 223580 492458 223632 492464
rect 223488 491972 223540 491978
rect 223488 491914 223540 491920
rect 222568 490612 222620 490618
rect 222568 490554 222620 490560
rect 221016 489886 221228 489914
rect 220912 459672 220964 459678
rect 221016 459649 221044 489886
rect 223592 475425 223620 492458
rect 223684 486470 223712 495023
rect 223776 495023 223974 495051
rect 223776 492522 223804 495023
rect 224420 492561 224448 495037
rect 224406 492552 224462 492561
rect 223764 492516 223816 492522
rect 224406 492487 224462 492496
rect 223764 492458 223816 492464
rect 224880 491881 224908 495037
rect 225370 495023 225644 495051
rect 225738 495023 226104 495051
rect 225616 492046 225644 495023
rect 226076 492182 226104 495023
rect 226168 492250 226196 495037
rect 226156 492244 226208 492250
rect 226156 492186 226208 492192
rect 226064 492176 226116 492182
rect 226064 492118 226116 492124
rect 225604 492040 225656 492046
rect 225604 491982 225656 491988
rect 224866 491872 224922 491881
rect 224866 491807 224922 491816
rect 226432 487348 226484 487354
rect 226432 487290 226484 487296
rect 226340 486804 226392 486810
rect 226340 486746 226392 486752
rect 223672 486464 223724 486470
rect 223672 486406 223724 486412
rect 223578 475416 223634 475425
rect 223578 475351 223634 475360
rect 226352 465798 226380 486746
rect 226444 467265 226472 487290
rect 226628 485774 226656 495037
rect 226720 495023 227102 495051
rect 227272 495023 227562 495051
rect 227824 495023 227930 495051
rect 228008 495023 228390 495051
rect 228560 495023 228850 495051
rect 226720 487354 226748 495023
rect 226708 487348 226760 487354
rect 226708 487290 226760 487296
rect 227272 486810 227300 495023
rect 227824 492674 227852 495023
rect 228008 492674 228036 495023
rect 227640 492646 227852 492674
rect 227916 492646 228036 492674
rect 227640 487830 227668 492646
rect 227916 487914 227944 492646
rect 227732 487886 227944 487914
rect 227628 487824 227680 487830
rect 227628 487766 227680 487772
rect 227260 486804 227312 486810
rect 227260 486746 227312 486752
rect 226536 485746 226656 485774
rect 226536 476814 226564 485746
rect 226524 476808 226576 476814
rect 226524 476750 226576 476756
rect 226430 467256 226486 467265
rect 226430 467191 226486 467200
rect 226340 465792 226392 465798
rect 226340 465734 226392 465740
rect 227732 465730 227760 487886
rect 227812 487824 227864 487830
rect 227812 487766 227864 487772
rect 227824 467158 227852 487766
rect 228560 485774 228588 495023
rect 229100 494964 229152 494970
rect 229100 494906 229152 494912
rect 227916 485746 228588 485774
rect 227916 475386 227944 485746
rect 229112 482322 229140 494906
rect 229312 494850 229340 495037
rect 229480 495023 229770 495051
rect 229848 495023 230138 495051
rect 230492 495023 230598 495051
rect 231074 495023 231440 495051
rect 231534 495023 231808 495051
rect 231902 495023 231992 495051
rect 229480 494970 229508 495023
rect 229468 494964 229520 494970
rect 229468 494906 229520 494912
rect 229312 494822 229508 494850
rect 229192 486872 229244 486878
rect 229192 486814 229244 486820
rect 229204 483721 229232 486814
rect 229480 485774 229508 494822
rect 229848 486878 229876 495023
rect 229836 486872 229888 486878
rect 229836 486814 229888 486820
rect 229296 485746 229508 485774
rect 229296 485110 229324 485746
rect 229284 485104 229336 485110
rect 229284 485046 229336 485052
rect 229190 483712 229246 483721
rect 229190 483647 229246 483656
rect 229100 482316 229152 482322
rect 229100 482258 229152 482264
rect 230492 480962 230520 495023
rect 231412 492250 231440 495023
rect 231400 492244 231452 492250
rect 231400 492186 231452 492192
rect 231780 492114 231808 495023
rect 231768 492108 231820 492114
rect 231768 492050 231820 492056
rect 231860 490408 231912 490414
rect 231860 490350 231912 490356
rect 230480 480956 230532 480962
rect 230480 480898 230532 480904
rect 231872 478145 231900 490350
rect 231964 479505 231992 495023
rect 232332 492017 232360 495037
rect 232424 495023 232806 495051
rect 232318 492008 232374 492017
rect 232318 491943 232374 491952
rect 232424 490414 232452 495023
rect 233252 492153 233280 495037
rect 233344 495023 233726 495051
rect 234110 495023 234200 495051
rect 233238 492144 233294 492153
rect 233238 492079 233294 492088
rect 232412 490408 232464 490414
rect 232412 490350 232464 490356
rect 233240 490408 233292 490414
rect 233240 490350 233292 490356
rect 231950 479496 232006 479505
rect 231950 479431 232006 479440
rect 231858 478136 231914 478145
rect 231858 478071 231914 478080
rect 227904 475380 227956 475386
rect 227904 475322 227956 475328
rect 227812 467152 227864 467158
rect 233252 467129 233280 490350
rect 233344 472569 233372 495023
rect 234172 491881 234200 495023
rect 234264 495023 234554 495051
rect 235030 495023 235304 495051
rect 235490 495023 235856 495051
rect 234158 491872 234214 491881
rect 234158 491807 234214 491816
rect 234264 490414 234292 495023
rect 235276 492289 235304 495023
rect 235828 492425 235856 495023
rect 235920 492561 235948 495037
rect 236318 495023 236592 495051
rect 235906 492552 235962 492561
rect 235906 492487 235962 492496
rect 235814 492416 235870 492425
rect 235814 492351 235870 492360
rect 235262 492280 235318 492289
rect 235262 492215 235318 492224
rect 234252 490408 234304 490414
rect 234252 490350 234304 490356
rect 236564 487801 236592 495023
rect 236748 489258 236776 495037
rect 236840 495023 237222 495051
rect 236736 489252 236788 489258
rect 236736 489194 236788 489200
rect 236550 487792 236606 487801
rect 236550 487727 236606 487736
rect 236840 485774 236868 495023
rect 237472 490476 237524 490482
rect 237472 490418 237524 490424
rect 237380 490408 237432 490414
rect 237380 490350 237432 490356
rect 236012 485746 236868 485774
rect 236012 482390 236040 485746
rect 236000 482384 236052 482390
rect 236000 482326 236052 482332
rect 233330 472560 233386 472569
rect 233330 472495 233386 472504
rect 227812 467094 227864 467100
rect 233238 467120 233294 467129
rect 233238 467055 233294 467064
rect 227720 465724 227772 465730
rect 227720 465666 227772 465672
rect 237392 460222 237420 490350
rect 237484 474026 237512 490418
rect 237668 485774 237696 495037
rect 237760 495023 238142 495051
rect 238220 495023 238510 495051
rect 238986 495023 239352 495051
rect 239446 495023 239720 495051
rect 239906 495023 240088 495051
rect 240274 495023 240640 495051
rect 240734 495023 240824 495051
rect 237760 490482 237788 495023
rect 237748 490476 237800 490482
rect 237748 490418 237800 490424
rect 238220 490414 238248 495023
rect 238208 490408 238260 490414
rect 238208 490350 238260 490356
rect 239324 489190 239352 495023
rect 239692 492454 239720 495023
rect 240060 492590 240088 495023
rect 240048 492584 240100 492590
rect 240048 492526 240100 492532
rect 239680 492448 239732 492454
rect 239680 492390 239732 492396
rect 240612 492318 240640 495023
rect 240796 492386 240824 495023
rect 240888 495023 241178 495051
rect 241532 495023 241638 495051
rect 240784 492380 240836 492386
rect 240784 492322 240836 492328
rect 240600 492312 240652 492318
rect 240600 492254 240652 492260
rect 239312 489184 239364 489190
rect 239312 489126 239364 489132
rect 240888 485774 240916 495023
rect 237576 485746 237696 485774
rect 240152 485746 240916 485774
rect 237576 483682 237604 485746
rect 237564 483676 237616 483682
rect 237564 483618 237616 483624
rect 237472 474020 237524 474026
rect 237472 473962 237524 473968
rect 240152 463010 240180 485746
rect 241532 463146 241560 495023
rect 242084 486538 242112 495037
rect 242176 495023 242466 495051
rect 242072 486532 242124 486538
rect 242072 486474 242124 486480
rect 242176 485774 242204 495023
rect 242928 494834 242956 495037
rect 243004 495023 243386 495051
rect 243464 495023 243846 495051
rect 244322 495023 244504 495051
rect 242916 494828 242968 494834
rect 242916 494770 242968 494776
rect 242900 490408 242952 490414
rect 242900 490350 242952 490356
rect 241624 485746 242204 485774
rect 241624 469946 241652 485746
rect 241612 469940 241664 469946
rect 241612 469882 241664 469888
rect 241520 463140 241572 463146
rect 241520 463082 241572 463088
rect 240140 463004 240192 463010
rect 240140 462946 240192 462952
rect 242912 460426 242940 490350
rect 243004 481098 243032 495023
rect 243084 494828 243136 494834
rect 243084 494770 243136 494776
rect 243096 485178 243124 494770
rect 243464 490414 243492 495023
rect 244372 494828 244424 494834
rect 244372 494770 244424 494776
rect 244384 490498 244412 494770
rect 244476 494714 244504 495023
rect 244568 495023 244674 495051
rect 244752 495023 245134 495051
rect 245304 495023 245594 495051
rect 245764 495023 246054 495051
rect 246438 495023 246528 495051
rect 244568 494834 244596 495023
rect 244556 494828 244608 494834
rect 244556 494770 244608 494776
rect 244476 494686 244688 494714
rect 244292 490470 244412 490498
rect 243452 490408 243504 490414
rect 243452 490350 243504 490356
rect 243084 485172 243136 485178
rect 243084 485114 243136 485120
rect 242992 481092 243044 481098
rect 242992 481034 243044 481040
rect 244292 474094 244320 490470
rect 244372 490408 244424 490414
rect 244372 490350 244424 490356
rect 244384 476882 244412 490350
rect 244660 490210 244688 494686
rect 244648 490204 244700 490210
rect 244648 490146 244700 490152
rect 244556 490000 244608 490006
rect 244556 489942 244608 489948
rect 244464 487824 244516 487830
rect 244464 487766 244516 487772
rect 244476 478174 244504 487766
rect 244568 479534 244596 489942
rect 244752 487830 244780 495023
rect 245304 490414 245332 495023
rect 245292 490408 245344 490414
rect 245292 490350 245344 490356
rect 245660 490408 245712 490414
rect 245660 490350 245712 490356
rect 244740 487824 244792 487830
rect 244740 487766 244792 487772
rect 244556 479528 244608 479534
rect 244556 479470 244608 479476
rect 244464 478168 244516 478174
rect 244464 478110 244516 478116
rect 244372 476876 244424 476882
rect 244372 476818 244424 476824
rect 244280 474088 244332 474094
rect 244280 474030 244332 474036
rect 242900 460420 242952 460426
rect 242900 460362 242952 460368
rect 237380 460216 237432 460222
rect 237380 460158 237432 460164
rect 220912 459614 220964 459620
rect 221002 459640 221058 459649
rect 220820 459604 220872 459610
rect 221002 459575 221058 459584
rect 220820 459546 220872 459552
rect 245672 458862 245700 490350
rect 245764 472734 245792 495023
rect 246500 490686 246528 495023
rect 246592 495023 246882 495051
rect 246488 490680 246540 490686
rect 246488 490622 246540 490628
rect 246592 490414 246620 495023
rect 246580 490408 246632 490414
rect 246580 490350 246632 490356
rect 247328 489326 247356 495037
rect 247420 495023 247802 495051
rect 247880 495023 248262 495051
rect 247316 489320 247368 489326
rect 247316 489262 247368 489268
rect 247420 489138 247448 495023
rect 247052 489110 247448 489138
rect 245752 472728 245804 472734
rect 245752 472670 245804 472676
rect 247052 458930 247080 489110
rect 247880 485774 247908 495023
rect 248616 492726 248644 495037
rect 248708 495023 249090 495051
rect 249168 495023 249550 495051
rect 249904 495023 250010 495051
rect 250088 495023 250470 495051
rect 250548 495023 250838 495051
rect 251192 495023 251298 495051
rect 251376 495023 251758 495051
rect 251928 495023 252218 495051
rect 248604 492720 248656 492726
rect 248604 492662 248656 492668
rect 248708 490362 248736 495023
rect 247144 485746 247908 485774
rect 248432 490334 248736 490362
rect 247144 468586 247172 485746
rect 247132 468580 247184 468586
rect 247132 468522 247184 468528
rect 248432 460630 248460 490334
rect 249168 485774 249196 495023
rect 249800 490408 249852 490414
rect 249800 490350 249852 490356
rect 248524 485746 249196 485774
rect 248420 460624 248472 460630
rect 248420 460566 248472 460572
rect 248524 460290 248552 485746
rect 249812 460562 249840 490350
rect 249800 460556 249852 460562
rect 249800 460498 249852 460504
rect 249904 460358 249932 495023
rect 250088 485774 250116 495023
rect 250548 490414 250576 495023
rect 250536 490408 250588 490414
rect 250536 490350 250588 490356
rect 249996 485746 250116 485774
rect 249996 460494 250024 485746
rect 251192 463078 251220 495023
rect 251376 490362 251404 495023
rect 251284 490334 251404 490362
rect 251284 470014 251312 490334
rect 251928 485774 251956 495023
rect 251376 485746 251956 485774
rect 251376 471306 251404 485746
rect 252572 475454 252600 495037
rect 252664 495023 253046 495051
rect 253216 495023 253506 495051
rect 252664 478242 252692 495023
rect 253216 485774 253244 495023
rect 253952 491910 253980 495037
rect 254044 495023 254426 495051
rect 254504 495023 254794 495051
rect 254872 495023 255254 495051
rect 255516 495023 255714 495051
rect 255792 495023 256174 495051
rect 256344 495023 256634 495051
rect 256896 495023 257002 495051
rect 257080 495023 257462 495051
rect 257632 495023 257922 495051
rect 258276 495023 258382 495051
rect 258552 495023 258842 495051
rect 258920 495023 259210 495051
rect 253940 491904 253992 491910
rect 253940 491846 253992 491852
rect 253940 491768 253992 491774
rect 253940 491710 253992 491716
rect 252756 485746 253244 485774
rect 252756 479602 252784 485746
rect 252744 479596 252796 479602
rect 252744 479538 252796 479544
rect 252652 478236 252704 478242
rect 252652 478178 252704 478184
rect 252560 475448 252612 475454
rect 252560 475390 252612 475396
rect 251364 471300 251416 471306
rect 251364 471242 251416 471248
rect 251272 470008 251324 470014
rect 251272 469950 251324 469956
rect 251180 463072 251232 463078
rect 251180 463014 251232 463020
rect 249984 460488 250036 460494
rect 249984 460430 250036 460436
rect 249892 460352 249944 460358
rect 249892 460294 249944 460300
rect 248512 460284 248564 460290
rect 248512 460226 248564 460232
rect 253952 458998 253980 491710
rect 254044 468926 254072 495023
rect 254504 492538 254532 495023
rect 254136 492510 254532 492538
rect 254032 468920 254084 468926
rect 254032 468862 254084 468868
rect 254136 468790 254164 492510
rect 254216 491904 254268 491910
rect 254216 491846 254268 491852
rect 254228 481030 254256 491846
rect 254872 491774 254900 495023
rect 255320 492652 255372 492658
rect 255320 492594 255372 492600
rect 254860 491768 254912 491774
rect 254860 491710 254912 491716
rect 254216 481024 254268 481030
rect 254216 480966 254268 480972
rect 255332 468858 255360 492594
rect 255412 492584 255464 492590
rect 255412 492526 255464 492532
rect 255320 468852 255372 468858
rect 255320 468794 255372 468800
rect 254124 468784 254176 468790
rect 254124 468726 254176 468732
rect 255424 468654 255452 492526
rect 255516 468722 255544 495023
rect 255792 492590 255820 495023
rect 256344 492658 256372 495023
rect 256332 492652 256384 492658
rect 256332 492594 256384 492600
rect 256700 492652 256752 492658
rect 256700 492594 256752 492600
rect 255780 492584 255832 492590
rect 255780 492526 255832 492532
rect 256712 476950 256740 492594
rect 256792 491904 256844 491910
rect 256792 491846 256844 491852
rect 256804 478310 256832 491846
rect 256896 485246 256924 495023
rect 257080 492658 257108 495023
rect 257068 492652 257120 492658
rect 257068 492594 257120 492600
rect 257632 491910 257660 495023
rect 258172 492720 258224 492726
rect 258172 492662 258224 492668
rect 258080 492652 258132 492658
rect 258080 492594 258132 492600
rect 257620 491904 257672 491910
rect 257620 491846 257672 491852
rect 256884 485240 256936 485246
rect 256884 485182 256936 485188
rect 256792 478304 256844 478310
rect 256792 478246 256844 478252
rect 256700 476944 256752 476950
rect 256700 476886 256752 476892
rect 255504 468716 255556 468722
rect 255504 468658 255556 468664
rect 255412 468648 255464 468654
rect 255412 468590 255464 468596
rect 258092 460698 258120 492594
rect 258184 462913 258212 492662
rect 258276 472802 258304 495023
rect 258552 492658 258580 495023
rect 258920 492726 258948 495023
rect 259552 494964 259604 494970
rect 259552 494906 259604 494912
rect 258908 492720 258960 492726
rect 258908 492662 258960 492668
rect 258540 492652 258592 492658
rect 258540 492594 258592 492600
rect 259460 492652 259512 492658
rect 259460 492594 259512 492600
rect 258264 472796 258316 472802
rect 258264 472738 258316 472744
rect 259472 468994 259500 492594
rect 259564 471374 259592 494906
rect 259672 494850 259700 495037
rect 259840 495023 260130 495051
rect 260208 495023 260590 495051
rect 259840 494970 259868 495023
rect 259828 494964 259880 494970
rect 259828 494906 259880 494912
rect 259672 494822 259868 494850
rect 259840 489954 259868 494822
rect 260208 492658 260236 495023
rect 260196 492652 260248 492658
rect 260196 492594 260248 492600
rect 260840 492652 260892 492658
rect 260840 492594 260892 492600
rect 259672 489926 259868 489954
rect 259672 489914 259700 489926
rect 259656 489886 259700 489914
rect 259656 474162 259684 489886
rect 259644 474156 259696 474162
rect 259644 474098 259696 474104
rect 259552 471368 259604 471374
rect 259552 471310 259604 471316
rect 259460 468988 259512 468994
rect 259460 468930 259512 468936
rect 260852 465866 260880 492594
rect 260944 490754 260972 495037
rect 261036 495023 261418 495051
rect 261496 495023 261878 495051
rect 262354 495023 262444 495051
rect 260932 490748 260984 490754
rect 260932 490690 260984 490696
rect 261036 489914 261064 495023
rect 261496 492658 261524 495023
rect 262416 492726 262444 495023
rect 262508 495023 262798 495051
rect 262876 495023 263166 495051
rect 262404 492720 262456 492726
rect 262404 492662 262456 492668
rect 261484 492652 261536 492658
rect 261484 492594 261536 492600
rect 262220 492652 262272 492658
rect 262220 492594 262272 492600
rect 260944 489886 261064 489914
rect 260944 487830 260972 489886
rect 260932 487824 260984 487830
rect 260932 487766 260984 487772
rect 260840 465860 260892 465866
rect 260840 465802 260892 465808
rect 262232 463214 262260 492594
rect 262508 492538 262536 495023
rect 262588 492720 262640 492726
rect 262588 492662 262640 492668
rect 262324 492510 262536 492538
rect 262324 475522 262352 492510
rect 262600 492402 262628 492662
rect 262876 492658 262904 495023
rect 262864 492652 262916 492658
rect 262864 492594 262916 492600
rect 262416 492374 262628 492402
rect 262416 482458 262444 492374
rect 262404 482452 262456 482458
rect 262404 482394 262456 482400
rect 262312 475516 262364 475522
rect 262312 475458 262364 475464
rect 263612 463282 263640 495037
rect 263704 495023 264086 495051
rect 264256 495023 264546 495051
rect 265022 495023 265112 495051
rect 263704 466070 263732 495023
rect 264256 489914 264284 495023
rect 264980 492652 265032 492658
rect 264980 492594 265032 492600
rect 263796 489886 264284 489914
rect 263796 466138 263824 489886
rect 263784 466132 263836 466138
rect 263784 466074 263836 466080
rect 263692 466064 263744 466070
rect 263692 466006 263744 466012
rect 263600 463276 263652 463282
rect 263600 463218 263652 463224
rect 262220 463208 262272 463214
rect 262220 463150 262272 463156
rect 258170 462904 258226 462913
rect 258170 462839 258226 462848
rect 258080 460692 258132 460698
rect 258080 460634 258132 460640
rect 264992 459066 265020 492594
rect 265084 465769 265112 495023
rect 265176 495023 265374 495051
rect 265544 495023 265834 495051
rect 265912 495023 266294 495051
rect 266372 495023 266754 495051
rect 265176 465934 265204 495023
rect 265544 489914 265572 495023
rect 265912 492658 265940 495023
rect 265900 492652 265952 492658
rect 265900 492594 265952 492600
rect 265268 489886 265572 489914
rect 265268 466002 265296 489886
rect 265256 465996 265308 466002
rect 265256 465938 265308 465944
rect 265164 465928 265216 465934
rect 265164 465870 265216 465876
rect 265070 465760 265126 465769
rect 265070 465695 265126 465704
rect 266372 460834 266400 495023
rect 267108 490822 267136 495037
rect 267200 495023 267582 495051
rect 267752 495023 268042 495051
rect 268120 495023 268502 495051
rect 268672 495023 268962 495051
rect 269224 495023 269330 495051
rect 269408 495023 269790 495051
rect 269960 495023 270250 495051
rect 270512 495023 270710 495051
rect 270880 495023 271170 495051
rect 271248 495023 271538 495051
rect 271892 495023 271998 495051
rect 272076 495023 272458 495051
rect 272536 495023 272918 495051
rect 267096 490816 267148 490822
rect 267096 490758 267148 490764
rect 267200 489914 267228 495023
rect 266464 489886 267228 489914
rect 266464 469130 266492 489886
rect 267752 471578 267780 495023
rect 267832 492652 267884 492658
rect 267832 492594 267884 492600
rect 267844 474570 267872 492594
rect 268120 489914 268148 495023
rect 268672 492658 268700 495023
rect 268660 492652 268712 492658
rect 268660 492594 268712 492600
rect 269120 492652 269172 492658
rect 269120 492594 269172 492600
rect 267936 489886 268148 489914
rect 267832 474564 267884 474570
rect 267832 474506 267884 474512
rect 267936 474434 267964 489886
rect 267924 474428 267976 474434
rect 267924 474370 267976 474376
rect 267740 471572 267792 471578
rect 267740 471514 267792 471520
rect 266452 469124 266504 469130
rect 266452 469066 266504 469072
rect 269132 463350 269160 492594
rect 269224 474230 269252 495023
rect 269408 489914 269436 495023
rect 269960 492658 269988 495023
rect 269948 492652 270000 492658
rect 269948 492594 270000 492600
rect 269316 489886 269436 489914
rect 269316 474298 269344 489886
rect 269304 474292 269356 474298
rect 269304 474234 269356 474240
rect 269212 474224 269264 474230
rect 269212 474166 269264 474172
rect 269120 463344 269172 463350
rect 269120 463286 269172 463292
rect 266360 460828 266412 460834
rect 266360 460770 266412 460776
rect 270512 459202 270540 495023
rect 270592 492652 270644 492658
rect 270592 492594 270644 492600
rect 270604 474366 270632 492594
rect 270880 489914 270908 495023
rect 271248 492658 271276 495023
rect 271236 492652 271288 492658
rect 271236 492594 271288 492600
rect 270696 489886 270908 489914
rect 270696 474502 270724 489886
rect 270684 474496 270736 474502
rect 270684 474438 270736 474444
rect 270592 474360 270644 474366
rect 270592 474302 270644 474308
rect 271892 461854 271920 495023
rect 271972 492652 272024 492658
rect 271972 492594 272024 492600
rect 271984 466206 272012 492594
rect 272076 471510 272104 495023
rect 272536 492658 272564 495023
rect 273288 494834 273316 495037
rect 273364 495023 273746 495051
rect 273824 495023 274206 495051
rect 274682 495023 274772 495051
rect 273276 494828 273328 494834
rect 273276 494770 273328 494776
rect 272524 492652 272576 492658
rect 272524 492594 272576 492600
rect 273260 490408 273312 490414
rect 273260 490350 273312 490356
rect 272064 471504 272116 471510
rect 272064 471446 272116 471452
rect 271972 466200 272024 466206
rect 271972 466142 272024 466148
rect 271880 461848 271932 461854
rect 271880 461790 271932 461796
rect 270500 459196 270552 459202
rect 270500 459138 270552 459144
rect 273272 459134 273300 490350
rect 273364 471442 273392 495023
rect 273444 494828 273496 494834
rect 273444 494770 273496 494776
rect 273456 471918 273484 494770
rect 273824 490414 273852 495023
rect 273812 490408 273864 490414
rect 273812 490350 273864 490356
rect 274640 490408 274692 490414
rect 274640 490350 274692 490356
rect 273444 471912 273496 471918
rect 273444 471854 273496 471860
rect 273352 471436 273404 471442
rect 273352 471378 273404 471384
rect 274652 459270 274680 490350
rect 274744 461650 274772 495023
rect 275020 495023 275126 495051
rect 275204 495023 275494 495051
rect 275664 495023 275954 495051
rect 276216 495023 276414 495051
rect 276584 495023 276874 495051
rect 276952 495023 277334 495051
rect 277412 495023 277702 495051
rect 277872 495023 278162 495051
rect 278240 495023 278622 495051
rect 278792 495023 279082 495051
rect 279160 495023 279542 495051
rect 279620 495023 279910 495051
rect 280264 495023 280370 495051
rect 280448 495023 280830 495051
rect 281000 495023 281290 495051
rect 274824 490476 274876 490482
rect 274824 490418 274876 490424
rect 274836 464438 274864 490418
rect 275020 485774 275048 495023
rect 275204 490482 275232 495023
rect 275192 490476 275244 490482
rect 275192 490418 275244 490424
rect 275664 490414 275692 495023
rect 276020 490476 276072 490482
rect 276020 490418 276072 490424
rect 275652 490408 275704 490414
rect 275652 490350 275704 490356
rect 274928 485746 275048 485774
rect 274928 471714 274956 485746
rect 274916 471708 274968 471714
rect 274916 471650 274968 471656
rect 274824 464432 274876 464438
rect 274824 464374 274876 464380
rect 276032 463418 276060 490418
rect 276112 490408 276164 490414
rect 276112 490350 276164 490356
rect 276124 469062 276152 490350
rect 276216 471850 276244 495023
rect 276584 490414 276612 495023
rect 276952 490482 276980 495023
rect 276940 490476 276992 490482
rect 276940 490418 276992 490424
rect 276572 490408 276624 490414
rect 276572 490350 276624 490356
rect 276204 471844 276256 471850
rect 276204 471786 276256 471792
rect 276112 469056 276164 469062
rect 276112 468998 276164 469004
rect 277412 463486 277440 495023
rect 277492 490408 277544 490414
rect 277492 490350 277544 490356
rect 277504 463622 277532 490350
rect 277872 485774 277900 495023
rect 278240 490414 278268 495023
rect 278228 490408 278280 490414
rect 278228 490350 278280 490356
rect 277596 485746 277900 485774
rect 277596 471782 277624 485746
rect 277584 471776 277636 471782
rect 277584 471718 277636 471724
rect 277492 463616 277544 463622
rect 277492 463558 277544 463564
rect 277400 463480 277452 463486
rect 277400 463422 277452 463428
rect 276020 463412 276072 463418
rect 276020 463354 276072 463360
rect 278792 462058 278820 495023
rect 279160 490362 279188 495023
rect 278884 490334 279188 490362
rect 278884 471209 278912 490334
rect 279620 485774 279648 495023
rect 280160 490408 280212 490414
rect 280160 490350 280212 490356
rect 278976 485746 279648 485774
rect 278976 474065 279004 485746
rect 278962 474056 279018 474065
rect 278962 473991 279018 474000
rect 278870 471200 278926 471209
rect 278870 471135 278926 471144
rect 278780 462052 278832 462058
rect 278780 461994 278832 462000
rect 274732 461644 274784 461650
rect 274732 461586 274784 461592
rect 280172 460154 280200 490350
rect 280264 461786 280292 495023
rect 280448 485774 280476 495023
rect 281000 490414 281028 495023
rect 281660 494850 281688 495037
rect 281920 495023 282118 495051
rect 282288 495023 282578 495051
rect 283054 495023 283144 495051
rect 281660 494822 281856 494850
rect 280988 490408 281040 490414
rect 280988 490350 281040 490356
rect 281828 489394 281856 494822
rect 281816 489388 281868 489394
rect 281816 489330 281868 489336
rect 281920 489274 281948 495023
rect 280356 485746 280476 485774
rect 281552 489246 281948 489274
rect 280356 466410 280384 485746
rect 280344 466404 280396 466410
rect 280344 466346 280396 466352
rect 280252 461780 280304 461786
rect 280252 461722 280304 461728
rect 281552 460766 281580 489246
rect 282288 485774 282316 495023
rect 283012 492720 283064 492726
rect 283012 492662 283064 492668
rect 282920 492652 282972 492658
rect 282920 492594 282972 492600
rect 281644 485746 282316 485774
rect 281644 477086 281672 485746
rect 281632 477080 281684 477086
rect 281632 477022 281684 477028
rect 281540 460760 281592 460766
rect 281540 460702 281592 460708
rect 280160 460148 280212 460154
rect 280160 460090 280212 460096
rect 282932 459406 282960 492594
rect 283024 462126 283052 492662
rect 283116 487898 283144 495023
rect 283208 495023 283498 495051
rect 283576 495023 283866 495051
rect 283208 492658 283236 495023
rect 283576 492726 283604 495023
rect 284328 494834 284356 495037
rect 284404 495023 284786 495051
rect 284864 495023 285246 495051
rect 285722 495023 285812 495051
rect 284316 494828 284368 494834
rect 284316 494770 284368 494776
rect 283564 492720 283616 492726
rect 283564 492662 283616 492668
rect 283196 492652 283248 492658
rect 283196 492594 283248 492600
rect 284300 492652 284352 492658
rect 284300 492594 284352 492600
rect 283104 487892 283156 487898
rect 283104 487834 283156 487840
rect 284312 470082 284340 492594
rect 284404 471646 284432 495023
rect 284484 494828 284536 494834
rect 284484 494770 284536 494776
rect 284496 479670 284524 494770
rect 284864 492658 284892 495023
rect 284852 492652 284904 492658
rect 284852 492594 284904 492600
rect 285680 492652 285732 492658
rect 285680 492594 285732 492600
rect 284484 479664 284536 479670
rect 284484 479606 284536 479612
rect 284392 471640 284444 471646
rect 284392 471582 284444 471588
rect 284300 470076 284352 470082
rect 284300 470018 284352 470024
rect 283012 462120 283064 462126
rect 283012 462062 283064 462068
rect 285692 461922 285720 492594
rect 285784 464370 285812 495023
rect 285876 495023 286074 495051
rect 286152 495023 286534 495051
rect 286704 495023 286994 495051
rect 287072 495023 287454 495051
rect 287532 495023 287822 495051
rect 287992 495023 288282 495051
rect 288544 495023 288742 495051
rect 288912 495023 289202 495051
rect 289280 495023 289662 495051
rect 289832 495023 290030 495051
rect 290108 495023 290490 495051
rect 290568 495023 290950 495051
rect 285876 469198 285904 495023
rect 286152 489914 286180 495023
rect 286704 492658 286732 495023
rect 286692 492652 286744 492658
rect 286692 492594 286744 492600
rect 285968 489886 286180 489914
rect 285968 477154 285996 489886
rect 285956 477148 286008 477154
rect 285956 477090 286008 477096
rect 285864 469192 285916 469198
rect 285864 469134 285916 469140
rect 285772 464364 285824 464370
rect 285772 464306 285824 464312
rect 287072 461990 287100 495023
rect 287532 492538 287560 495023
rect 287164 492510 287560 492538
rect 287164 464506 287192 492510
rect 287992 489914 288020 495023
rect 288440 492652 288492 492658
rect 288440 492594 288492 492600
rect 287256 489886 288020 489914
rect 287256 479738 287284 489886
rect 287244 479732 287296 479738
rect 287244 479674 287296 479680
rect 287152 464500 287204 464506
rect 287152 464442 287204 464448
rect 287060 461984 287112 461990
rect 287060 461926 287112 461932
rect 285680 461916 285732 461922
rect 285680 461858 285732 461864
rect 282920 459400 282972 459406
rect 282920 459342 282972 459348
rect 288452 459338 288480 492594
rect 288544 463554 288572 495023
rect 288912 489914 288940 495023
rect 289280 492658 289308 495023
rect 289268 492652 289320 492658
rect 289268 492594 289320 492600
rect 288636 489886 288940 489914
rect 288636 468450 288664 489886
rect 288624 468444 288676 468450
rect 288624 468386 288676 468392
rect 289832 466274 289860 495023
rect 290108 492538 290136 495023
rect 289924 492510 290136 492538
rect 289924 474638 289952 492510
rect 290568 489914 290596 495023
rect 291200 492720 291252 492726
rect 291200 492662 291252 492668
rect 290016 489886 290596 489914
rect 290016 477018 290044 489886
rect 290004 477012 290056 477018
rect 290004 476954 290056 476960
rect 289912 474632 289964 474638
rect 289912 474574 289964 474580
rect 289820 466268 289872 466274
rect 289820 466210 289872 466216
rect 288532 463548 288584 463554
rect 288532 463490 288584 463496
rect 291212 459474 291240 492662
rect 291292 492652 291344 492658
rect 291292 492594 291344 492600
rect 291304 477222 291332 492594
rect 291396 477290 291424 495037
rect 291488 495023 291870 495051
rect 291948 495023 292238 495051
rect 291488 492658 291516 495023
rect 291948 492726 291976 495023
rect 291936 492720 291988 492726
rect 291936 492662 291988 492668
rect 291476 492652 291528 492658
rect 291476 492594 291528 492600
rect 292580 491836 292632 491842
rect 292580 491778 292632 491784
rect 291384 477284 291436 477290
rect 291384 477226 291436 477232
rect 291292 477216 291344 477222
rect 291292 477158 291344 477164
rect 292592 476785 292620 491778
rect 292684 477494 292712 495037
rect 292776 495023 293158 495051
rect 293328 495023 293618 495051
rect 292776 491842 292804 495023
rect 292764 491836 292816 491842
rect 292764 491778 292816 491784
rect 293328 489914 293356 495023
rect 292776 489886 293356 489914
rect 292776 483750 292804 489886
rect 292764 483744 292816 483750
rect 292764 483686 292816 483692
rect 292672 477488 292724 477494
rect 292672 477430 292724 477436
rect 293972 477358 294000 495037
rect 294064 495023 294446 495051
rect 294616 495023 294906 495051
rect 295382 495023 295472 495051
rect 294064 477426 294092 495023
rect 294616 489914 294644 495023
rect 295340 492720 295392 492726
rect 295340 492662 295392 492668
rect 294156 489886 294644 489914
rect 294156 479942 294184 489886
rect 295352 480078 295380 492662
rect 295444 480146 295472 495023
rect 295628 495023 295826 495051
rect 295904 495023 296194 495051
rect 296272 495023 296654 495051
rect 296824 495023 297114 495051
rect 297192 495023 297574 495051
rect 297744 495023 298034 495051
rect 298112 495023 298402 495051
rect 298480 495023 298862 495051
rect 299032 495023 299322 495051
rect 295524 492652 295576 492658
rect 295524 492594 295576 492600
rect 295432 480140 295484 480146
rect 295432 480082 295484 480088
rect 295340 480072 295392 480078
rect 295340 480014 295392 480020
rect 295536 480010 295564 492594
rect 295628 481166 295656 495023
rect 295904 492726 295932 495023
rect 295892 492720 295944 492726
rect 295892 492662 295944 492668
rect 296272 492658 296300 495023
rect 296260 492652 296312 492658
rect 296260 492594 296312 492600
rect 296720 492652 296772 492658
rect 296720 492594 296772 492600
rect 295616 481160 295668 481166
rect 295616 481102 295668 481108
rect 295524 480004 295576 480010
rect 295524 479946 295576 479952
rect 294144 479936 294196 479942
rect 294144 479878 294196 479884
rect 294052 477420 294104 477426
rect 294052 477362 294104 477368
rect 293960 477352 294012 477358
rect 293960 477294 294012 477300
rect 292578 476776 292634 476785
rect 292578 476711 292634 476720
rect 296732 463049 296760 492594
rect 296824 479874 296852 495023
rect 297192 489914 297220 495023
rect 297744 492658 297772 495023
rect 297732 492652 297784 492658
rect 297732 492594 297784 492600
rect 296916 489886 297220 489914
rect 296916 480214 296944 489886
rect 296904 480208 296956 480214
rect 296904 480150 296956 480156
rect 296812 479868 296864 479874
rect 296812 479810 296864 479816
rect 296718 463040 296774 463049
rect 296718 462975 296774 462984
rect 298112 460193 298140 495023
rect 298192 492652 298244 492658
rect 298192 492594 298244 492600
rect 298204 466342 298232 492594
rect 298480 489914 298508 495023
rect 299032 492658 299060 495023
rect 299020 492652 299072 492658
rect 299020 492594 299072 492600
rect 299860 489914 299888 495094
rect 298296 489886 298508 489914
rect 299492 489886 299888 489914
rect 298296 479806 298324 489886
rect 298284 479800 298336 479806
rect 298284 479742 298336 479748
rect 298192 466336 298244 466342
rect 298192 466278 298244 466284
rect 299492 460902 299520 489886
rect 307036 472666 307064 630634
rect 309796 568002 309824 647391
rect 311164 625184 311216 625190
rect 311164 625126 311216 625132
rect 309784 567996 309836 568002
rect 309784 567938 309836 567944
rect 311176 565282 311204 625126
rect 312556 572150 312584 648042
rect 313924 647896 313976 647902
rect 313924 647838 313976 647844
rect 312544 572144 312596 572150
rect 312544 572086 312596 572092
rect 313936 566574 313964 647838
rect 315304 647692 315356 647698
rect 315304 647634 315356 647640
rect 314016 647556 314068 647562
rect 314016 647498 314068 647504
rect 314028 566642 314056 647498
rect 315316 573578 315344 647634
rect 316696 582729 316724 684490
rect 318800 652044 318852 652050
rect 318800 651986 318852 651992
rect 318248 648168 318300 648174
rect 318248 648110 318300 648116
rect 316868 647828 316920 647834
rect 316868 647770 316920 647776
rect 316776 647420 316828 647426
rect 316776 647362 316828 647368
rect 316682 582720 316738 582729
rect 316682 582655 316738 582664
rect 315304 573572 315356 573578
rect 315304 573514 315356 573520
rect 314016 566636 314068 566642
rect 314016 566578 314068 566584
rect 313924 566568 313976 566574
rect 313924 566510 313976 566516
rect 311164 565276 311216 565282
rect 311164 565218 311216 565224
rect 315488 559904 315540 559910
rect 315488 559846 315540 559852
rect 312728 559496 312780 559502
rect 312728 559438 312780 559444
rect 309784 559428 309836 559434
rect 309784 559370 309836 559376
rect 309796 534070 309824 559370
rect 312544 559360 312596 559366
rect 312544 559302 312596 559308
rect 311164 558136 311216 558142
rect 311164 558078 311216 558084
rect 309784 534064 309836 534070
rect 309784 534006 309836 534012
rect 311176 532166 311204 558078
rect 311164 532160 311216 532166
rect 311164 532102 311216 532108
rect 312556 529922 312584 559302
rect 312636 557592 312688 557598
rect 312636 557534 312688 557540
rect 312648 531282 312676 557534
rect 312740 533798 312768 559438
rect 312820 559292 312872 559298
rect 312820 559234 312872 559240
rect 312832 535294 312860 559234
rect 315304 559224 315356 559230
rect 315304 559166 315356 559172
rect 312912 558952 312964 558958
rect 312912 558894 312964 558900
rect 312924 535430 312952 558894
rect 313096 555756 313148 555762
rect 313096 555698 313148 555704
rect 313004 555348 313056 555354
rect 313004 555290 313056 555296
rect 312912 535424 312964 535430
rect 312912 535366 312964 535372
rect 312820 535288 312872 535294
rect 312820 535230 312872 535236
rect 312728 533792 312780 533798
rect 312728 533734 312780 533740
rect 313016 532642 313044 555290
rect 313108 535362 313136 555698
rect 313096 535356 313148 535362
rect 313096 535298 313148 535304
rect 313004 532636 313056 532642
rect 313004 532578 313056 532584
rect 312636 531276 312688 531282
rect 312636 531218 312688 531224
rect 312544 529916 312596 529922
rect 312544 529858 312596 529864
rect 315316 529854 315344 559166
rect 315396 559088 315448 559094
rect 315396 559030 315448 559036
rect 315304 529848 315356 529854
rect 315304 529790 315356 529796
rect 315408 529786 315436 559030
rect 315500 531214 315528 559846
rect 316788 559774 316816 647362
rect 316880 561134 316908 647770
rect 318156 647488 318208 647494
rect 318156 647430 318208 647436
rect 318064 647352 318116 647358
rect 318064 647294 318116 647300
rect 317602 645280 317658 645289
rect 317602 645215 317658 645224
rect 317616 644502 317644 645215
rect 317604 644496 317656 644502
rect 317604 644438 317656 644444
rect 317694 640520 317750 640529
rect 317694 640455 317750 640464
rect 317708 640354 317736 640455
rect 317696 640348 317748 640354
rect 317696 640290 317748 640296
rect 317970 635760 318026 635769
rect 317970 635695 318026 635704
rect 317984 634846 318012 635695
rect 317972 634840 318024 634846
rect 317972 634782 318024 634788
rect 317418 631000 317474 631009
rect 317418 630935 317474 630944
rect 317432 630698 317460 630935
rect 317420 630692 317472 630698
rect 317420 630634 317472 630640
rect 317970 626240 318026 626249
rect 317970 626175 318026 626184
rect 317984 625190 318012 626175
rect 317972 625184 318024 625190
rect 317972 625126 318024 625132
rect 317970 621480 318026 621489
rect 317970 621415 318026 621424
rect 317984 621042 318012 621415
rect 317972 621036 318024 621042
rect 317972 620978 318024 620984
rect 317418 616720 317474 616729
rect 317418 616655 317474 616664
rect 317432 615534 317460 616655
rect 317420 615528 317472 615534
rect 317420 615470 317472 615476
rect 317970 611960 318026 611969
rect 317970 611895 318026 611904
rect 317984 611386 318012 611895
rect 317972 611380 318024 611386
rect 317972 611322 318024 611328
rect 317970 602440 318026 602449
rect 317970 602375 318026 602384
rect 317984 601730 318012 602375
rect 317972 601724 318024 601730
rect 317972 601666 318024 601672
rect 317970 597680 318026 597689
rect 317970 597615 318026 597624
rect 317984 597582 318012 597615
rect 317972 597576 318024 597582
rect 317972 597518 318024 597524
rect 317970 592920 318026 592929
rect 317970 592855 318026 592864
rect 317984 592074 318012 592855
rect 317972 592068 318024 592074
rect 317972 592010 318024 592016
rect 317420 586560 317472 586566
rect 317418 586528 317420 586537
rect 317472 586528 317474 586537
rect 317418 586463 317474 586472
rect 317510 577960 317566 577969
rect 317510 577895 317566 577904
rect 317524 570654 317552 577895
rect 317970 573200 318026 573209
rect 317970 573135 318026 573144
rect 317984 572762 318012 573135
rect 317972 572756 318024 572762
rect 317972 572698 318024 572704
rect 317512 570648 317564 570654
rect 317512 570590 317564 570596
rect 317970 568440 318026 568449
rect 317970 568375 318026 568384
rect 317984 567254 318012 568375
rect 317972 567248 318024 567254
rect 317972 567190 318024 567196
rect 317972 564392 318024 564398
rect 317972 564334 318024 564340
rect 317984 563689 318012 564334
rect 317970 563680 318026 563689
rect 317970 563615 318026 563624
rect 318076 562358 318104 647294
rect 318168 565214 318196 647430
rect 318260 575006 318288 648110
rect 318812 607209 318840 651986
rect 332600 648100 332652 648106
rect 332600 648042 332652 648048
rect 319720 647964 319772 647970
rect 319720 647906 319772 647912
rect 319534 647592 319590 647601
rect 319534 647527 319590 647536
rect 319444 646332 319496 646338
rect 319444 646274 319496 646280
rect 318798 607200 318854 607209
rect 318798 607135 318854 607144
rect 318248 575000 318300 575006
rect 318248 574942 318300 574948
rect 318156 565208 318208 565214
rect 318156 565150 318208 565156
rect 318064 562352 318116 562358
rect 318064 562294 318116 562300
rect 316868 561128 316920 561134
rect 316868 561070 316920 561076
rect 316776 559768 316828 559774
rect 316776 559710 316828 559716
rect 315580 559156 315632 559162
rect 315580 559098 315632 559104
rect 315592 535022 315620 559098
rect 318248 559020 318300 559026
rect 318248 558962 318300 558968
rect 317970 558920 318026 558929
rect 317970 558855 318026 558864
rect 316684 557864 316736 557870
rect 316684 557806 316736 557812
rect 315672 555688 315724 555694
rect 315672 555630 315724 555636
rect 315580 535016 315632 535022
rect 315580 534958 315632 534964
rect 315684 533730 315712 555630
rect 315672 533724 315724 533730
rect 315672 533666 315724 533672
rect 316696 531962 316724 557806
rect 317984 557734 318012 558855
rect 318064 558340 318116 558346
rect 318064 558282 318116 558288
rect 317972 557728 318024 557734
rect 317972 557670 318024 557676
rect 316868 556572 316920 556578
rect 316868 556514 316920 556520
rect 316776 556300 316828 556306
rect 316776 556242 316828 556248
rect 316788 533662 316816 556242
rect 316880 534954 316908 556514
rect 317972 554736 318024 554742
rect 317972 554678 318024 554684
rect 317984 554169 318012 554678
rect 317970 554160 318026 554169
rect 317970 554095 318026 554104
rect 317420 550588 317472 550594
rect 317420 550530 317472 550536
rect 317432 549409 317460 550530
rect 317418 549400 317474 549409
rect 317418 549335 317474 549344
rect 317972 545080 318024 545086
rect 317972 545022 318024 545028
rect 317984 544649 318012 545022
rect 317970 544640 318026 544649
rect 317970 544575 318026 544584
rect 316868 534948 316920 534954
rect 316868 534890 316920 534896
rect 316776 533656 316828 533662
rect 316776 533598 316828 533604
rect 316684 531956 316736 531962
rect 316684 531898 316736 531904
rect 318076 531758 318104 558282
rect 318156 557932 318208 557938
rect 318156 557874 318208 557880
rect 318168 532302 318196 557874
rect 318260 534750 318288 558962
rect 318616 557388 318668 557394
rect 318616 557330 318668 557336
rect 318338 556336 318394 556345
rect 318338 556271 318394 556280
rect 318248 534744 318300 534750
rect 318248 534686 318300 534692
rect 318352 534002 318380 556271
rect 318432 555144 318484 555150
rect 318432 555086 318484 555092
rect 318340 533996 318392 534002
rect 318340 533938 318392 533944
rect 318156 532296 318208 532302
rect 318156 532238 318208 532244
rect 318444 531894 318472 555086
rect 318522 554840 318578 554849
rect 318522 554775 318578 554784
rect 318536 532030 318564 554775
rect 318628 534886 318656 557330
rect 319352 557252 319404 557258
rect 319352 557194 319404 557200
rect 318708 555484 318760 555490
rect 318708 555426 318760 555432
rect 318720 539889 318748 555426
rect 319260 543040 319312 543046
rect 319260 542982 319312 542988
rect 318706 539880 318762 539889
rect 318706 539815 318762 539824
rect 319168 536308 319220 536314
rect 319168 536250 319220 536256
rect 318616 534880 318668 534886
rect 318616 534822 318668 534828
rect 319180 532098 319208 536250
rect 319272 532506 319300 542982
rect 319364 534818 319392 557194
rect 319456 556850 319484 646274
rect 319548 560998 319576 647527
rect 319628 647284 319680 647290
rect 319628 647226 319680 647232
rect 319640 562426 319668 647226
rect 319732 563718 319760 647906
rect 319812 647760 319864 647766
rect 319812 647702 319864 647708
rect 319824 572082 319852 647702
rect 323492 647284 323544 647290
rect 323492 647226 323544 647232
rect 323504 645946 323532 647226
rect 328090 646232 328146 646241
rect 328090 646167 328146 646176
rect 328104 645946 328132 646167
rect 332612 645946 332640 648042
rect 355140 647964 355192 647970
rect 355140 647906 355192 647912
rect 350540 647624 350592 647630
rect 350540 647566 350592 647572
rect 337108 647352 337160 647358
rect 337108 647294 337160 647300
rect 337120 645946 337148 647294
rect 341524 646672 341576 646678
rect 341524 646614 341576 646620
rect 341536 645946 341564 646614
rect 346582 646096 346638 646105
rect 346582 646031 346638 646040
rect 346596 645946 346624 646031
rect 323504 645918 323886 645946
rect 328104 645918 328394 645946
rect 332612 645918 332902 645946
rect 337120 645918 337410 645946
rect 341536 645918 341918 645946
rect 346426 645918 346624 645946
rect 350552 645946 350580 647566
rect 355152 645946 355180 647906
rect 375392 647902 375420 703582
rect 376312 703474 376340 703582
rect 376454 703520 376566 704960
rect 391818 703520 391930 704960
rect 407182 703520 407294 704960
rect 422546 703520 422658 704960
rect 437910 703520 438022 704960
rect 453274 703520 453386 704960
rect 468638 703520 468750 704960
rect 484002 703520 484114 704960
rect 498212 703582 499252 703610
rect 376496 703474 376524 703520
rect 376312 703446 376524 703474
rect 407224 701010 407252 703520
rect 407212 701004 407264 701010
rect 407212 700946 407264 700952
rect 437952 699718 437980 703520
rect 468680 701010 468708 703520
rect 468668 701004 468720 701010
rect 468668 700946 468720 700952
rect 436744 699712 436796 699718
rect 436744 699654 436796 699660
rect 437940 699712 437992 699718
rect 437940 699654 437992 699660
rect 400220 698964 400272 698970
rect 400220 698906 400272 698912
rect 400232 654134 400260 698906
rect 400232 654106 400720 654134
rect 378324 648032 378376 648038
rect 378324 647974 378376 647980
rect 359556 647896 359608 647902
rect 359556 647838 359608 647844
rect 375380 647896 375432 647902
rect 375380 647838 375432 647844
rect 359568 645946 359596 647838
rect 364340 647828 364392 647834
rect 364340 647770 364392 647776
rect 364352 645946 364380 647770
rect 373172 647760 373224 647766
rect 373172 647702 373224 647708
rect 368572 647692 368624 647698
rect 368572 647634 368624 647640
rect 368584 645946 368612 647634
rect 373184 645946 373212 647702
rect 378336 645946 378364 647974
rect 391938 647592 391994 647601
rect 382740 647556 382792 647562
rect 391938 647527 391994 647536
rect 382740 647498 382792 647504
rect 382752 645946 382780 647498
rect 387340 647488 387392 647494
rect 387340 647430 387392 647436
rect 387352 645946 387380 647430
rect 391952 645946 391980 647527
rect 396356 647420 396408 647426
rect 396356 647362 396408 647368
rect 396368 645946 396396 647362
rect 400692 645946 400720 654106
rect 429292 650684 429344 650690
rect 429292 650626 429344 650632
rect 427820 648168 427872 648174
rect 427820 648110 427872 648116
rect 423864 647896 423916 647902
rect 423864 647838 423916 647844
rect 418802 647456 418858 647465
rect 418802 647391 418858 647400
rect 409880 645992 409932 645998
rect 405370 645960 405426 645969
rect 350552 645918 350934 645946
rect 355152 645918 355442 645946
rect 359568 645918 359950 645946
rect 364352 645918 364458 645946
rect 368584 645918 368966 645946
rect 373184 645918 373474 645946
rect 378336 645918 378626 645946
rect 382752 645918 383134 645946
rect 387352 645918 387642 645946
rect 391952 645918 392150 645946
rect 396368 645918 396658 645946
rect 400692 645918 401166 645946
rect 405426 645918 405674 645946
rect 418816 645946 418844 647391
rect 409932 645940 410182 645946
rect 409880 645934 410182 645940
rect 409892 645918 410182 645934
rect 414400 645930 414690 645946
rect 414388 645924 414690 645930
rect 405370 645895 405426 645904
rect 414440 645918 414690 645924
rect 418816 645918 419198 645946
rect 414388 645866 414440 645872
rect 423876 645810 423904 647838
rect 427832 645946 427860 648110
rect 428464 646468 428516 646474
rect 428464 646410 428516 646416
rect 427832 645918 428214 645946
rect 423706 645782 423904 645810
rect 428476 634778 428504 646410
rect 428464 634772 428516 634778
rect 428464 634714 428516 634720
rect 429198 598360 429254 598369
rect 429198 598295 429254 598304
rect 428370 573336 428426 573345
rect 428370 573271 428426 573280
rect 319812 572076 319864 572082
rect 319812 572018 319864 572024
rect 319812 569220 319864 569226
rect 319812 569162 319864 569168
rect 319720 563712 319772 563718
rect 319720 563654 319772 563660
rect 319628 562420 319680 562426
rect 319628 562362 319680 562368
rect 319536 560992 319588 560998
rect 319536 560934 319588 560940
rect 319628 557796 319680 557802
rect 319628 557738 319680 557744
rect 319536 557660 319588 557666
rect 319536 557602 319588 557608
rect 319444 556844 319496 556850
rect 319444 556786 319496 556792
rect 319444 555076 319496 555082
rect 319444 555018 319496 555024
rect 319456 543046 319484 555018
rect 319444 543040 319496 543046
rect 319444 542982 319496 542988
rect 319548 536314 319576 557602
rect 319536 536308 319588 536314
rect 319536 536250 319588 536256
rect 319640 536194 319668 557738
rect 319720 556640 319772 556646
rect 319720 556582 319772 556588
rect 319456 536166 319668 536194
rect 319352 534812 319404 534818
rect 319352 534754 319404 534760
rect 319456 532574 319484 536166
rect 319732 536058 319760 556582
rect 319548 536030 319760 536058
rect 319548 533934 319576 536030
rect 319824 535378 319852 569162
rect 319902 556200 319958 556209
rect 319902 556135 319958 556144
rect 319916 535401 319944 556135
rect 319640 535350 319852 535378
rect 319902 535392 319958 535401
rect 319640 535106 319668 535350
rect 319902 535327 319958 535336
rect 356086 535214 356284 535242
rect 319640 535078 319760 535106
rect 319536 533928 319588 533934
rect 319536 533870 319588 533876
rect 319732 532681 319760 535078
rect 319916 535078 320022 535106
rect 324530 535078 324912 535106
rect 319718 532672 319774 532681
rect 319628 532636 319680 532642
rect 319916 532658 319944 535078
rect 324884 534041 324912 535078
rect 328656 535078 329038 535106
rect 333256 535078 333546 535106
rect 337672 535078 338054 535106
rect 342272 535078 342562 535106
rect 346688 535078 347070 535106
rect 351288 535078 351578 535106
rect 324870 534032 324926 534041
rect 324870 533967 324926 533976
rect 328656 533186 328684 535078
rect 328644 533180 328696 533186
rect 328644 533122 328696 533128
rect 319718 532607 319774 532616
rect 319824 532630 319944 532658
rect 319628 532578 319680 532584
rect 319444 532568 319496 532574
rect 319444 532510 319496 532516
rect 319640 532522 319668 532578
rect 319824 532522 319852 532630
rect 333256 532574 333284 535078
rect 337672 532681 337700 535078
rect 342272 532710 342300 535078
rect 342260 532704 342312 532710
rect 337658 532672 337714 532681
rect 342260 532646 342312 532652
rect 346688 532642 346716 535078
rect 351288 534206 351316 535078
rect 351276 534200 351328 534206
rect 351276 534142 351328 534148
rect 337658 532607 337714 532616
rect 346676 532636 346728 532642
rect 346676 532578 346728 532584
rect 319260 532500 319312 532506
rect 319640 532494 319852 532522
rect 333244 532568 333296 532574
rect 333244 532510 333296 532516
rect 319904 532500 319956 532506
rect 319260 532442 319312 532448
rect 319904 532442 319956 532448
rect 319168 532092 319220 532098
rect 319168 532034 319220 532040
rect 318524 532024 318576 532030
rect 318524 531966 318576 531972
rect 319916 531962 319944 532442
rect 356256 532030 356284 535214
rect 360304 535078 360594 535106
rect 364720 535078 365102 535106
rect 369320 535078 369610 535106
rect 374472 535078 374762 535106
rect 378152 535078 379270 535106
rect 383672 535078 383778 535106
rect 387904 535078 388286 535106
rect 391952 535078 392794 535106
rect 396920 535078 397302 535106
rect 401612 535078 401810 535106
rect 405936 535078 406318 535106
rect 410536 535078 410826 535106
rect 414952 535078 415334 535106
rect 419552 535078 419842 535106
rect 423968 535078 424350 535106
rect 360304 532098 360332 535078
rect 364720 532166 364748 535078
rect 369320 534138 369348 535078
rect 369308 534132 369360 534138
rect 369308 534074 369360 534080
rect 374472 532234 374500 535078
rect 374460 532228 374512 532234
rect 374460 532170 374512 532176
rect 364708 532160 364760 532166
rect 364708 532102 364760 532108
rect 360292 532092 360344 532098
rect 360292 532034 360344 532040
rect 356244 532024 356296 532030
rect 356244 531966 356296 531972
rect 319904 531956 319956 531962
rect 319904 531898 319956 531904
rect 319996 531956 320048 531962
rect 319996 531898 320048 531904
rect 318432 531888 318484 531894
rect 318432 531830 318484 531836
rect 320008 531758 320036 531898
rect 318064 531752 318116 531758
rect 318064 531694 318116 531700
rect 319996 531752 320048 531758
rect 319996 531694 320048 531700
rect 315488 531208 315540 531214
rect 315488 531150 315540 531156
rect 315396 529780 315448 529786
rect 315396 529722 315448 529728
rect 356796 492584 356848 492590
rect 356796 492526 356848 492532
rect 356704 492176 356756 492182
rect 356704 492118 356756 492124
rect 307024 472660 307076 472666
rect 307024 472602 307076 472608
rect 339684 461712 339736 461718
rect 339684 461654 339736 461660
rect 339696 461281 339724 461654
rect 339682 461272 339738 461281
rect 339682 461207 339738 461216
rect 339696 461106 339724 461207
rect 339684 461100 339736 461106
rect 339684 461042 339736 461048
rect 338304 461032 338356 461038
rect 338302 461000 338304 461009
rect 338356 461000 338358 461009
rect 338302 460935 338358 460944
rect 350998 461000 351054 461009
rect 350998 460935 351000 460944
rect 351052 460935 351054 460944
rect 351000 460906 351052 460912
rect 299480 460896 299532 460902
rect 299480 460838 299532 460844
rect 298098 460184 298154 460193
rect 298098 460119 298154 460128
rect 291200 459468 291252 459474
rect 291200 459410 291252 459416
rect 288440 459332 288492 459338
rect 288440 459274 288492 459280
rect 274640 459264 274692 459270
rect 274640 459206 274692 459212
rect 273260 459128 273312 459134
rect 273260 459070 273312 459076
rect 264980 459060 265032 459066
rect 264980 459002 265032 459008
rect 253940 458992 253992 458998
rect 253940 458934 253992 458940
rect 247040 458924 247092 458930
rect 247040 458866 247092 458872
rect 245660 458856 245712 458862
rect 245660 458798 245712 458804
rect 263690 375048 263746 375057
rect 263690 374983 263746 374992
rect 311806 375048 311862 375057
rect 311806 374983 311862 374992
rect 244278 374504 244334 374513
rect 244278 374439 244280 374448
rect 244332 374439 244334 374448
rect 248694 374504 248750 374513
rect 248694 374439 248750 374448
rect 250074 374504 250130 374513
rect 250074 374439 250130 374448
rect 244280 374410 244332 374416
rect 248708 374406 248736 374439
rect 241244 374400 241296 374406
rect 241244 374342 241296 374348
rect 248696 374400 248748 374406
rect 248696 374342 248748 374348
rect 241152 374332 241204 374338
rect 241152 374274 241204 374280
rect 222016 374128 222068 374134
rect 222016 374070 222068 374076
rect 220728 372836 220780 372842
rect 220728 372778 220780 372784
rect 220740 372638 220768 372778
rect 220912 372768 220964 372774
rect 220832 372728 220912 372756
rect 220728 372632 220780 372638
rect 220728 372574 220780 372580
rect 220832 372450 220860 372728
rect 220912 372710 220964 372716
rect 220740 372422 220860 372450
rect 220544 372224 220596 372230
rect 220544 372166 220596 372172
rect 220452 372156 220504 372162
rect 220452 372098 220504 372104
rect 220464 371958 220492 372098
rect 220452 371952 220504 371958
rect 220452 371894 220504 371900
rect 220556 371686 220584 372166
rect 220636 372020 220688 372026
rect 220636 371962 220688 371968
rect 220544 371680 220596 371686
rect 220544 371622 220596 371628
rect 220648 371550 220676 371962
rect 220636 371544 220688 371550
rect 220636 371486 220688 371492
rect 220740 371113 220768 372422
rect 220820 372088 220872 372094
rect 220820 372030 220872 372036
rect 221924 372088 221976 372094
rect 221924 372030 221976 372036
rect 220726 371104 220782 371113
rect 220726 371039 220782 371048
rect 220832 350538 220860 372030
rect 221936 371550 221964 372030
rect 221924 371544 221976 371550
rect 220910 371512 220966 371521
rect 221924 371486 221976 371492
rect 220910 371447 220966 371456
rect 220820 350532 220872 350538
rect 220820 350474 220872 350480
rect 220924 349246 220952 371447
rect 222028 371385 222056 374070
rect 236458 373688 236514 373697
rect 236458 373623 236514 373632
rect 236472 373590 236500 373623
rect 236460 373584 236512 373590
rect 236460 373526 236512 373532
rect 224224 373516 224276 373522
rect 224224 373458 224276 373464
rect 222106 372056 222162 372065
rect 222106 371991 222162 372000
rect 222120 371521 222148 371991
rect 224236 371890 224264 373458
rect 238114 372600 238170 372609
rect 238114 372535 238170 372544
rect 239126 372600 239182 372609
rect 239126 372535 239182 372544
rect 224224 371884 224276 371890
rect 224224 371826 224276 371832
rect 222106 371512 222162 371521
rect 222106 371447 222162 371456
rect 238128 371414 238156 372535
rect 239140 371822 239168 372535
rect 241164 371958 241192 374274
rect 241256 372026 241284 374342
rect 250088 374338 250116 374439
rect 250076 374332 250128 374338
rect 250076 374274 250128 374280
rect 263704 374270 263732 374983
rect 281448 374808 281500 374814
rect 281448 374750 281500 374756
rect 271142 374504 271198 374513
rect 271142 374439 271198 374448
rect 275834 374504 275890 374513
rect 275834 374439 275890 374448
rect 263692 374264 263744 374270
rect 263692 374206 263744 374212
rect 271156 374202 271184 374439
rect 271144 374196 271196 374202
rect 271144 374138 271196 374144
rect 275848 374134 275876 374439
rect 270316 374128 270368 374134
rect 270316 374070 270368 374076
rect 275836 374128 275888 374134
rect 275836 374070 275888 374076
rect 258078 373960 258134 373969
rect 258078 373895 258134 373904
rect 242898 373688 242954 373697
rect 242898 373623 242954 373632
rect 242912 373454 242940 373623
rect 242900 373448 242952 373454
rect 242900 373390 242952 373396
rect 253938 373280 253994 373289
rect 253938 373215 253940 373224
rect 253992 373215 253994 373224
rect 255410 373280 255466 373289
rect 255410 373215 255466 373224
rect 256698 373280 256754 373289
rect 256698 373215 256754 373224
rect 253940 373186 253992 373192
rect 255424 373182 255452 373215
rect 255412 373176 255464 373182
rect 247130 373144 247186 373153
rect 255412 373118 255464 373124
rect 247130 373079 247186 373088
rect 244278 372600 244334 372609
rect 244278 372535 244334 372544
rect 244292 372298 244320 372535
rect 244280 372292 244332 372298
rect 244280 372234 244332 372240
rect 241244 372020 241296 372026
rect 241244 371962 241296 371968
rect 241152 371952 241204 371958
rect 241152 371894 241204 371900
rect 245658 371920 245714 371929
rect 245658 371855 245714 371864
rect 246026 371920 246082 371929
rect 247144 371890 247172 373079
rect 256712 373046 256740 373215
rect 258092 373114 258120 373895
rect 269210 373416 269266 373425
rect 269210 373351 269266 373360
rect 269224 373318 269252 373351
rect 269212 373312 269264 373318
rect 269212 373254 269264 373260
rect 261298 373144 261354 373153
rect 258080 373108 258132 373114
rect 261298 373079 261354 373088
rect 264978 373144 265034 373153
rect 264978 373079 265034 373088
rect 258080 373050 258132 373056
rect 256700 373040 256752 373046
rect 256700 372982 256752 372988
rect 259644 372972 259696 372978
rect 259644 372914 259696 372920
rect 259460 372904 259512 372910
rect 259460 372846 259512 372852
rect 259472 372609 259500 372846
rect 259656 372609 259684 372914
rect 261312 372706 261340 373079
rect 264992 372842 265020 373079
rect 264980 372836 265032 372842
rect 264980 372778 265032 372784
rect 266360 372768 266412 372774
rect 266360 372710 266412 372716
rect 261300 372700 261352 372706
rect 261300 372642 261352 372648
rect 262220 372632 262272 372638
rect 251178 372600 251234 372609
rect 251178 372535 251234 372544
rect 252558 372600 252614 372609
rect 252558 372535 252614 372544
rect 259458 372600 259514 372609
rect 259458 372535 259514 372544
rect 259642 372600 259698 372609
rect 259642 372535 259698 372544
rect 262218 372600 262220 372609
rect 266372 372609 266400 372710
rect 262272 372600 262274 372609
rect 262218 372535 262274 372544
rect 266358 372600 266414 372609
rect 266358 372535 266414 372544
rect 251192 372230 251220 372535
rect 251180 372224 251232 372230
rect 251180 372166 251232 372172
rect 246026 371855 246082 371864
rect 247132 371884 247184 371890
rect 239128 371816 239180 371822
rect 239128 371758 239180 371764
rect 240048 371816 240100 371822
rect 240048 371758 240100 371764
rect 240060 371414 240088 371758
rect 245672 371754 245700 371855
rect 245660 371748 245712 371754
rect 245660 371690 245712 371696
rect 246040 371657 246068 371855
rect 247132 371826 247184 371832
rect 251180 371680 251232 371686
rect 246026 371648 246082 371657
rect 246026 371583 246082 371592
rect 251178 371648 251180 371657
rect 251232 371648 251234 371657
rect 251178 371583 251234 371592
rect 252572 371550 252600 372535
rect 258170 371648 258226 371657
rect 258170 371583 258226 371592
rect 252560 371544 252612 371550
rect 247038 371512 247094 371521
rect 247038 371447 247094 371456
rect 249798 371512 249854 371521
rect 252560 371486 252612 371492
rect 252650 371512 252706 371521
rect 249798 371447 249854 371456
rect 252650 371447 252706 371456
rect 255318 371512 255374 371521
rect 255318 371447 255374 371456
rect 238116 371408 238168 371414
rect 222014 371376 222070 371385
rect 238116 371350 238168 371356
rect 240048 371408 240100 371414
rect 240048 371350 240100 371356
rect 222014 371311 222070 371320
rect 247052 369034 247080 371447
rect 249812 369238 249840 371447
rect 249800 369232 249852 369238
rect 249800 369174 249852 369180
rect 247040 369028 247092 369034
rect 247040 368970 247092 368976
rect 252664 368966 252692 371447
rect 255332 369102 255360 371447
rect 258184 369442 258212 371583
rect 260838 371512 260894 371521
rect 260838 371447 260894 371456
rect 263598 371512 263654 371521
rect 263598 371447 263654 371456
rect 264978 371512 265034 371521
rect 264978 371447 265034 371456
rect 267738 371512 267794 371521
rect 267738 371447 267794 371456
rect 258172 369436 258224 369442
rect 258172 369378 258224 369384
rect 260852 369170 260880 371447
rect 263612 369306 263640 371447
rect 264992 370326 265020 371447
rect 264980 370320 265032 370326
rect 264980 370262 265032 370268
rect 267752 369510 267780 371447
rect 270328 371385 270356 374070
rect 275848 372638 275876 374070
rect 275836 372632 275888 372638
rect 271878 372600 271934 372609
rect 271878 372535 271934 372544
rect 273258 372600 273314 372609
rect 275836 372574 275888 372580
rect 281460 372570 281488 374750
rect 311820 374746 311848 374983
rect 314566 374776 314622 374785
rect 311808 374740 311860 374746
rect 314566 374711 314622 374720
rect 311808 374682 311860 374688
rect 314580 374678 314608 374711
rect 314568 374672 314620 374678
rect 314568 374614 314620 374620
rect 320914 374504 320970 374513
rect 320914 374439 320970 374448
rect 320928 374066 320956 374439
rect 320916 374060 320968 374066
rect 320916 374002 320968 374008
rect 300858 373144 300914 373153
rect 300858 373079 300914 373088
rect 273258 372535 273260 372544
rect 271892 372502 271920 372535
rect 273312 372535 273314 372544
rect 281448 372564 281500 372570
rect 273260 372506 273312 372512
rect 281448 372506 281500 372512
rect 271880 372496 271932 372502
rect 271880 372438 271932 372444
rect 280066 372464 280122 372473
rect 280066 372399 280122 372408
rect 276018 371784 276074 371793
rect 276018 371719 276074 371728
rect 274640 371680 274692 371686
rect 274640 371622 274692 371628
rect 270314 371376 270370 371385
rect 270314 371311 270370 371320
rect 270498 371376 270554 371385
rect 270498 371311 270554 371320
rect 273258 371376 273314 371385
rect 273258 371311 273314 371320
rect 270512 370462 270540 371311
rect 270500 370456 270552 370462
rect 270500 370398 270552 370404
rect 267740 369504 267792 369510
rect 267740 369446 267792 369452
rect 273272 369374 273300 371311
rect 274652 370530 274680 371622
rect 276032 371550 276060 371719
rect 280080 371618 280108 372399
rect 292578 372192 292634 372201
rect 292578 372127 292634 372136
rect 280068 371612 280120 371618
rect 280068 371554 280120 371560
rect 276020 371544 276072 371550
rect 276020 371486 276072 371492
rect 277306 371512 277362 371521
rect 277306 371447 277362 371456
rect 276018 371376 276074 371385
rect 276018 371311 276074 371320
rect 274640 370524 274692 370530
rect 274640 370466 274692 370472
rect 276032 370394 276060 371311
rect 276020 370388 276072 370394
rect 276020 370330 276072 370336
rect 273260 369368 273312 369374
rect 273260 369310 273312 369316
rect 263600 369300 263652 369306
rect 263600 369242 263652 369248
rect 260840 369164 260892 369170
rect 260840 369106 260892 369112
rect 255320 369096 255372 369102
rect 255320 369038 255372 369044
rect 252652 368960 252704 368966
rect 252652 368902 252704 368908
rect 277320 349858 277348 371447
rect 277398 371376 277454 371385
rect 277398 371311 277454 371320
rect 280158 371376 280214 371385
rect 280158 371311 280214 371320
rect 282918 371376 282974 371385
rect 282918 371311 282974 371320
rect 285678 371376 285734 371385
rect 285678 371311 285734 371320
rect 287242 371376 287298 371385
rect 287242 371311 287298 371320
rect 289818 371376 289874 371385
rect 289818 371311 289874 371320
rect 277412 370598 277440 371311
rect 277400 370592 277452 370598
rect 277400 370534 277452 370540
rect 280172 369646 280200 371311
rect 280160 369640 280212 369646
rect 280160 369582 280212 369588
rect 282932 369578 282960 371311
rect 285692 370666 285720 371311
rect 287256 371006 287284 371311
rect 287244 371000 287296 371006
rect 287244 370942 287296 370948
rect 289832 370734 289860 371311
rect 292592 370802 292620 372127
rect 295338 371376 295394 371385
rect 295338 371311 295394 371320
rect 298098 371376 298154 371385
rect 298098 371311 298154 371320
rect 295352 370870 295380 371311
rect 298112 371142 298140 371311
rect 298100 371136 298152 371142
rect 298100 371078 298152 371084
rect 300872 370938 300900 373079
rect 356612 372632 356664 372638
rect 326066 372600 326122 372609
rect 356612 372574 356664 372580
rect 326066 372535 326068 372544
rect 326120 372535 326122 372544
rect 326068 372506 326120 372512
rect 343178 372192 343234 372201
rect 343178 372127 343234 372136
rect 343454 372192 343510 372201
rect 343454 372127 343510 372136
rect 302238 371784 302294 371793
rect 302238 371719 302294 371728
rect 302252 371686 302280 371719
rect 302240 371680 302292 371686
rect 302240 371622 302292 371628
rect 304998 371376 305054 371385
rect 304998 371311 305054 371320
rect 307758 371376 307814 371385
rect 307758 371311 307814 371320
rect 310518 371376 310574 371385
rect 310518 371311 310574 371320
rect 313278 371376 313334 371385
rect 313278 371311 313334 371320
rect 322938 371376 322994 371385
rect 343192 371346 343220 372127
rect 322938 371311 322994 371320
rect 343180 371340 343232 371346
rect 305012 371210 305040 371311
rect 305000 371204 305052 371210
rect 305000 371146 305052 371152
rect 307772 371074 307800 371311
rect 307760 371068 307812 371074
rect 307760 371010 307812 371016
rect 300860 370932 300912 370938
rect 300860 370874 300912 370880
rect 295340 370864 295392 370870
rect 295340 370806 295392 370812
rect 292580 370796 292632 370802
rect 292580 370738 292632 370744
rect 289820 370728 289872 370734
rect 289820 370670 289872 370676
rect 285680 370660 285732 370666
rect 285680 370602 285732 370608
rect 310532 369714 310560 371311
rect 313292 369782 313320 371311
rect 322952 369850 322980 371311
rect 343180 371282 343232 371288
rect 343468 371278 343496 372127
rect 343456 371272 343508 371278
rect 343456 371214 343508 371220
rect 322940 369844 322992 369850
rect 322940 369786 322992 369792
rect 313280 369776 313332 369782
rect 313280 369718 313332 369724
rect 310520 369708 310572 369714
rect 310520 369650 310572 369656
rect 282920 369572 282972 369578
rect 282920 369514 282972 369520
rect 338488 351348 338540 351354
rect 338488 351290 338540 351296
rect 338500 350577 338528 351290
rect 340512 351280 340564 351286
rect 340512 351222 340564 351228
rect 340524 350577 340552 351222
rect 351644 351212 351696 351218
rect 351644 351154 351696 351160
rect 351656 350577 351684 351154
rect 338486 350568 338542 350577
rect 338486 350503 338542 350512
rect 340510 350568 340566 350577
rect 340510 350503 340566 350512
rect 351642 350568 351698 350577
rect 351642 350503 351698 350512
rect 277308 349852 277360 349858
rect 277308 349794 277360 349800
rect 220912 349240 220964 349246
rect 220912 349182 220964 349188
rect 250442 265024 250498 265033
rect 250442 264959 250498 264968
rect 274178 265024 274234 265033
rect 274178 264959 274234 264968
rect 221188 264920 221240 264926
rect 221188 264862 221240 264868
rect 221096 264852 221148 264858
rect 221096 264794 221148 264800
rect 221004 264784 221056 264790
rect 221004 264726 221056 264732
rect 220912 264648 220964 264654
rect 220912 264590 220964 264596
rect 220820 264104 220872 264110
rect 220820 264046 220872 264052
rect 220268 241256 220320 241262
rect 220268 241198 220320 241204
rect 220084 241120 220136 241126
rect 220084 241062 220136 241068
rect 220096 240281 220124 241062
rect 220280 240310 220308 241198
rect 220636 241188 220688 241194
rect 220636 241130 220688 241136
rect 220268 240304 220320 240310
rect 220082 240272 220138 240281
rect 220268 240246 220320 240252
rect 220648 240242 220676 241130
rect 220728 241052 220780 241058
rect 220728 240994 220780 241000
rect 220740 240446 220768 240994
rect 220728 240440 220780 240446
rect 220728 240382 220780 240388
rect 220082 240207 220138 240216
rect 220636 240236 220688 240242
rect 220636 240178 220688 240184
rect 220832 239902 220860 264046
rect 220820 239896 220872 239902
rect 220820 239838 220872 239844
rect 220728 239828 220780 239834
rect 220728 239770 220780 239776
rect 220740 239714 220768 239770
rect 220740 239686 220860 239714
rect 220924 239698 220952 264590
rect 220832 239578 220860 239686
rect 220912 239692 220964 239698
rect 220912 239634 220964 239640
rect 221016 239578 221044 264726
rect 221108 240106 221136 264794
rect 221200 241398 221228 264862
rect 250456 264722 250484 264959
rect 250444 264716 250496 264722
rect 250444 264658 250496 264664
rect 274192 264654 274220 264959
rect 224224 264648 224276 264654
rect 224224 264590 224276 264596
rect 274180 264648 274232 264654
rect 274180 264590 274232 264596
rect 291842 264616 291898 264625
rect 224236 264178 224264 264590
rect 280804 264580 280856 264586
rect 291842 264551 291898 264560
rect 293406 264616 293462 264625
rect 293406 264551 293462 264560
rect 280804 264522 280856 264528
rect 280816 264353 280844 264522
rect 285956 264512 286008 264518
rect 285956 264454 286008 264460
rect 283380 264444 283432 264450
rect 283380 264386 283432 264392
rect 283392 264353 283420 264386
rect 285968 264353 285996 264454
rect 290924 264376 290976 264382
rect 280802 264344 280858 264353
rect 280802 264279 280858 264288
rect 283378 264344 283434 264353
rect 283378 264279 283434 264288
rect 285954 264344 286010 264353
rect 285954 264279 286010 264288
rect 288162 264344 288218 264353
rect 288162 264279 288164 264288
rect 288216 264279 288218 264288
rect 290922 264344 290924 264353
rect 291856 264353 291884 264551
rect 290976 264344 290978 264353
rect 290922 264279 290978 264288
rect 291842 264344 291898 264353
rect 291842 264279 291898 264288
rect 288164 264250 288216 264256
rect 293420 264246 293448 264551
rect 293408 264240 293460 264246
rect 293408 264182 293460 264188
rect 224224 264172 224276 264178
rect 224224 264114 224276 264120
rect 273260 263628 273312 263634
rect 273260 263570 273312 263576
rect 279240 263628 279292 263634
rect 279240 263570 279292 263576
rect 273272 263537 273300 263570
rect 279252 263537 279280 263570
rect 308404 263560 308456 263566
rect 235998 263528 236054 263537
rect 235998 263463 236054 263472
rect 238758 263528 238814 263537
rect 238758 263463 238814 263472
rect 243082 263528 243138 263537
rect 243082 263463 243138 263472
rect 247130 263528 247186 263537
rect 247130 263463 247186 263472
rect 247682 263528 247738 263537
rect 247682 263463 247738 263472
rect 253570 263528 253626 263537
rect 253570 263463 253626 263472
rect 256146 263528 256202 263537
rect 256146 263463 256202 263472
rect 258170 263528 258226 263537
rect 258170 263463 258226 263472
rect 260838 263528 260894 263537
rect 260838 263463 260894 263472
rect 262218 263528 262274 263537
rect 262218 263463 262274 263472
rect 263598 263528 263654 263537
rect 263598 263463 263654 263472
rect 264978 263528 265034 263537
rect 264978 263463 265034 263472
rect 265898 263528 265954 263537
rect 265898 263463 265954 263472
rect 268290 263528 268346 263537
rect 268290 263463 268346 263472
rect 269762 263528 269818 263537
rect 269762 263463 269818 263472
rect 270866 263528 270922 263537
rect 270866 263463 270922 263472
rect 271234 263528 271290 263537
rect 271234 263463 271290 263472
rect 272062 263528 272118 263537
rect 272062 263463 272118 263472
rect 273258 263528 273314 263537
rect 273258 263463 273314 263472
rect 275926 263528 275982 263537
rect 275926 263463 275982 263472
rect 276110 263528 276166 263537
rect 276110 263463 276166 263472
rect 279238 263528 279294 263537
rect 279238 263463 279294 263472
rect 305826 263528 305882 263537
rect 305826 263463 305828 263472
rect 236012 260166 236040 263463
rect 237378 262304 237434 262313
rect 237378 262239 237434 262248
rect 236000 260160 236052 260166
rect 236000 260102 236052 260108
rect 221188 241392 221240 241398
rect 221188 241334 221240 241340
rect 237392 240990 237420 262239
rect 237380 240984 237432 240990
rect 237380 240926 237432 240932
rect 238772 240650 238800 263463
rect 240138 262304 240194 262313
rect 240138 262239 240194 262248
rect 241518 262304 241574 262313
rect 241518 262239 241574 262248
rect 240152 241466 240180 262239
rect 240140 241460 240192 241466
rect 240140 241402 240192 241408
rect 241532 240786 241560 262239
rect 243096 260778 243124 263463
rect 244370 262984 244426 262993
rect 244370 262919 244426 262928
rect 244278 262304 244334 262313
rect 244278 262239 244334 262248
rect 243084 260772 243136 260778
rect 243084 260714 243136 260720
rect 244292 240854 244320 262239
rect 244384 260846 244412 262919
rect 245658 262304 245714 262313
rect 245658 262239 245714 262248
rect 244372 260840 244424 260846
rect 244372 260782 244424 260788
rect 245672 240922 245700 262239
rect 247144 241330 247172 263463
rect 247696 262750 247724 263463
rect 253584 262886 253612 263463
rect 256160 263158 256188 263463
rect 256148 263152 256200 263158
rect 256148 263094 256200 263100
rect 253572 262880 253624 262886
rect 253572 262822 253624 262828
rect 247684 262744 247736 262750
rect 247684 262686 247736 262692
rect 251178 262440 251234 262449
rect 251178 262375 251234 262384
rect 248418 262304 248474 262313
rect 248418 262239 248474 262248
rect 249798 262304 249854 262313
rect 249798 262239 249854 262248
rect 247132 241324 247184 241330
rect 247132 241266 247184 241272
rect 248432 241058 248460 262239
rect 249812 241126 249840 262239
rect 251192 241262 251220 262375
rect 251270 262304 251326 262313
rect 251270 262239 251326 262248
rect 252650 262304 252706 262313
rect 252650 262239 252706 262248
rect 253938 262304 253994 262313
rect 253938 262239 253994 262248
rect 255318 262304 255374 262313
rect 255318 262239 255374 262248
rect 256698 262304 256754 262313
rect 256698 262239 256754 262248
rect 251180 241256 251232 241262
rect 251180 241198 251232 241204
rect 251284 241194 251312 262239
rect 251272 241188 251324 241194
rect 251272 241130 251324 241136
rect 249800 241120 249852 241126
rect 249800 241062 249852 241068
rect 248420 241052 248472 241058
rect 248420 240994 248472 241000
rect 245660 240916 245712 240922
rect 245660 240858 245712 240864
rect 244280 240848 244332 240854
rect 244280 240790 244332 240796
rect 241520 240780 241572 240786
rect 241520 240722 241572 240728
rect 252664 240718 252692 262239
rect 253952 241398 253980 262239
rect 253940 241392 253992 241398
rect 253940 241334 253992 241340
rect 252652 240712 252704 240718
rect 252652 240654 252704 240660
rect 238760 240644 238812 240650
rect 238760 240586 238812 240592
rect 221096 240100 221148 240106
rect 221096 240042 221148 240048
rect 222108 240100 222160 240106
rect 222108 240042 222160 240048
rect 221108 239902 221136 240042
rect 221096 239896 221148 239902
rect 221096 239838 221148 239844
rect 222120 239834 222148 240042
rect 222108 239828 222160 239834
rect 222108 239770 222160 239776
rect 222200 239828 222252 239834
rect 222200 239770 222252 239776
rect 222212 239714 222240 239770
rect 220832 239550 221044 239578
rect 222120 239686 222240 239714
rect 220832 239290 220860 239550
rect 222120 239290 222148 239686
rect 255332 239358 255360 262239
rect 256712 239562 256740 262239
rect 258184 239630 258212 263463
rect 258354 262984 258410 262993
rect 258354 262919 258410 262928
rect 258368 262818 258396 262919
rect 258356 262812 258408 262818
rect 258356 262754 258408 262760
rect 259550 262440 259606 262449
rect 259550 262375 259606 262384
rect 259458 262304 259514 262313
rect 259458 262239 259514 262248
rect 258172 239624 258224 239630
rect 258172 239566 258224 239572
rect 256700 239556 256752 239562
rect 256700 239498 256752 239504
rect 259472 239494 259500 262239
rect 259564 239766 259592 262375
rect 259552 239760 259604 239766
rect 259552 239702 259604 239708
rect 259460 239488 259512 239494
rect 259460 239430 259512 239436
rect 260852 239426 260880 263463
rect 260932 263084 260984 263090
rect 260932 263026 260984 263032
rect 260944 262993 260972 263026
rect 260930 262984 260986 262993
rect 260930 262919 260986 262928
rect 262232 239970 262260 263463
rect 263612 262954 263640 263463
rect 263600 262948 263652 262954
rect 263600 262890 263652 262896
rect 263598 262304 263654 262313
rect 263598 262239 263654 262248
rect 262220 239964 262272 239970
rect 262220 239906 262272 239912
rect 263612 239698 263640 262239
rect 264992 240038 265020 263463
rect 265912 263226 265940 263463
rect 268304 263430 268332 263463
rect 268292 263424 268344 263430
rect 268292 263366 268344 263372
rect 265900 263220 265952 263226
rect 265900 263162 265952 263168
rect 266358 262440 266414 262449
rect 266358 262375 266414 262384
rect 264980 240032 265032 240038
rect 264980 239974 265032 239980
rect 266372 239834 266400 262375
rect 266450 262304 266506 262313
rect 266450 262239 266506 262248
rect 267738 262304 267794 262313
rect 267738 262239 267794 262248
rect 266464 239902 266492 262239
rect 267752 240106 267780 262239
rect 269776 261594 269804 263463
rect 270880 263294 270908 263463
rect 270868 263288 270920 263294
rect 270868 263230 270920 263236
rect 269764 261588 269816 261594
rect 269764 261530 269816 261536
rect 271248 261526 271276 263463
rect 272076 262274 272104 263463
rect 273352 263016 273404 263022
rect 273350 262984 273352 262993
rect 273404 262984 273406 262993
rect 273350 262919 273406 262928
rect 272064 262268 272116 262274
rect 272064 262210 272116 262216
rect 271236 261520 271288 261526
rect 271236 261462 271288 261468
rect 275940 241466 275968 263463
rect 276124 263362 276152 263463
rect 305880 263463 305882 263472
rect 308402 263528 308404 263537
rect 308456 263528 308458 263537
rect 308402 263463 308458 263472
rect 323030 263528 323086 263537
rect 323030 263463 323086 263472
rect 325790 263528 325846 263537
rect 325790 263463 325846 263472
rect 343454 263528 343510 263537
rect 343454 263463 343510 263472
rect 305828 263434 305880 263440
rect 276112 263356 276164 263362
rect 276112 263298 276164 263304
rect 277306 262304 277362 262313
rect 277306 262239 277362 262248
rect 278686 262304 278742 262313
rect 278686 262239 278742 262248
rect 275928 241460 275980 241466
rect 275928 241402 275980 241408
rect 277320 241398 277348 262239
rect 277308 241392 277360 241398
rect 277308 241334 277360 241340
rect 278700 241330 278728 262239
rect 323044 262138 323072 263463
rect 325804 262206 325832 263463
rect 343468 262886 343496 263463
rect 343546 263120 343602 263129
rect 343546 263055 343602 263064
rect 343560 263022 343588 263055
rect 343548 263016 343600 263022
rect 343548 262958 343600 262964
rect 343456 262880 343508 262886
rect 343456 262822 343508 262828
rect 325792 262200 325844 262206
rect 325792 262142 325844 262148
rect 323032 262132 323084 262138
rect 323032 262074 323084 262080
rect 343560 258074 343588 262958
rect 343468 258046 343588 258074
rect 278688 241324 278740 241330
rect 278688 241266 278740 241272
rect 339408 241256 339460 241262
rect 339408 241198 339460 241204
rect 339420 240281 339448 241198
rect 343468 240922 343496 258046
rect 356624 241466 356652 372574
rect 356612 241460 356664 241466
rect 356612 241402 356664 241408
rect 343456 240916 343508 240922
rect 343456 240858 343508 240864
rect 340052 240848 340104 240854
rect 340052 240790 340104 240796
rect 340064 240281 340092 240790
rect 351552 240780 351604 240786
rect 351552 240722 351604 240728
rect 351564 240281 351592 240722
rect 339406 240272 339462 240281
rect 339406 240207 339462 240216
rect 340050 240272 340106 240281
rect 340050 240207 340106 240216
rect 351550 240272 351606 240281
rect 351550 240207 351606 240216
rect 267740 240100 267792 240106
rect 267740 240042 267792 240048
rect 266452 239896 266504 239902
rect 266452 239838 266504 239844
rect 266360 239828 266412 239834
rect 266360 239770 266412 239776
rect 263600 239692 263652 239698
rect 263600 239634 263652 239640
rect 260840 239420 260892 239426
rect 260840 239362 260892 239368
rect 255320 239352 255372 239358
rect 255320 239294 255372 239300
rect 220820 239284 220872 239290
rect 220820 239226 220872 239232
rect 222108 239284 222160 239290
rect 222108 239226 222160 239232
rect 261022 154592 261078 154601
rect 261022 154527 261078 154536
rect 273534 154592 273590 154601
rect 273534 154527 273590 154536
rect 261036 154290 261064 154527
rect 261024 154284 261076 154290
rect 261024 154226 261076 154232
rect 273548 154222 273576 154527
rect 273536 154216 273588 154222
rect 273536 154158 273588 154164
rect 287978 154184 288034 154193
rect 287978 154119 288034 154128
rect 288162 154184 288218 154193
rect 288162 154119 288218 154128
rect 293314 154184 293370 154193
rect 293314 154119 293316 154128
rect 287992 153921 288020 154119
rect 288176 154086 288204 154119
rect 293368 154119 293370 154128
rect 293316 154090 293368 154096
rect 288164 154080 288216 154086
rect 288164 154022 288216 154028
rect 298466 154048 298522 154057
rect 298466 153983 298468 153992
rect 298520 153983 298522 153992
rect 303434 154048 303490 154057
rect 303434 153983 303490 153992
rect 298468 153954 298520 153960
rect 303448 153950 303476 153983
rect 303436 153944 303488 153950
rect 287978 153912 288034 153921
rect 303436 153886 303488 153892
rect 308402 153912 308458 153921
rect 287978 153847 288034 153856
rect 308402 153847 308404 153856
rect 308456 153847 308458 153856
rect 308404 153818 308456 153824
rect 300860 153196 300912 153202
rect 300860 153138 300912 153144
rect 285680 153128 285732 153134
rect 236090 153096 236146 153105
rect 236090 153031 236146 153040
rect 237378 153096 237434 153105
rect 237378 153031 237434 153040
rect 240138 153096 240194 153105
rect 240138 153031 240194 153040
rect 241518 153096 241574 153105
rect 241518 153031 241574 153040
rect 242898 153096 242954 153105
rect 242898 153031 242954 153040
rect 244278 153096 244334 153105
rect 244278 153031 244334 153040
rect 245658 153096 245714 153105
rect 245658 153031 245714 153040
rect 247038 153096 247094 153105
rect 247038 153031 247094 153040
rect 248418 153096 248474 153105
rect 248418 153031 248474 153040
rect 249798 153096 249854 153105
rect 249798 153031 249854 153040
rect 250258 153096 250314 153105
rect 250258 153031 250314 153040
rect 251178 153096 251234 153105
rect 251178 153031 251234 153040
rect 252558 153096 252614 153105
rect 252558 153031 252614 153040
rect 253570 153096 253626 153105
rect 253570 153031 253626 153040
rect 253938 153096 253994 153105
rect 253938 153031 253994 153040
rect 255318 153096 255374 153105
rect 255318 153031 255374 153040
rect 255962 153096 256018 153105
rect 255962 153031 256018 153040
rect 256698 153096 256754 153105
rect 256698 153031 256754 153040
rect 258078 153096 258134 153105
rect 258078 153031 258134 153040
rect 259550 153096 259606 153105
rect 259550 153031 259606 153040
rect 261206 153096 261262 153105
rect 261206 153031 261262 153040
rect 262218 153096 262274 153105
rect 262218 153031 262274 153040
rect 263598 153096 263654 153105
rect 263598 153031 263654 153040
rect 264978 153096 265034 153105
rect 264978 153031 265034 153040
rect 266358 153096 266414 153105
rect 266358 153031 266414 153040
rect 267738 153096 267794 153105
rect 267738 153031 267794 153040
rect 269118 153096 269174 153105
rect 269118 153031 269174 153040
rect 270498 153096 270554 153105
rect 270498 153031 270554 153040
rect 271878 153096 271934 153105
rect 271878 153031 271934 153040
rect 273258 153096 273314 153105
rect 273258 153031 273314 153040
rect 274730 153096 274786 153105
rect 274730 153031 274786 153040
rect 277950 153096 278006 153105
rect 277950 153031 278006 153040
rect 280066 153096 280122 153105
rect 280066 153031 280122 153040
rect 280250 153096 280306 153105
rect 280250 153031 280306 153040
rect 282918 153096 282974 153105
rect 282918 153031 282974 153040
rect 285678 153096 285680 153105
rect 300872 153105 300900 153138
rect 285732 153096 285734 153105
rect 285678 153031 285734 153040
rect 289818 153096 289874 153105
rect 289818 153031 289820 153040
rect 235998 152416 236054 152425
rect 235998 152351 236054 152360
rect 236012 130354 236040 152351
rect 236104 150414 236132 153031
rect 236092 150408 236144 150414
rect 236092 150350 236144 150356
rect 236000 130348 236052 130354
rect 236000 130290 236052 130296
rect 236104 130286 236132 150350
rect 237392 130529 237420 153031
rect 238758 152008 238814 152017
rect 238758 151943 238814 151952
rect 238772 133754 238800 151943
rect 240152 133822 240180 153031
rect 240140 133816 240192 133822
rect 240140 133758 240192 133764
rect 238760 133748 238812 133754
rect 238760 133690 238812 133696
rect 241532 133278 241560 153031
rect 241520 133272 241572 133278
rect 241520 133214 241572 133220
rect 242912 130626 242940 153031
rect 242900 130620 242952 130626
rect 242900 130562 242952 130568
rect 237378 130520 237434 130529
rect 244292 130490 244320 153031
rect 244370 152416 244426 152425
rect 244370 152351 244426 152360
rect 244384 130694 244412 152351
rect 245672 131102 245700 153031
rect 245660 131096 245712 131102
rect 245660 131038 245712 131044
rect 244372 130688 244424 130694
rect 244372 130630 244424 130636
rect 247052 130558 247080 153031
rect 247130 152416 247186 152425
rect 247130 152351 247132 152360
rect 247184 152351 247186 152360
rect 247132 152322 247184 152328
rect 248432 130762 248460 153031
rect 249812 130937 249840 153031
rect 250272 152454 250300 153031
rect 250260 152448 250312 152454
rect 250260 152390 250312 152396
rect 249798 130928 249854 130937
rect 249798 130863 249854 130872
rect 251192 130830 251220 153031
rect 251270 152416 251326 152425
rect 251270 152351 251326 152360
rect 251284 130898 251312 152351
rect 252572 130966 252600 153031
rect 253584 152590 253612 153031
rect 253572 152584 253624 152590
rect 253572 152526 253624 152532
rect 253952 131034 253980 153031
rect 253940 131028 253992 131034
rect 253940 130970 253992 130976
rect 252560 130960 252612 130966
rect 252560 130902 252612 130908
rect 251272 130892 251324 130898
rect 251272 130834 251324 130840
rect 251180 130824 251232 130830
rect 251180 130766 251232 130772
rect 248420 130756 248472 130762
rect 248420 130698 248472 130704
rect 247040 130552 247092 130558
rect 247040 130494 247092 130500
rect 237378 130455 237434 130464
rect 244280 130484 244332 130490
rect 244280 130426 244332 130432
rect 236092 130280 236144 130286
rect 236092 130222 236144 130228
rect 255332 130218 255360 153031
rect 255976 152726 256004 153031
rect 255964 152720 256016 152726
rect 255964 152662 256016 152668
rect 256712 130422 256740 153031
rect 258092 151230 258120 153031
rect 259458 152688 259514 152697
rect 259458 152623 259514 152632
rect 258262 152552 258318 152561
rect 258262 152487 258264 152496
rect 258316 152487 258318 152496
rect 258264 152458 258316 152464
rect 259472 151434 259500 152623
rect 259460 151428 259512 151434
rect 259460 151370 259512 151376
rect 258080 151224 258132 151230
rect 258080 151166 258132 151172
rect 259564 151026 259592 153031
rect 261220 151366 261248 153031
rect 262232 151502 262260 153031
rect 262220 151496 262272 151502
rect 262220 151438 262272 151444
rect 261208 151360 261260 151366
rect 261208 151302 261260 151308
rect 263612 151298 263640 153031
rect 264992 151570 265020 153031
rect 265070 152688 265126 152697
rect 265070 152623 265072 152632
rect 265124 152623 265126 152632
rect 265072 152594 265124 152600
rect 266372 151638 266400 153031
rect 266450 152688 266506 152697
rect 266450 152623 266506 152632
rect 266360 151632 266412 151638
rect 266360 151574 266412 151580
rect 264980 151564 265032 151570
rect 264980 151506 265032 151512
rect 263600 151292 263652 151298
rect 263600 151234 263652 151240
rect 266464 151162 266492 152623
rect 267752 151706 267780 153031
rect 268016 152788 268068 152794
rect 268016 152730 268068 152736
rect 268028 152697 268056 152730
rect 268014 152688 268070 152697
rect 268014 152623 268070 152632
rect 267740 151700 267792 151706
rect 267740 151642 267792 151648
rect 266452 151156 266504 151162
rect 266452 151098 266504 151104
rect 259552 151020 259604 151026
rect 259552 150962 259604 150968
rect 256700 130416 256752 130422
rect 269132 130393 269160 153031
rect 270512 149734 270540 153031
rect 271892 151094 271920 153031
rect 271880 151088 271932 151094
rect 271880 151030 271932 151036
rect 270500 149728 270552 149734
rect 270500 149670 270552 149676
rect 273272 133890 273300 153031
rect 274638 152688 274694 152697
rect 274638 152623 274694 152632
rect 273260 133884 273312 133890
rect 273260 133826 273312 133832
rect 274652 131073 274680 152623
rect 274744 131170 274772 153031
rect 277964 152998 277992 153031
rect 277952 152992 278004 152998
rect 277952 152934 278004 152940
rect 277398 152008 277454 152017
rect 277398 151943 277454 151952
rect 277412 151706 277440 151943
rect 278686 151872 278742 151881
rect 278686 151807 278742 151816
rect 277400 151700 277452 151706
rect 277400 151642 277452 151648
rect 278044 151700 278096 151706
rect 278044 151642 278096 151648
rect 278056 133210 278084 151642
rect 278044 133204 278096 133210
rect 278044 133146 278096 133152
rect 274732 131164 274784 131170
rect 274732 131106 274784 131112
rect 274638 131064 274694 131073
rect 274638 130999 274694 131008
rect 274744 130422 274772 131106
rect 278700 130490 278728 151807
rect 280080 133210 280108 153031
rect 280264 152930 280292 153031
rect 280252 152924 280304 152930
rect 280252 152866 280304 152872
rect 282932 152862 282960 153031
rect 289872 153031 289874 153040
rect 300858 153096 300914 153105
rect 300858 153031 300914 153040
rect 320178 153096 320234 153105
rect 320178 153031 320234 153040
rect 289820 153002 289872 153008
rect 282920 152856 282972 152862
rect 282920 152798 282972 152804
rect 320192 151774 320220 153031
rect 343546 152824 343602 152833
rect 343546 152759 343602 152768
rect 343560 152658 343588 152759
rect 343548 152652 343600 152658
rect 343548 152594 343600 152600
rect 343546 152552 343602 152561
rect 343546 152487 343548 152496
rect 343600 152487 343602 152496
rect 343548 152458 343600 152464
rect 320180 151768 320232 151774
rect 320180 151710 320232 151716
rect 280068 133204 280120 133210
rect 280068 133146 280120 133152
rect 306380 133204 306432 133210
rect 306380 133146 306432 133152
rect 306392 131850 306420 133146
rect 306380 131844 306432 131850
rect 306380 131786 306432 131792
rect 338488 131096 338540 131102
rect 338488 131038 338540 131044
rect 278688 130484 278740 130490
rect 278688 130426 278740 130432
rect 302240 130484 302292 130490
rect 302240 130426 302292 130432
rect 274732 130416 274784 130422
rect 256700 130358 256752 130364
rect 269118 130384 269174 130393
rect 274732 130358 274784 130364
rect 300768 130416 300820 130422
rect 300768 130358 300820 130364
rect 269118 130319 269174 130328
rect 255320 130212 255372 130218
rect 255320 130154 255372 130160
rect 300780 129742 300808 130358
rect 300768 129736 300820 129742
rect 300768 129678 300820 129684
rect 302252 129062 302280 130426
rect 338500 129849 338528 131038
rect 340604 131028 340656 131034
rect 340604 130970 340656 130976
rect 340616 129849 340644 130970
rect 343560 130490 343588 152458
rect 343548 130484 343600 130490
rect 343548 130426 343600 130432
rect 351736 130416 351788 130422
rect 351736 130358 351788 130364
rect 351748 129849 351776 130358
rect 338486 129840 338542 129849
rect 338486 129775 338542 129784
rect 340602 129840 340658 129849
rect 340602 129775 340658 129784
rect 351734 129840 351790 129849
rect 351734 129775 351790 129784
rect 356624 129742 356652 241402
rect 356612 129736 356664 129742
rect 356612 129678 356664 129684
rect 302240 129056 302292 129062
rect 302240 128998 302292 129004
rect 235998 44840 236054 44849
rect 235998 44775 236054 44784
rect 237102 44840 237158 44849
rect 237102 44775 237158 44784
rect 243082 44840 243138 44849
rect 243082 44775 243138 44784
rect 244278 44840 244334 44849
rect 244278 44775 244334 44784
rect 236012 44606 236040 44775
rect 236000 44600 236052 44606
rect 236000 44542 236052 44548
rect 237116 44538 237144 44775
rect 237104 44532 237156 44538
rect 237104 44474 237156 44480
rect 243096 44470 243124 44775
rect 243084 44464 243136 44470
rect 243084 44406 243136 44412
rect 244292 44062 244320 44775
rect 255870 44704 255926 44713
rect 255870 44639 255926 44648
rect 256974 44704 257030 44713
rect 256974 44639 257030 44648
rect 258078 44704 258134 44713
rect 258078 44639 258134 44648
rect 262862 44704 262918 44713
rect 262862 44639 262918 44648
rect 315854 44704 315910 44713
rect 315854 44639 315910 44648
rect 255884 44402 255912 44639
rect 255872 44396 255924 44402
rect 255872 44338 255924 44344
rect 256988 44334 257016 44639
rect 256976 44328 257028 44334
rect 256976 44270 257028 44276
rect 258092 44266 258120 44639
rect 259458 44568 259514 44577
rect 259458 44503 259514 44512
rect 260654 44568 260710 44577
rect 260654 44503 260710 44512
rect 261758 44568 261814 44577
rect 261758 44503 261814 44512
rect 258080 44260 258132 44266
rect 258080 44202 258132 44208
rect 244280 44056 244332 44062
rect 244280 43998 244332 44004
rect 259472 43994 259500 44503
rect 259460 43988 259512 43994
rect 259460 43930 259512 43936
rect 260668 43790 260696 44503
rect 261772 43858 261800 44503
rect 262876 44198 262904 44639
rect 263874 44568 263930 44577
rect 263874 44503 263930 44512
rect 308494 44568 308550 44577
rect 308494 44503 308550 44512
rect 262864 44192 262916 44198
rect 262864 44134 262916 44140
rect 263888 43926 263916 44503
rect 300858 44160 300914 44169
rect 300858 44095 300914 44104
rect 263876 43920 263928 43926
rect 263876 43862 263928 43868
rect 279238 43888 279294 43897
rect 261760 43852 261812 43858
rect 279238 43823 279294 43832
rect 261760 43794 261812 43800
rect 279252 43790 279280 43823
rect 260656 43784 260708 43790
rect 260656 43726 260708 43732
rect 279240 43784 279292 43790
rect 279240 43726 279292 43732
rect 300872 43518 300900 44095
rect 308508 43722 308536 44503
rect 308496 43716 308548 43722
rect 308496 43658 308548 43664
rect 315868 43654 315896 44639
rect 356716 43722 356744 492118
rect 356808 154018 356836 492526
rect 358360 492516 358412 492522
rect 358360 492458 358412 492464
rect 358268 492448 358320 492454
rect 358268 492390 358320 492396
rect 358176 492244 358228 492250
rect 358176 492186 358228 492192
rect 357164 477488 357216 477494
rect 357164 477430 357216 477436
rect 356888 466132 356940 466138
rect 356888 466074 356940 466080
rect 356900 264246 356928 466074
rect 357072 461032 357124 461038
rect 357072 460974 357124 460980
rect 356980 371544 357032 371550
rect 356980 371486 357032 371492
rect 356888 264240 356940 264246
rect 356888 264182 356940 264188
rect 356888 242684 356940 242690
rect 356888 242626 356940 242632
rect 356900 240854 356928 242626
rect 356992 241398 357020 371486
rect 357084 351354 357112 460974
rect 357176 369374 357204 477430
rect 357256 466404 357308 466410
rect 357256 466346 357308 466352
rect 357268 369782 357296 466346
rect 357348 463616 357400 463622
rect 357348 463558 357400 463564
rect 357360 371142 357388 463558
rect 357900 462052 357952 462058
rect 357900 461994 357952 462000
rect 357440 371272 357492 371278
rect 357440 371214 357492 371220
rect 357348 371136 357400 371142
rect 357348 371078 357400 371084
rect 357256 369776 357308 369782
rect 357256 369718 357308 369724
rect 357164 369368 357216 369374
rect 357164 369310 357216 369316
rect 357072 351348 357124 351354
rect 357072 351290 357124 351296
rect 357084 248414 357112 351290
rect 357452 263022 357480 371214
rect 357912 371210 357940 461994
rect 358084 460828 358136 460834
rect 358084 460770 358136 460776
rect 357992 460148 358044 460154
rect 357992 460090 358044 460096
rect 357900 371204 357952 371210
rect 357900 371146 357952 371152
rect 358004 369850 358032 460090
rect 357992 369844 358044 369850
rect 357992 369786 358044 369792
rect 357532 349852 357584 349858
rect 357532 349794 357584 349800
rect 357440 263016 357492 263022
rect 357440 262958 357492 262964
rect 357084 248386 357296 248414
rect 357268 241534 357296 248386
rect 357256 241528 357308 241534
rect 357256 241470 357308 241476
rect 356980 241392 357032 241398
rect 356980 241334 357032 241340
rect 356888 240848 356940 240854
rect 356888 240790 356940 240796
rect 356796 154012 356848 154018
rect 356796 153954 356848 153960
rect 356900 131034 356928 240790
rect 356992 151706 357020 241334
rect 357268 241262 357296 241470
rect 357544 241330 357572 349794
rect 358096 276010 358124 460770
rect 358084 276004 358136 276010
rect 358084 275946 358136 275952
rect 358084 273284 358136 273290
rect 358084 273226 358136 273232
rect 357716 263628 357768 263634
rect 357716 263570 357768 263576
rect 357532 241324 357584 241330
rect 357532 241266 357584 241272
rect 357256 241256 357308 241262
rect 357256 241198 357308 241204
rect 356980 151700 357032 151706
rect 356980 151642 357032 151648
rect 356980 131844 357032 131850
rect 356980 131786 357032 131792
rect 356992 131646 357020 131786
rect 356980 131640 357032 131646
rect 356980 131582 357032 131588
rect 356888 131028 356940 131034
rect 356888 130970 356940 130976
rect 356796 129056 356848 129062
rect 356796 128998 356848 129004
rect 356704 43716 356756 43722
rect 356704 43658 356756 43664
rect 315856 43648 315908 43654
rect 315856 43590 315908 43596
rect 300860 43512 300912 43518
rect 300860 43454 300912 43460
rect 265162 43208 265218 43217
rect 265162 43143 265218 43152
rect 272154 43208 272210 43217
rect 272154 43143 272210 43152
rect 325882 43208 325938 43217
rect 325882 43143 325938 43152
rect 238114 42800 238170 42809
rect 238114 42735 238170 42744
rect 239126 42800 239182 42809
rect 239126 42735 239182 42744
rect 240506 42800 240562 42809
rect 240506 42735 240562 42744
rect 241610 42800 241666 42809
rect 241610 42735 241666 42744
rect 245290 42800 245346 42809
rect 245290 42735 245346 42744
rect 246394 42800 246450 42809
rect 246394 42735 246450 42744
rect 250074 42800 250130 42809
rect 250074 42735 250130 42744
rect 251178 42800 251234 42809
rect 251178 42735 251234 42744
rect 253386 42800 253442 42809
rect 253386 42735 253442 42744
rect 260930 42800 260986 42809
rect 260930 42735 260986 42744
rect 219992 41404 220044 41410
rect 219992 41346 220044 41352
rect 238128 39982 238156 42735
rect 239140 40730 239168 42735
rect 239128 40724 239180 40730
rect 239128 40666 239180 40672
rect 240520 40050 240548 42735
rect 241624 40662 241652 42735
rect 245304 40798 245332 42735
rect 246408 40866 246436 42735
rect 248602 41984 248658 41993
rect 248602 41919 248658 41928
rect 247682 41848 247738 41857
rect 247682 41783 247738 41792
rect 246396 40860 246448 40866
rect 246396 40802 246448 40808
rect 245292 40792 245344 40798
rect 245292 40734 245344 40740
rect 241612 40656 241664 40662
rect 241612 40598 241664 40604
rect 240508 40044 240560 40050
rect 240508 39986 240560 39992
rect 238116 39976 238168 39982
rect 238116 39918 238168 39924
rect 219900 39704 219952 39710
rect 219900 39646 219952 39652
rect 219716 39636 219768 39642
rect 219716 39578 219768 39584
rect 247696 39438 247724 41783
rect 248616 39506 248644 41919
rect 250088 39953 250116 42735
rect 251192 40934 251220 42735
rect 251730 41984 251786 41993
rect 251730 41919 251786 41928
rect 251180 40928 251232 40934
rect 251180 40870 251232 40876
rect 250074 39944 250130 39953
rect 250074 39879 250130 39888
rect 251744 39574 251772 41919
rect 253400 41002 253428 42735
rect 254122 42120 254178 42129
rect 260944 42090 260972 42735
rect 254122 42055 254178 42064
rect 260932 42084 260984 42090
rect 253388 40996 253440 41002
rect 253388 40938 253440 40944
rect 254136 39642 254164 42055
rect 260932 42026 260984 42032
rect 265176 41070 265204 43143
rect 268198 42800 268254 42809
rect 268198 42735 268254 42744
rect 268474 42800 268530 42809
rect 268474 42735 268530 42744
rect 271234 42800 271290 42809
rect 271234 42735 271290 42744
rect 266358 42392 266414 42401
rect 266358 42327 266414 42336
rect 266634 42392 266690 42401
rect 266634 42327 266690 42336
rect 265164 41064 265216 41070
rect 265164 41006 265216 41012
rect 266372 39710 266400 42327
rect 266648 39778 266676 42327
rect 268212 42158 268240 42735
rect 268200 42152 268252 42158
rect 268200 42094 268252 42100
rect 268488 41138 268516 42735
rect 269762 42392 269818 42401
rect 269762 42327 269818 42336
rect 268476 41132 268528 41138
rect 268476 41074 268528 41080
rect 269776 39846 269804 42327
rect 271248 41206 271276 42735
rect 271236 41200 271288 41206
rect 271236 41142 271288 41148
rect 272168 39914 272196 43143
rect 273258 42800 273314 42809
rect 273258 42735 273314 42744
rect 276110 42800 276166 42809
rect 276110 42735 276166 42744
rect 276938 42800 276994 42809
rect 276938 42735 276994 42744
rect 278318 42800 278374 42809
rect 278318 42735 278374 42744
rect 293314 42800 293370 42809
rect 293314 42735 293370 42744
rect 298466 42800 298522 42809
rect 298466 42735 298522 42744
rect 302514 42800 302570 42809
rect 302514 42735 302570 42744
rect 310978 42800 311034 42809
rect 310978 42735 311034 42744
rect 313370 42800 313426 42809
rect 313370 42735 313426 42744
rect 318338 42800 318394 42809
rect 318338 42735 318394 42744
rect 320914 42800 320970 42809
rect 320914 42735 320916 42744
rect 273272 41274 273300 42735
rect 273534 42256 273590 42265
rect 273534 42191 273590 42200
rect 274730 42256 274786 42265
rect 276124 42226 276152 42735
rect 274730 42191 274786 42200
rect 276112 42220 276164 42226
rect 273260 41268 273312 41274
rect 273260 41210 273312 41216
rect 272156 39908 272208 39914
rect 272156 39850 272208 39856
rect 269764 39840 269816 39846
rect 269764 39782 269816 39788
rect 266636 39772 266688 39778
rect 266636 39714 266688 39720
rect 266360 39704 266412 39710
rect 266360 39646 266412 39652
rect 254124 39636 254176 39642
rect 254124 39578 254176 39584
rect 251732 39568 251784 39574
rect 251732 39510 251784 39516
rect 248604 39500 248656 39506
rect 248604 39442 248656 39448
rect 219164 39432 219216 39438
rect 219164 39374 219216 39380
rect 247684 39432 247736 39438
rect 247684 39374 247736 39380
rect 213552 39364 213604 39370
rect 213552 39306 213604 39312
rect 273548 39302 273576 42191
rect 274744 39370 274772 42191
rect 276112 42162 276164 42168
rect 276952 41342 276980 42735
rect 278332 42226 278360 42735
rect 293328 42362 293356 42735
rect 298480 42430 298508 42735
rect 298468 42424 298520 42430
rect 298468 42366 298520 42372
rect 293316 42356 293368 42362
rect 293316 42298 293368 42304
rect 302528 42294 302556 42735
rect 310992 42566 311020 42735
rect 310980 42560 311032 42566
rect 310980 42502 311032 42508
rect 313384 42498 313412 42735
rect 318352 42634 318380 42735
rect 320968 42735 320970 42744
rect 320916 42706 320968 42712
rect 325896 42702 325924 43143
rect 343178 42800 343234 42809
rect 343178 42735 343180 42744
rect 343232 42735 343234 42744
rect 343454 42800 343510 42809
rect 343454 42735 343510 42744
rect 343180 42706 343232 42712
rect 343468 42702 343496 42735
rect 325884 42696 325936 42702
rect 325884 42638 325936 42644
rect 343456 42696 343508 42702
rect 343456 42638 343508 42644
rect 318340 42628 318392 42634
rect 318340 42570 318392 42576
rect 313372 42492 313424 42498
rect 313372 42434 313424 42440
rect 302516 42288 302568 42294
rect 302516 42230 302568 42236
rect 356808 42226 356836 128998
rect 356992 43790 357020 131582
rect 357440 130484 357492 130490
rect 357440 130426 357492 130432
rect 356980 43784 357032 43790
rect 356980 43726 357032 43732
rect 357452 42702 357480 130426
rect 357544 129062 357572 241266
rect 357624 154420 357676 154426
rect 357624 154362 357676 154368
rect 357636 152658 357664 154362
rect 357624 152652 357676 152658
rect 357624 152594 357676 152600
rect 357532 129056 357584 129062
rect 357532 128998 357584 129004
rect 357636 42770 357664 152594
rect 357728 131646 357756 263570
rect 358096 240786 358124 273226
rect 358084 240780 358136 240786
rect 358084 240722 358136 240728
rect 358096 163538 358124 240722
rect 358084 163532 358136 163538
rect 358084 163474 358136 163480
rect 357716 131640 357768 131646
rect 357716 131582 357768 131588
rect 358096 130422 358124 163474
rect 358084 130416 358136 130422
rect 358084 130358 358136 130364
rect 358084 52488 358136 52494
rect 358084 52430 358136 52436
rect 358096 44130 358124 52430
rect 358084 44124 358136 44130
rect 358084 44066 358136 44072
rect 358188 43518 358216 492186
rect 358280 154562 358308 492390
rect 358268 154556 358320 154562
rect 358268 154498 358320 154504
rect 358372 154494 358400 492458
rect 362316 492380 362368 492386
rect 362316 492322 362368 492328
rect 362224 492040 362276 492046
rect 362224 491982 362276 491988
rect 359464 490816 359516 490822
rect 359464 490758 359516 490764
rect 358636 480208 358688 480214
rect 358636 480150 358688 480156
rect 358452 474088 358504 474094
rect 358452 474030 358504 474036
rect 358360 154488 358412 154494
rect 358360 154430 358412 154436
rect 358464 153134 358492 474030
rect 358544 463140 358596 463146
rect 358544 463082 358596 463088
rect 358452 153128 358504 153134
rect 358452 153070 358504 153076
rect 358556 151745 358584 463082
rect 358648 374746 358676 480150
rect 358728 466200 358780 466206
rect 358728 466142 358780 466148
rect 358636 374740 358688 374746
rect 358636 374682 358688 374688
rect 358740 370938 358768 466142
rect 358820 458312 358872 458318
rect 358820 458254 358872 458260
rect 358832 454753 358860 458254
rect 358818 454744 358874 454753
rect 358818 454679 358874 454688
rect 358728 370932 358780 370938
rect 358728 370874 358780 370880
rect 358832 354674 358860 454679
rect 358910 393816 358966 393825
rect 358910 393751 358966 393760
rect 358924 363662 358952 393751
rect 359002 390824 359058 390833
rect 359002 390759 359058 390768
rect 359016 368014 359044 390759
rect 359094 388104 359150 388113
rect 359094 388039 359150 388048
rect 359004 368008 359056 368014
rect 359004 367950 359056 367956
rect 359016 367810 359044 367950
rect 359004 367804 359056 367810
rect 359004 367746 359056 367752
rect 359108 366353 359136 388039
rect 359476 383586 359504 490758
rect 359556 489388 359608 489394
rect 359556 489330 359608 489336
rect 359568 385014 359596 489330
rect 359832 487892 359884 487898
rect 359832 487834 359884 487840
rect 359648 474564 359700 474570
rect 359648 474506 359700 474512
rect 359556 385008 359608 385014
rect 359556 384950 359608 384956
rect 359464 383580 359516 383586
rect 359464 383522 359516 383528
rect 359280 371612 359332 371618
rect 359280 371554 359332 371560
rect 359094 366344 359150 366353
rect 359094 366279 359150 366288
rect 359108 364334 359136 366279
rect 359108 364306 359228 364334
rect 358912 363656 358964 363662
rect 358912 363598 358964 363604
rect 358924 359582 358952 363598
rect 358912 359576 358964 359582
rect 358912 359518 358964 359524
rect 359096 359508 359148 359514
rect 359096 359450 359148 359456
rect 359004 356720 359056 356726
rect 359004 356662 359056 356668
rect 358832 354646 358952 354674
rect 358924 344185 358952 354646
rect 358910 344176 358966 344185
rect 358910 344111 358966 344120
rect 358818 284336 358874 284345
rect 358818 284271 358874 284280
rect 358832 175001 358860 284271
rect 358924 234025 358952 344111
rect 359016 280129 359044 356662
rect 359108 287054 359136 359450
rect 359200 358766 359228 364306
rect 359188 358760 359240 358766
rect 359188 358702 359240 358708
rect 359108 287026 359228 287054
rect 359200 282441 359228 287026
rect 359186 282432 359242 282441
rect 359186 282367 359242 282376
rect 359002 280120 359058 280129
rect 359002 280055 359058 280064
rect 359094 278760 359150 278769
rect 359094 278695 359150 278704
rect 358910 234016 358966 234025
rect 358910 233951 358966 233960
rect 358818 174992 358874 175001
rect 358818 174927 358874 174936
rect 358818 172408 358874 172417
rect 358818 172343 358874 172352
rect 358832 171329 358860 172343
rect 358818 171320 358874 171329
rect 358818 171255 358874 171264
rect 358542 151736 358598 151745
rect 358542 151671 358598 151680
rect 358728 130416 358780 130422
rect 358728 130358 358780 130364
rect 358740 53106 358768 130358
rect 358832 61985 358860 171255
rect 359108 171134 359136 278695
rect 359200 172689 359228 282367
rect 359292 263634 359320 371554
rect 359660 370870 359688 474506
rect 359740 471912 359792 471918
rect 359740 471854 359792 471860
rect 359752 374814 359780 471854
rect 359844 403646 359872 487834
rect 360936 482316 360988 482322
rect 360936 482258 360988 482264
rect 360752 469124 360804 469130
rect 360752 469066 360804 469072
rect 360108 461100 360160 461106
rect 360108 461042 360160 461048
rect 359924 459400 359976 459406
rect 359924 459342 359976 459348
rect 359936 405006 359964 459342
rect 359924 405000 359976 405006
rect 359924 404942 359976 404948
rect 359832 403640 359884 403646
rect 359832 403582 359884 403588
rect 359922 392184 359978 392193
rect 359922 392119 359978 392128
rect 359830 389328 359886 389337
rect 359830 389263 359886 389272
rect 359740 374808 359792 374814
rect 359740 374750 359792 374756
rect 359648 370864 359700 370870
rect 359648 370806 359700 370812
rect 359556 368008 359608 368014
rect 359556 367950 359608 367956
rect 359464 358760 359516 358766
rect 359464 358702 359516 358708
rect 359476 358086 359504 358702
rect 359464 358080 359516 358086
rect 359464 358022 359516 358028
rect 359370 280120 359426 280129
rect 359370 280055 359426 280064
rect 359280 263628 359332 263634
rect 359280 263570 359332 263576
rect 359278 234016 359334 234025
rect 359278 233951 359334 233960
rect 359186 172680 359242 172689
rect 359186 172615 359242 172624
rect 359016 171106 359136 171134
rect 358910 169824 358966 169833
rect 358910 169759 358966 169768
rect 358818 61976 358874 61985
rect 358818 61911 358874 61920
rect 358924 60489 358952 169759
rect 359016 168609 359044 171106
rect 359002 168600 359058 168609
rect 359002 168535 359058 168544
rect 358910 60480 358966 60489
rect 358910 60415 358966 60424
rect 359016 59265 359044 168535
rect 359200 63345 359228 172615
rect 359292 124137 359320 233951
rect 359384 169833 359412 280055
rect 359476 278769 359504 358022
rect 359568 356794 359596 367950
rect 359844 360874 359872 389263
rect 359936 366382 359964 392119
rect 360120 389366 360148 461042
rect 360660 459468 360712 459474
rect 360660 459410 360712 459416
rect 360108 389360 360160 389366
rect 360108 389302 360160 389308
rect 360292 371340 360344 371346
rect 360292 371282 360344 371288
rect 359924 366376 359976 366382
rect 359924 366318 359976 366324
rect 359832 360868 359884 360874
rect 359832 360810 359884 360816
rect 359648 359576 359700 359582
rect 359648 359518 359700 359524
rect 359556 356788 359608 356794
rect 359556 356730 359608 356736
rect 359568 281489 359596 356730
rect 359660 284345 359688 359518
rect 359844 356726 359872 360810
rect 359936 359514 359964 366318
rect 359924 359508 359976 359514
rect 359924 359450 359976 359456
rect 359832 356720 359884 356726
rect 359832 356662 359884 356668
rect 360200 351280 360252 351286
rect 360200 351222 360252 351228
rect 359646 284336 359702 284345
rect 359646 284271 359702 284280
rect 359554 281480 359610 281489
rect 359554 281415 359610 281424
rect 359462 278760 359518 278769
rect 359462 278695 359518 278704
rect 359568 277394 359596 281415
rect 359568 277366 359688 277394
rect 359464 240916 359516 240922
rect 359464 240858 359516 240864
rect 359370 169824 359426 169833
rect 359370 169759 359426 169768
rect 359476 152522 359504 240858
rect 359554 174992 359610 175001
rect 359554 174927 359610 174936
rect 359464 152516 359516 152522
rect 359464 152458 359516 152464
rect 359278 124128 359334 124137
rect 359278 124063 359334 124072
rect 359568 64705 359596 174927
rect 359660 172417 359688 277366
rect 360212 274650 360240 351222
rect 360200 274644 360252 274650
rect 360200 274586 360252 274592
rect 360212 273290 360240 274586
rect 360200 273284 360252 273290
rect 360200 273226 360252 273232
rect 360304 262886 360332 371282
rect 360672 369238 360700 459410
rect 360764 374610 360792 469066
rect 360844 462120 360896 462126
rect 360844 462062 360896 462068
rect 360856 406434 360884 462062
rect 360844 406428 360896 406434
rect 360844 406370 360896 406376
rect 360844 382288 360896 382294
rect 360844 382230 360896 382236
rect 360752 374604 360804 374610
rect 360752 374546 360804 374552
rect 360660 369232 360712 369238
rect 360660 369174 360712 369180
rect 360856 351286 360884 382230
rect 360844 351280 360896 351286
rect 360844 351222 360896 351228
rect 360292 262880 360344 262886
rect 360292 262822 360344 262828
rect 360200 241528 360252 241534
rect 360200 241470 360252 241476
rect 359646 172408 359702 172417
rect 359646 172343 359702 172352
rect 360212 131102 360240 241470
rect 360304 154426 360332 262822
rect 360292 154420 360344 154426
rect 360292 154362 360344 154368
rect 360200 131096 360252 131102
rect 360200 131038 360252 131044
rect 359554 64696 359610 64705
rect 359554 64631 359610 64640
rect 359186 63336 359242 63345
rect 359186 63271 359242 63280
rect 359002 59256 359058 59265
rect 359002 59191 359058 59200
rect 358728 53100 358780 53106
rect 358728 53042 358780 53048
rect 358740 52494 358768 53042
rect 358728 52488 358780 52494
rect 358728 52430 358780 52436
rect 358176 43512 358228 43518
rect 358176 43454 358228 43460
rect 357624 42764 357676 42770
rect 357624 42706 357676 42712
rect 357440 42696 357492 42702
rect 357440 42638 357492 42644
rect 360948 42634 360976 482258
rect 361304 478304 361356 478310
rect 361304 478246 361356 478252
rect 361120 472728 361172 472734
rect 361120 472670 361172 472676
rect 361028 465792 361080 465798
rect 361028 465734 361080 465740
rect 360936 42628 360988 42634
rect 360936 42570 360988 42576
rect 361040 42430 361068 465734
rect 361132 153202 361160 472670
rect 361212 463004 361264 463010
rect 361212 462946 361264 462952
rect 361120 153196 361172 153202
rect 361120 153138 361172 153144
rect 361224 151609 361252 462946
rect 361316 263294 361344 478246
rect 361396 474428 361448 474434
rect 361396 474370 361448 474376
rect 361408 370802 361436 474370
rect 361488 471572 361540 471578
rect 361488 471514 361540 471520
rect 361500 374542 361528 471514
rect 361580 460964 361632 460970
rect 361580 460906 361632 460912
rect 361592 383654 361620 460906
rect 361672 389360 361724 389366
rect 361672 389302 361724 389308
rect 361580 383648 361632 383654
rect 361580 383590 361632 383596
rect 361592 382294 361620 383590
rect 361580 382288 361632 382294
rect 361580 382230 361632 382236
rect 361488 374536 361540 374542
rect 361488 374478 361540 374484
rect 361396 370796 361448 370802
rect 361396 370738 361448 370744
rect 361684 354674 361712 389302
rect 361592 354646 361712 354674
rect 361592 351354 361620 354646
rect 361580 351348 361632 351354
rect 361580 351290 361632 351296
rect 361304 263288 361356 263294
rect 361304 263230 361356 263236
rect 361592 242690 361620 351290
rect 361580 242684 361632 242690
rect 361580 242626 361632 242632
rect 361210 151600 361266 151609
rect 361210 151535 361266 151544
rect 362236 44441 362264 491982
rect 362328 154426 362356 492322
rect 366548 492312 366600 492318
rect 366548 492254 366600 492260
rect 366364 492108 366416 492114
rect 366364 492050 366416 492056
rect 363604 491972 363656 491978
rect 363604 491914 363656 491920
rect 362684 480140 362736 480146
rect 362684 480082 362736 480088
rect 362408 470008 362460 470014
rect 362408 469950 362460 469956
rect 362420 165578 362448 469950
rect 362500 468988 362552 468994
rect 362500 468930 362552 468936
rect 362512 263566 362540 468930
rect 362592 468920 362644 468926
rect 362592 468862 362644 468868
rect 362604 264722 362632 468862
rect 362696 367946 362724 480082
rect 362776 474496 362828 474502
rect 362776 474438 362828 474444
rect 362788 369578 362816 474438
rect 363512 461848 363564 461854
rect 363512 461790 363564 461796
rect 362868 459264 362920 459270
rect 362868 459206 362920 459212
rect 362880 373386 362908 459206
rect 363420 459196 363472 459202
rect 363420 459138 363472 459144
rect 363432 373726 363460 459138
rect 363524 374270 363552 461790
rect 363512 374264 363564 374270
rect 363512 374206 363564 374212
rect 363420 373720 363472 373726
rect 363420 373662 363472 373668
rect 362868 373380 362920 373386
rect 362868 373322 362920 373328
rect 362776 369572 362828 369578
rect 362776 369514 362828 369520
rect 362684 367940 362736 367946
rect 362684 367882 362736 367888
rect 362592 264716 362644 264722
rect 362592 264658 362644 264664
rect 362500 263560 362552 263566
rect 362500 263502 362552 263508
rect 362408 165572 362460 165578
rect 362408 165514 362460 165520
rect 362316 154420 362368 154426
rect 362316 154362 362368 154368
rect 362222 44432 362278 44441
rect 362222 44367 362278 44376
rect 363616 44198 363644 491914
rect 363696 486464 363748 486470
rect 363696 486406 363748 486412
rect 363604 44192 363656 44198
rect 363604 44134 363656 44140
rect 361028 42424 361080 42430
rect 361028 42366 361080 42372
rect 278320 42220 278372 42226
rect 278320 42162 278372 42168
rect 356796 42220 356848 42226
rect 356796 42162 356848 42168
rect 363708 42158 363736 486406
rect 364984 485104 365036 485110
rect 364984 485046 365036 485052
rect 363788 481092 363840 481098
rect 363788 481034 363840 481040
rect 363800 152862 363828 481034
rect 364156 480072 364208 480078
rect 364156 480014 364208 480020
rect 363972 471300 364024 471306
rect 363972 471242 364024 471248
rect 363880 463276 363932 463282
rect 363880 463218 363932 463224
rect 363892 264450 363920 463218
rect 363984 273222 364012 471242
rect 364064 460692 364116 460698
rect 364064 460634 364116 460640
rect 363972 273216 364024 273222
rect 363972 273158 364024 273164
rect 363880 264444 363932 264450
rect 363880 264386 363932 264392
rect 364076 263362 364104 460634
rect 364168 367878 364196 480014
rect 364892 474360 364944 474366
rect 364892 474302 364944 474308
rect 364248 471844 364300 471850
rect 364248 471786 364300 471792
rect 364260 373318 364288 471786
rect 364800 464432 364852 464438
rect 364800 464374 364852 464380
rect 364812 373522 364840 464374
rect 364800 373516 364852 373522
rect 364800 373458 364852 373464
rect 364248 373312 364300 373318
rect 364248 373254 364300 373260
rect 364904 369646 364932 474302
rect 364892 369640 364944 369646
rect 364892 369582 364944 369588
rect 364156 367872 364208 367878
rect 364156 367814 364208 367820
rect 364064 263356 364116 263362
rect 364064 263298 364116 263304
rect 363788 152856 363840 152862
rect 363788 152798 363840 152804
rect 364996 42566 365024 485046
rect 365076 480956 365128 480962
rect 365076 480898 365128 480904
rect 365088 42702 365116 480898
rect 365628 479936 365680 479942
rect 365628 479878 365680 479884
rect 365352 476944 365404 476950
rect 365352 476886 365404 476892
rect 365168 469940 365220 469946
rect 365168 469882 365220 469888
rect 365180 152726 365208 469882
rect 365260 460420 365312 460426
rect 365260 460362 365312 460368
rect 365272 154358 365300 460362
rect 365364 263158 365392 476886
rect 365444 468852 365496 468858
rect 365444 468794 365496 468800
rect 365352 263152 365404 263158
rect 365352 263094 365404 263100
rect 365456 262206 365484 468794
rect 365536 463208 365588 463214
rect 365536 463150 365588 463156
rect 365548 264654 365576 463150
rect 365640 373250 365668 479878
rect 366272 463480 366324 463486
rect 366272 463422 366324 463428
rect 366180 463344 366232 463350
rect 366180 463286 366232 463292
rect 366192 373862 366220 463286
rect 366180 373856 366232 373862
rect 366180 373798 366232 373804
rect 365628 373244 365680 373250
rect 365628 373186 365680 373192
rect 366284 371074 366312 463422
rect 366272 371068 366324 371074
rect 366272 371010 366324 371016
rect 365536 264648 365588 264654
rect 365536 264590 365588 264596
rect 365444 262200 365496 262206
rect 365444 262142 365496 262148
rect 365260 154352 365312 154358
rect 365260 154294 365312 154300
rect 365168 152720 365220 152726
rect 365168 152662 365220 152668
rect 366376 43654 366404 492050
rect 366456 489252 366508 489258
rect 366456 489194 366508 489200
rect 366468 55214 366496 489194
rect 366560 153814 366588 492254
rect 368112 490748 368164 490754
rect 368112 490690 368164 490696
rect 366732 487824 366784 487830
rect 366732 487766 366784 487772
rect 366640 460624 366692 460630
rect 366640 460566 366692 460572
rect 366652 154154 366680 460566
rect 366744 262721 366772 487766
rect 367836 482384 367888 482390
rect 367836 482326 367888 482332
rect 366916 480004 366968 480010
rect 366916 479946 366968 479952
rect 366824 466064 366876 466070
rect 366824 466006 366876 466012
rect 366836 264518 366864 466006
rect 366928 367810 366956 479946
rect 367744 475380 367796 475386
rect 367744 475322 367796 475328
rect 367652 471708 367704 471714
rect 367652 471650 367704 471656
rect 367008 471504 367060 471510
rect 367008 471446 367060 471452
rect 367020 374338 367048 471446
rect 367560 468444 367612 468450
rect 367560 468386 367612 468392
rect 367008 374332 367060 374338
rect 367008 374274 367060 374280
rect 367572 372094 367600 468386
rect 367664 373658 367692 471650
rect 367652 373652 367704 373658
rect 367652 373594 367704 373600
rect 367560 372088 367612 372094
rect 367560 372030 367612 372036
rect 366916 367804 366968 367810
rect 366916 367746 366968 367752
rect 366824 264512 366876 264518
rect 366824 264454 366876 264460
rect 366730 262712 366786 262721
rect 366730 262647 366786 262656
rect 366640 154148 366692 154154
rect 366640 154090 366692 154096
rect 366548 153808 366600 153814
rect 366548 153750 366600 153756
rect 366456 55208 366508 55214
rect 366456 55150 366508 55156
rect 366364 43648 366416 43654
rect 366364 43590 366416 43596
rect 365076 42696 365128 42702
rect 365076 42638 365128 42644
rect 364984 42560 365036 42566
rect 364984 42502 365036 42508
rect 367756 42498 367784 475322
rect 367848 164218 367876 482326
rect 368020 460556 368072 460562
rect 368020 460498 368072 460504
rect 367928 458924 367980 458930
rect 367928 458866 367980 458872
rect 367836 164212 367888 164218
rect 367836 164154 367888 164160
rect 367940 152289 367968 458866
rect 368032 153950 368060 460498
rect 368124 263498 368152 490690
rect 376116 490680 376168 490686
rect 376116 490622 376168 490628
rect 376024 490612 376076 490618
rect 376024 490554 376076 490560
rect 370596 489320 370648 489326
rect 370596 489262 370648 489268
rect 369308 485240 369360 485246
rect 369308 485182 369360 485188
rect 369124 479528 369176 479534
rect 369124 479470 369176 479476
rect 368388 477420 368440 477426
rect 368388 477362 368440 477368
rect 368296 477080 368348 477086
rect 368296 477022 368348 477028
rect 368204 468784 368256 468790
rect 368204 468726 368256 468732
rect 368216 264858 368244 468726
rect 368308 370734 368336 477022
rect 368400 373794 368428 477362
rect 369032 471776 369084 471782
rect 369032 471718 369084 471724
rect 368940 463548 368992 463554
rect 368940 463490 368992 463496
rect 368388 373788 368440 373794
rect 368388 373730 368440 373736
rect 368952 372366 368980 463490
rect 368940 372360 368992 372366
rect 368940 372302 368992 372308
rect 368386 372056 368442 372065
rect 368386 371991 368442 372000
rect 368296 370728 368348 370734
rect 368296 370670 368348 370676
rect 368204 264852 368256 264858
rect 368204 264794 368256 264800
rect 368112 263492 368164 263498
rect 368112 263434 368164 263440
rect 368400 243574 368428 371991
rect 369044 371006 369072 471718
rect 369032 371000 369084 371006
rect 369032 370942 369084 370948
rect 368388 243568 368440 243574
rect 368388 243510 368440 243516
rect 368020 153944 368072 153950
rect 368020 153886 368072 153892
rect 369136 152930 369164 479470
rect 369216 460488 369268 460494
rect 369216 460430 369268 460436
rect 369228 154086 369256 460430
rect 369320 263022 369348 485182
rect 369584 479868 369636 479874
rect 369584 479810 369636 479816
rect 369400 478236 369452 478242
rect 369400 478178 369452 478184
rect 369308 263016 369360 263022
rect 369308 262958 369360 262964
rect 369412 262954 369440 478178
rect 369492 459060 369544 459066
rect 369492 459002 369544 459008
rect 369504 264314 369532 459002
rect 369596 369102 369624 479810
rect 369676 474292 369728 474298
rect 369676 474234 369728 474240
rect 369688 373930 369716 474234
rect 370412 469192 370464 469198
rect 370412 469134 370464 469140
rect 370320 464500 370372 464506
rect 370320 464442 370372 464448
rect 369676 373924 369728 373930
rect 369676 373866 369728 373872
rect 369768 372632 369820 372638
rect 369768 372574 369820 372580
rect 369676 371816 369728 371822
rect 369676 371758 369728 371764
rect 369584 369096 369636 369102
rect 369584 369038 369636 369044
rect 369492 264308 369544 264314
rect 369492 264250 369544 264256
rect 369400 262948 369452 262954
rect 369400 262890 369452 262896
rect 369688 240718 369716 371758
rect 369676 240712 369728 240718
rect 369676 240654 369728 240660
rect 369780 239902 369808 372574
rect 370332 372570 370360 464442
rect 370320 372564 370372 372570
rect 370320 372506 370372 372512
rect 370424 370394 370452 469134
rect 370504 465724 370556 465730
rect 370504 465666 370556 465672
rect 370412 370388 370464 370394
rect 370412 370330 370464 370336
rect 369768 239896 369820 239902
rect 369768 239838 369820 239844
rect 369216 154080 369268 154086
rect 369216 154022 369268 154028
rect 369124 152924 369176 152930
rect 369124 152866 369176 152872
rect 367926 152280 367982 152289
rect 367926 152215 367982 152224
rect 367744 42492 367796 42498
rect 367744 42434 367796 42440
rect 370516 42362 370544 465666
rect 370608 152969 370636 489262
rect 370688 486532 370740 486538
rect 370688 486474 370740 486480
rect 370594 152960 370650 152969
rect 370594 152895 370650 152904
rect 370700 152590 370728 486474
rect 371976 485172 372028 485178
rect 371976 485114 372028 485120
rect 371148 477352 371200 477358
rect 371148 477294 371200 477300
rect 370872 471368 370924 471374
rect 370872 471310 370924 471316
rect 370780 463072 370832 463078
rect 370780 463014 370832 463020
rect 370792 153882 370820 463014
rect 370884 263430 370912 471310
rect 371056 461644 371108 461650
rect 371056 461586 371108 461592
rect 370964 458992 371016 458998
rect 370964 458934 371016 458940
rect 370976 264178 371004 458934
rect 371068 374134 371096 461586
rect 371056 374128 371108 374134
rect 371056 374070 371108 374076
rect 371056 371952 371108 371958
rect 371056 371894 371108 371900
rect 371068 371414 371096 371894
rect 371056 371408 371108 371414
rect 371056 371350 371108 371356
rect 370964 264172 371016 264178
rect 370964 264114 371016 264120
rect 370872 263424 370924 263430
rect 370872 263366 370924 263372
rect 371068 243710 371096 371350
rect 371160 369170 371188 477294
rect 371792 477148 371844 477154
rect 371792 477090 371844 477096
rect 371700 463412 371752 463418
rect 371700 463354 371752 463360
rect 371712 373454 371740 463354
rect 371700 373448 371752 373454
rect 371700 373390 371752 373396
rect 371804 370326 371832 477090
rect 371884 467152 371936 467158
rect 371884 467094 371936 467100
rect 371792 370320 371844 370326
rect 371792 370262 371844 370268
rect 371148 369164 371200 369170
rect 371148 369106 371200 369112
rect 371792 369096 371844 369102
rect 371792 369038 371844 369044
rect 371148 367804 371200 367810
rect 371148 367746 371200 367752
rect 371056 243704 371108 243710
rect 371056 243646 371108 243652
rect 371160 240106 371188 367746
rect 371804 263634 371832 369038
rect 371792 263628 371844 263634
rect 371792 263570 371844 263576
rect 371148 240100 371200 240106
rect 371148 240042 371200 240048
rect 370780 153876 370832 153882
rect 370780 153818 370832 153824
rect 370688 152584 370740 152590
rect 370688 152526 370740 152532
rect 370504 42356 370556 42362
rect 370504 42298 370556 42304
rect 371896 42294 371924 467094
rect 371988 152658 372016 485114
rect 373448 482452 373500 482458
rect 373448 482394 373500 482400
rect 373264 476876 373316 476882
rect 373264 476818 373316 476824
rect 373172 474632 373224 474638
rect 373172 474574 373224 474580
rect 372436 474224 372488 474230
rect 372436 474166 372488 474172
rect 372252 474156 372304 474162
rect 372252 474098 372304 474104
rect 372068 474020 372120 474026
rect 372068 473962 372120 473968
rect 371976 152652 372028 152658
rect 371976 152594 372028 152600
rect 372080 152386 372108 473962
rect 372160 460284 372212 460290
rect 372160 460226 372212 460232
rect 372172 154290 372200 460226
rect 372264 263226 372292 474098
rect 372344 465996 372396 466002
rect 372344 465938 372396 465944
rect 372356 264382 372384 465938
rect 372448 374678 372476 474166
rect 373080 466268 373132 466274
rect 373080 466210 373132 466216
rect 372528 461984 372580 461990
rect 372528 461926 372580 461932
rect 372436 374672 372488 374678
rect 372436 374614 372488 374620
rect 372434 371920 372490 371929
rect 372540 371890 372568 461926
rect 372988 459128 373040 459134
rect 372988 459070 373040 459076
rect 372896 374740 372948 374746
rect 372896 374682 372948 374688
rect 372908 374474 372936 374682
rect 372896 374468 372948 374474
rect 372896 374410 372948 374416
rect 373000 374202 373028 459070
rect 372988 374196 373040 374202
rect 372988 374138 373040 374144
rect 373092 372162 373120 466210
rect 373080 372156 373132 372162
rect 373080 372098 373132 372104
rect 373184 372042 373212 474574
rect 373092 372014 373212 372042
rect 372434 371855 372490 371864
rect 372528 371884 372580 371890
rect 372344 264376 372396 264382
rect 372344 264318 372396 264324
rect 372252 263220 372304 263226
rect 372252 263162 372304 263168
rect 372448 244254 372476 371855
rect 372528 371826 372580 371832
rect 372436 244248 372488 244254
rect 372436 244190 372488 244196
rect 372540 240922 372568 371826
rect 373092 370666 373120 372014
rect 373172 371476 373224 371482
rect 373172 371418 373224 371424
rect 373080 370660 373132 370666
rect 373080 370602 373132 370608
rect 373080 369232 373132 369238
rect 373080 369174 373132 369180
rect 372986 369064 373042 369073
rect 372986 368999 373042 369008
rect 373000 262002 373028 368999
rect 373092 364334 373120 369174
rect 373184 368014 373212 371418
rect 373172 368008 373224 368014
rect 373172 367950 373224 367956
rect 373092 364306 373212 364334
rect 373080 264784 373132 264790
rect 373080 264726 373132 264732
rect 372988 261996 373040 262002
rect 372988 261938 373040 261944
rect 372528 240916 372580 240922
rect 372528 240858 372580 240864
rect 372528 240712 372580 240718
rect 372528 240654 372580 240660
rect 372436 238808 372488 238814
rect 372436 238750 372488 238756
rect 372160 154284 372212 154290
rect 372160 154226 372212 154232
rect 372068 152380 372120 152386
rect 372068 152322 372120 152328
rect 372448 151094 372476 238750
rect 372436 151088 372488 151094
rect 372436 151030 372488 151036
rect 372436 133612 372488 133618
rect 372436 133554 372488 133560
rect 371884 42288 371936 42294
rect 371884 42230 371936 42236
rect 363696 42152 363748 42158
rect 363696 42094 363748 42100
rect 276940 41336 276992 41342
rect 276940 41278 276992 41284
rect 372448 39506 372476 133554
rect 372540 130354 372568 240654
rect 372528 130348 372580 130354
rect 372528 130290 372580 130296
rect 373092 129742 373120 264726
rect 373184 262070 373212 364306
rect 373172 262064 373224 262070
rect 373172 262006 373224 262012
rect 373172 240100 373224 240106
rect 373172 240042 373224 240048
rect 373184 239426 373212 240042
rect 373172 239420 373224 239426
rect 373172 239362 373224 239368
rect 373184 151162 373212 239362
rect 373276 152998 373304 476818
rect 373356 460352 373408 460358
rect 373356 460294 373408 460300
rect 373368 154222 373396 460294
rect 373460 263401 373488 482394
rect 373724 479732 373776 479738
rect 373724 479674 373776 479680
rect 373540 472796 373592 472802
rect 373540 472738 373592 472744
rect 373446 263392 373502 263401
rect 373446 263327 373502 263336
rect 373552 263090 373580 472738
rect 373632 468716 373684 468722
rect 373632 468658 373684 468664
rect 373644 264926 373672 468658
rect 373736 371482 373764 479674
rect 374828 479596 374880 479602
rect 374828 479538 374880 479544
rect 374644 478168 374696 478174
rect 374644 478110 374696 478116
rect 374460 477284 374512 477290
rect 374460 477226 374512 477232
rect 374000 461916 374052 461922
rect 374000 461858 374052 461864
rect 374012 374490 374040 461858
rect 373816 374468 373868 374474
rect 373816 374410 373868 374416
rect 373920 374462 374040 374490
rect 373724 371476 373776 371482
rect 373724 371418 373776 371424
rect 373724 369436 373776 369442
rect 373724 369378 373776 369384
rect 373736 364334 373764 369378
rect 373828 369186 373856 374410
rect 373920 374066 373948 374462
rect 373908 374060 373960 374066
rect 373908 374002 373960 374008
rect 373920 369442 373948 374002
rect 374472 370530 374500 477226
rect 374552 459332 374604 459338
rect 374552 459274 374604 459280
rect 374564 371686 374592 459274
rect 374552 371680 374604 371686
rect 374552 371622 374604 371628
rect 374552 370728 374604 370734
rect 374552 370670 374604 370676
rect 374564 370598 374592 370670
rect 374552 370592 374604 370598
rect 374552 370534 374604 370540
rect 374460 370524 374512 370530
rect 374460 370466 374512 370472
rect 373908 369436 373960 369442
rect 373908 369378 373960 369384
rect 373828 369158 373948 369186
rect 373736 364306 373856 364334
rect 373632 264920 373684 264926
rect 373632 264862 373684 264868
rect 373632 263628 373684 263634
rect 373632 263570 373684 263576
rect 373540 263084 373592 263090
rect 373540 263026 373592 263032
rect 373540 243704 373592 243710
rect 373540 243646 373592 243652
rect 373448 243568 373500 243574
rect 373448 243510 373500 243516
rect 373356 154216 373408 154222
rect 373356 154158 373408 154164
rect 373264 152992 373316 152998
rect 373264 152934 373316 152940
rect 373172 151156 373224 151162
rect 373172 151098 373224 151104
rect 373460 133618 373488 243510
rect 373448 133612 373500 133618
rect 373448 133554 373500 133560
rect 373552 133210 373580 243646
rect 373644 153270 373672 263570
rect 373828 241194 373856 364306
rect 373920 263702 373948 369158
rect 374460 367872 374512 367878
rect 374460 367814 374512 367820
rect 374472 264790 374500 367814
rect 374460 264784 374512 264790
rect 374460 264726 374512 264732
rect 373908 263696 373960 263702
rect 373908 263638 373960 263644
rect 374368 263696 374420 263702
rect 374368 263638 374420 263644
rect 373816 241188 373868 241194
rect 373816 241130 373868 241136
rect 373828 238754 373856 241130
rect 373736 238726 373856 238754
rect 373632 153264 373684 153270
rect 373632 153206 373684 153212
rect 373540 133204 373592 133210
rect 373540 133146 373592 133152
rect 373736 130490 373764 238726
rect 373816 153264 373868 153270
rect 373816 153206 373868 153212
rect 373724 130484 373776 130490
rect 373724 130426 373776 130432
rect 373080 129736 373132 129742
rect 373080 129678 373132 129684
rect 373828 39846 373856 153206
rect 374380 133793 374408 263638
rect 374564 248414 374592 370534
rect 374472 248386 374592 248414
rect 374472 241466 374500 248386
rect 374552 244248 374604 244254
rect 374552 244190 374604 244196
rect 374564 243642 374592 244190
rect 374552 243636 374604 243642
rect 374552 243578 374604 243584
rect 374460 241460 374512 241466
rect 374460 241402 374512 241408
rect 374552 240644 374604 240650
rect 374552 240586 374604 240592
rect 374460 151088 374512 151094
rect 374460 151030 374512 151036
rect 374366 133784 374422 133793
rect 374366 133719 374422 133728
rect 373908 132524 373960 132530
rect 373908 132466 373960 132472
rect 373920 41070 373948 132466
rect 373908 41064 373960 41070
rect 373908 41006 373960 41012
rect 374472 39914 374500 151030
rect 374564 150958 374592 240586
rect 374656 152794 374684 478110
rect 374736 460216 374788 460222
rect 374736 460158 374788 460164
rect 374644 152788 374696 152794
rect 374644 152730 374696 152736
rect 374748 152454 374776 460158
rect 374840 262886 374868 479538
rect 374920 475448 374972 475454
rect 374920 475390 374972 475396
rect 374828 262880 374880 262886
rect 374828 262822 374880 262828
rect 374932 262750 374960 475390
rect 375104 469056 375156 469062
rect 375104 468998 375156 469004
rect 375012 465928 375064 465934
rect 375012 465870 375064 465876
rect 375024 264586 375052 465870
rect 375116 373590 375144 468998
rect 375748 461780 375800 461786
rect 375748 461722 375800 461728
rect 375194 373960 375250 373969
rect 375194 373895 375250 373904
rect 375104 373584 375156 373590
rect 375104 373526 375156 373532
rect 375104 372564 375156 372570
rect 375104 372506 375156 372512
rect 375116 371618 375144 372506
rect 375104 371612 375156 371618
rect 375104 371554 375156 371560
rect 375012 264580 375064 264586
rect 375012 264522 375064 264528
rect 374920 262744 374972 262750
rect 374920 262686 374972 262692
rect 374920 262132 374972 262138
rect 374920 262074 374972 262080
rect 374828 243636 374880 243642
rect 374828 243578 374880 243584
rect 374736 152448 374788 152454
rect 374736 152390 374788 152396
rect 374552 150952 374604 150958
rect 374552 150894 374604 150900
rect 374840 133686 374868 243578
rect 374932 150822 374960 262074
rect 375012 260840 375064 260846
rect 375012 260782 375064 260788
rect 374920 150816 374972 150822
rect 374920 150758 374972 150764
rect 374828 133680 374880 133686
rect 374828 133622 374880 133628
rect 374840 132530 374868 133622
rect 374828 132524 374880 132530
rect 374828 132466 374880 132472
rect 374736 130484 374788 130490
rect 374736 130426 374788 130432
rect 374644 129804 374696 129810
rect 374644 129746 374696 129752
rect 374656 44606 374684 129746
rect 374644 44600 374696 44606
rect 374644 44542 374696 44548
rect 374748 44062 374776 130426
rect 374828 130348 374880 130354
rect 374828 130290 374880 130296
rect 374736 44056 374788 44062
rect 374736 43998 374788 44004
rect 374840 41002 374868 130290
rect 374932 44334 374960 150758
rect 375024 133822 375052 260782
rect 375116 240854 375144 371554
rect 375208 260846 375236 373895
rect 375286 372736 375342 372745
rect 375286 372671 375342 372680
rect 375196 260840 375248 260846
rect 375196 260782 375248 260788
rect 375196 241460 375248 241466
rect 375196 241402 375248 241408
rect 375104 240848 375156 240854
rect 375104 240790 375156 240796
rect 375012 133816 375064 133822
rect 375012 133758 375064 133764
rect 374920 44328 374972 44334
rect 374920 44270 374972 44276
rect 374828 40996 374880 41002
rect 374828 40938 374880 40944
rect 374460 39908 374512 39914
rect 374460 39850 374512 39856
rect 373816 39840 373868 39846
rect 373816 39782 373868 39788
rect 372436 39500 372488 39506
rect 372436 39442 372488 39448
rect 375024 39438 375052 133758
rect 375116 130150 375144 240790
rect 375208 240514 375236 241402
rect 375196 240508 375248 240514
rect 375196 240450 375248 240456
rect 375208 150890 375236 240450
rect 375300 240038 375328 372671
rect 375760 369714 375788 461722
rect 375748 369708 375800 369714
rect 375748 369650 375800 369656
rect 375840 369232 375892 369238
rect 375840 369174 375892 369180
rect 375852 262138 375880 369174
rect 375932 369164 375984 369170
rect 375932 369106 375984 369112
rect 375840 262132 375892 262138
rect 375840 262074 375892 262080
rect 375852 261594 375880 262074
rect 375840 261588 375892 261594
rect 375840 261530 375892 261536
rect 375944 260846 375972 369106
rect 375932 260840 375984 260846
rect 375932 260782 375984 260788
rect 375748 241460 375800 241466
rect 375748 241402 375800 241408
rect 375656 240780 375708 240786
rect 375656 240722 375708 240728
rect 375288 240032 375340 240038
rect 375288 239974 375340 239980
rect 375300 238814 375328 239974
rect 375288 238808 375340 238814
rect 375288 238750 375340 238756
rect 375288 151156 375340 151162
rect 375288 151098 375340 151104
rect 375196 150884 375248 150890
rect 375196 150826 375248 150832
rect 375196 133204 375248 133210
rect 375196 133146 375248 133152
rect 375104 130144 375156 130150
rect 375104 130086 375156 130092
rect 375208 40050 375236 133146
rect 375196 40044 375248 40050
rect 375196 39986 375248 39992
rect 375300 39778 375328 151098
rect 375668 130082 375696 240722
rect 375760 130558 375788 241402
rect 375838 239864 375894 239873
rect 375838 239799 375894 239808
rect 375852 151638 375880 239799
rect 375932 239284 375984 239290
rect 375932 239226 375984 239232
rect 375944 151774 375972 239226
rect 375932 151768 375984 151774
rect 375932 151710 375984 151716
rect 375840 151632 375892 151638
rect 375840 151574 375892 151580
rect 375748 130552 375800 130558
rect 375748 130494 375800 130500
rect 375656 130076 375708 130082
rect 375656 130018 375708 130024
rect 375668 129810 375696 130018
rect 375656 129804 375708 129810
rect 375656 129746 375708 129752
rect 375760 128722 375788 130494
rect 375748 128716 375800 128722
rect 375748 128658 375800 128664
rect 375852 43790 375880 151574
rect 375944 150550 375972 151710
rect 375932 150544 375984 150550
rect 375932 150486 375984 150492
rect 375932 129804 375984 129810
rect 375932 129746 375984 129752
rect 375840 43784 375892 43790
rect 375840 43726 375892 43732
rect 375944 43314 375972 129746
rect 376036 53145 376064 490554
rect 376128 153066 376156 490622
rect 376208 489184 376260 489190
rect 376208 489126 376260 489132
rect 376116 153060 376168 153066
rect 376116 153002 376168 153008
rect 376220 152522 376248 489126
rect 376760 481160 376812 481166
rect 376760 481102 376812 481108
rect 376484 477216 376536 477222
rect 376484 477158 376536 477164
rect 376300 468648 376352 468654
rect 376300 468590 376352 468596
rect 376312 262138 376340 468590
rect 376392 465860 376444 465866
rect 376392 465802 376444 465808
rect 376404 263129 376432 465802
rect 376496 369510 376524 477158
rect 376576 466336 376628 466342
rect 376576 466278 376628 466284
rect 376588 372570 376616 466278
rect 376576 372564 376628 372570
rect 376576 372506 376628 372512
rect 376772 372502 376800 481102
rect 377404 479664 377456 479670
rect 377404 479606 377456 479612
rect 377220 477012 377272 477018
rect 377220 476954 377272 476960
rect 377034 407824 377090 407833
rect 377034 407759 377090 407768
rect 376944 385008 376996 385014
rect 376942 384976 376944 384985
rect 376996 384976 376998 384985
rect 376942 384911 376998 384920
rect 376944 383648 376996 383654
rect 376944 383590 376996 383596
rect 376852 383580 376904 383586
rect 376852 383522 376904 383528
rect 376864 383081 376892 383522
rect 376956 383353 376984 383590
rect 376942 383344 376998 383353
rect 376942 383279 376998 383288
rect 376850 383072 376906 383081
rect 376850 383007 376906 383016
rect 376852 373788 376904 373794
rect 376852 373730 376904 373736
rect 376864 372638 376892 373730
rect 376852 372632 376904 372638
rect 376852 372574 376904 372580
rect 376760 372496 376812 372502
rect 376760 372438 376812 372444
rect 376760 372088 376812 372094
rect 376760 372030 376812 372036
rect 376772 371482 376800 372030
rect 376760 371476 376812 371482
rect 376760 371418 376812 371424
rect 376668 370388 376720 370394
rect 376668 370330 376720 370336
rect 376484 369504 376536 369510
rect 376484 369446 376536 369452
rect 376496 369238 376524 369446
rect 376484 369232 376536 369238
rect 376484 369174 376536 369180
rect 376576 368484 376628 368490
rect 376576 368426 376628 368432
rect 376484 368008 376536 368014
rect 376484 367950 376536 367956
rect 376390 263120 376446 263129
rect 376390 263055 376446 263064
rect 376300 262132 376352 262138
rect 376300 262074 376352 262080
rect 376392 262064 376444 262070
rect 376392 262006 376444 262012
rect 376300 261996 376352 262002
rect 376300 261938 376352 261944
rect 376312 260982 376340 261938
rect 376300 260976 376352 260982
rect 376300 260918 376352 260924
rect 376208 152516 376260 152522
rect 376208 152458 376260 152464
rect 376312 151298 376340 260918
rect 376404 260914 376432 262006
rect 376392 260908 376444 260914
rect 376392 260850 376444 260856
rect 376404 151570 376432 260850
rect 376496 241466 376524 367950
rect 376484 241460 376536 241466
rect 376484 241402 376536 241408
rect 376484 241324 376536 241330
rect 376484 241266 376536 241272
rect 376392 151564 376444 151570
rect 376392 151506 376444 151512
rect 376300 151292 376352 151298
rect 376300 151234 376352 151240
rect 376208 150476 376260 150482
rect 376208 150418 376260 150424
rect 376116 129736 376168 129742
rect 376116 129678 376168 129684
rect 376022 53136 376078 53145
rect 376022 53071 376078 53080
rect 375932 43308 375984 43314
rect 375932 43250 375984 43256
rect 376128 41342 376156 129678
rect 376220 44402 376248 150418
rect 376208 44396 376260 44402
rect 376208 44338 376260 44344
rect 376312 43926 376340 151234
rect 376404 150482 376432 151506
rect 376392 150476 376444 150482
rect 376392 150418 376444 150424
rect 376496 130830 376524 241266
rect 376588 240106 376616 368426
rect 376680 241058 376708 370330
rect 377048 306374 377076 407759
rect 377128 370728 377180 370734
rect 377128 370670 377180 370676
rect 377140 370530 377168 370670
rect 377128 370524 377180 370530
rect 377128 370466 377180 370472
rect 377140 370433 377168 370466
rect 377126 370424 377182 370433
rect 377126 370359 377182 370368
rect 377232 369442 377260 476954
rect 377310 410000 377366 410009
rect 377310 409935 377366 409944
rect 377220 369436 377272 369442
rect 377220 369378 377272 369384
rect 377324 306374 377352 409935
rect 377416 407833 377444 479606
rect 377680 471640 377732 471646
rect 377680 471582 377732 471588
rect 377496 471436 377548 471442
rect 377496 471378 377548 471384
rect 377402 407824 377458 407833
rect 377402 407759 377458 407768
rect 377404 406428 377456 406434
rect 377404 406370 377456 406376
rect 377416 406065 377444 406370
rect 377402 406056 377458 406065
rect 377402 405991 377458 406000
rect 377508 374406 377536 471378
rect 377588 464364 377640 464370
rect 377588 464306 377640 464312
rect 377600 411913 377628 464306
rect 377586 411904 377642 411913
rect 377586 411839 377642 411848
rect 377496 374400 377548 374406
rect 377496 374342 377548 374348
rect 377496 370320 377548 370326
rect 377496 370262 377548 370268
rect 377048 306346 377260 306374
rect 377324 306346 377444 306374
rect 377232 302002 377260 306346
rect 377232 301974 377352 302002
rect 377218 301880 377274 301889
rect 377218 301815 377274 301824
rect 376850 300928 376906 300937
rect 376850 300863 376906 300872
rect 376758 295352 376814 295361
rect 376758 295287 376814 295296
rect 376772 274802 376800 295287
rect 376864 276162 376892 300863
rect 376942 298752 376998 298761
rect 376942 298687 376998 298696
rect 376956 276282 376984 298687
rect 377126 293992 377182 294001
rect 377126 293927 377182 293936
rect 376944 276276 376996 276282
rect 376944 276218 376996 276224
rect 376864 276134 377076 276162
rect 376944 276072 376996 276078
rect 376944 276014 376996 276020
rect 376852 276004 376904 276010
rect 376852 275946 376904 275952
rect 376864 274961 376892 275946
rect 376850 274952 376906 274961
rect 376850 274887 376906 274896
rect 376772 274774 376892 274802
rect 376760 274644 376812 274650
rect 376760 274586 376812 274592
rect 376772 273329 376800 274586
rect 376758 273320 376814 273329
rect 376758 273255 376814 273264
rect 376760 273216 376812 273222
rect 376760 273158 376812 273164
rect 376772 273057 376800 273158
rect 376758 273048 376814 273057
rect 376758 272983 376814 272992
rect 376864 272626 376892 274774
rect 376772 272598 376892 272626
rect 376668 241052 376720 241058
rect 376668 240994 376720 241000
rect 376680 240786 376708 240994
rect 376668 240780 376720 240786
rect 376668 240722 376720 240728
rect 376576 240100 376628 240106
rect 376576 240042 376628 240048
rect 376588 239290 376616 240042
rect 376576 239284 376628 239290
rect 376576 239226 376628 239232
rect 376772 185994 376800 272598
rect 376852 272536 376904 272542
rect 376852 272478 376904 272484
rect 376864 191729 376892 272478
rect 376850 191720 376906 191729
rect 376850 191655 376906 191664
rect 376956 188737 376984 276014
rect 377048 272542 377076 276134
rect 377036 272536 377088 272542
rect 377036 272478 377088 272484
rect 377036 260840 377088 260846
rect 377036 260782 377088 260788
rect 377048 260234 377076 260782
rect 377036 260228 377088 260234
rect 377036 260170 377088 260176
rect 376942 188728 376998 188737
rect 376942 188663 376998 188672
rect 376956 187921 376984 188663
rect 376942 187912 376998 187921
rect 376942 187847 376998 187856
rect 376942 186008 376998 186017
rect 376772 185966 376942 185994
rect 376942 185943 376998 185952
rect 376956 171134 376984 185943
rect 376864 171106 376984 171134
rect 376760 164212 376812 164218
rect 376760 164154 376812 164160
rect 376772 163169 376800 164154
rect 376758 163160 376814 163169
rect 376758 163095 376814 163104
rect 376864 161474 376892 171106
rect 376944 165572 376996 165578
rect 376944 165514 376996 165520
rect 376956 165073 376984 165514
rect 376942 165064 376998 165073
rect 376942 164999 376998 165008
rect 376944 163532 376996 163538
rect 376944 163474 376996 163480
rect 376956 163441 376984 163474
rect 376942 163432 376998 163441
rect 376942 163367 376998 163376
rect 376864 161446 376984 161474
rect 376668 150544 376720 150550
rect 376668 150486 376720 150492
rect 376484 130824 376536 130830
rect 376484 130766 376536 130772
rect 376392 129872 376444 129878
rect 376392 129814 376444 129820
rect 376404 44130 376432 129814
rect 376496 129810 376524 130766
rect 376574 130384 376630 130393
rect 376574 130319 376630 130328
rect 376484 129804 376536 129810
rect 376484 129746 376536 129752
rect 376588 129742 376616 130319
rect 376576 129736 376628 129742
rect 376576 129678 376628 129684
rect 376576 128716 376628 128722
rect 376576 128658 376628 128664
rect 376392 44124 376444 44130
rect 376392 44066 376444 44072
rect 376300 43920 376352 43926
rect 376300 43862 376352 43868
rect 376116 41336 376168 41342
rect 376116 41278 376168 41284
rect 375288 39772 375340 39778
rect 375288 39714 375340 39720
rect 376588 39574 376616 128658
rect 376680 39982 376708 150486
rect 376956 76129 376984 161446
rect 377048 150550 377076 260170
rect 377140 185065 377168 293927
rect 377232 193225 377260 301815
rect 377324 297809 377352 301974
rect 377416 300937 377444 306346
rect 377402 300928 377458 300937
rect 377402 300863 377458 300872
rect 377310 297800 377366 297809
rect 377310 297735 377366 297744
rect 377218 193216 377274 193225
rect 377218 193151 377274 193160
rect 377218 187912 377274 187921
rect 377218 187847 377274 187856
rect 377126 185056 377182 185065
rect 377126 184991 377182 185000
rect 377036 150544 377088 150550
rect 377036 150486 377088 150492
rect 376942 76120 376998 76129
rect 376942 76055 376998 76064
rect 377140 75041 377168 184991
rect 377232 180794 377260 187847
rect 377324 187785 377352 297735
rect 377508 241330 377536 370262
rect 377600 301889 377628 411839
rect 377692 408762 377720 471582
rect 377772 470076 377824 470082
rect 377772 470018 377824 470024
rect 377784 410961 377812 470018
rect 378152 468518 378180 535078
rect 383672 532370 383700 535078
rect 387904 532438 387932 535078
rect 387892 532432 387944 532438
rect 387892 532374 387944 532380
rect 383660 532364 383712 532370
rect 383660 532306 383712 532312
rect 379980 483744 380032 483750
rect 379980 483686 380032 483692
rect 378876 483676 378928 483682
rect 378876 483618 378928 483624
rect 378784 476808 378836 476814
rect 378784 476750 378836 476756
rect 378140 468512 378192 468518
rect 378140 468454 378192 468460
rect 377770 410952 377826 410961
rect 377770 410887 377826 410896
rect 377784 410009 377812 410887
rect 377770 410000 377826 410009
rect 377770 409935 377826 409944
rect 377862 408776 377918 408785
rect 377692 408734 377862 408762
rect 377862 408711 377918 408720
rect 377680 405000 377732 405006
rect 377678 404968 377680 404977
rect 377732 404968 377734 404977
rect 377678 404903 377734 404912
rect 377586 301880 377642 301889
rect 377586 301815 377642 301824
rect 377692 294953 377720 404903
rect 377772 403640 377824 403646
rect 377772 403582 377824 403588
rect 377784 403209 377812 403582
rect 377770 403200 377826 403209
rect 377770 403135 377826 403144
rect 377678 294944 377734 294953
rect 377678 294879 377734 294888
rect 377692 294001 377720 294879
rect 377678 293992 377734 294001
rect 377678 293927 377734 293936
rect 377784 293185 377812 403135
rect 377876 298761 377904 408711
rect 377954 406056 378010 406065
rect 377954 405991 378010 406000
rect 377968 402974 377996 405991
rect 377968 402946 378088 402974
rect 378060 379514 378088 402946
rect 377968 379486 378088 379514
rect 377862 298752 377918 298761
rect 377862 298687 377918 298696
rect 377968 296041 377996 379486
rect 378046 372736 378102 372745
rect 378046 372671 378102 372680
rect 378060 372638 378088 372671
rect 378048 372632 378100 372638
rect 378048 372574 378100 372580
rect 378048 371476 378100 371482
rect 378048 371418 378100 371424
rect 377954 296032 378010 296041
rect 377954 295967 378010 295976
rect 377968 295361 377996 295967
rect 377954 295352 378010 295361
rect 377954 295287 378010 295296
rect 377770 293176 377826 293185
rect 377770 293111 377826 293120
rect 377496 241324 377548 241330
rect 377496 241266 377548 241272
rect 377508 240990 377536 241266
rect 377588 241256 377640 241262
rect 377588 241198 377640 241204
rect 377496 240984 377548 240990
rect 377496 240926 377548 240932
rect 377310 187776 377366 187785
rect 377310 187711 377366 187720
rect 377494 183560 377550 183569
rect 377494 183495 377550 183504
rect 377232 180766 377352 180794
rect 377218 129840 377274 129849
rect 377218 129775 377274 129784
rect 377126 75032 377182 75041
rect 377126 74967 377182 74976
rect 376944 55208 376996 55214
rect 376944 55150 376996 55156
rect 376956 55049 376984 55150
rect 376942 55040 376998 55049
rect 376942 54975 376998 54984
rect 376942 53272 376998 53281
rect 376942 53207 376998 53216
rect 376956 53106 376984 53207
rect 376944 53100 376996 53106
rect 376944 53042 376996 53048
rect 377232 44470 377260 129775
rect 377324 78849 377352 180766
rect 377310 78840 377366 78849
rect 377310 78775 377366 78784
rect 377508 73273 377536 183495
rect 377600 131034 377628 241198
rect 377680 241120 377732 241126
rect 377680 241062 377732 241068
rect 377692 151814 377720 241062
rect 377784 183569 377812 293111
rect 378060 241398 378088 371418
rect 378692 369436 378744 369442
rect 378692 369378 378744 369384
rect 378600 349580 378652 349586
rect 378600 349522 378652 349528
rect 378506 262984 378562 262993
rect 378506 262919 378562 262928
rect 378048 241392 378100 241398
rect 378048 241334 378100 241340
rect 378048 239964 378100 239970
rect 378048 239906 378100 239912
rect 378060 239873 378088 239906
rect 378046 239864 378102 239873
rect 378046 239799 378102 239808
rect 377954 193216 378010 193225
rect 377954 193151 378010 193160
rect 377968 191865 377996 193151
rect 377954 191856 378010 191865
rect 377954 191791 378010 191800
rect 377862 191720 377918 191729
rect 377862 191655 377918 191664
rect 377876 190913 377904 191655
rect 377862 190904 377918 190913
rect 377862 190839 377918 190848
rect 377770 183560 377826 183569
rect 377770 183495 377826 183504
rect 377772 165164 377824 165170
rect 377772 165106 377824 165112
rect 377784 156670 377812 165106
rect 377772 156664 377824 156670
rect 377772 156606 377824 156612
rect 377692 151786 377812 151814
rect 377678 133784 377734 133793
rect 377678 133719 377734 133728
rect 377692 133550 377720 133719
rect 377680 133544 377732 133550
rect 377680 133486 377732 133492
rect 377784 132494 377812 151786
rect 377692 132466 377812 132494
rect 377588 131028 377640 131034
rect 377588 130970 377640 130976
rect 377494 73264 377550 73273
rect 377494 73199 377550 73208
rect 377220 44464 377272 44470
rect 377220 44406 377272 44412
rect 376668 39976 376720 39982
rect 376668 39918 376720 39924
rect 377600 39710 377628 130970
rect 377692 130898 377720 132466
rect 377680 130892 377732 130898
rect 377680 130834 377732 130840
rect 377692 41138 377720 130834
rect 377876 81025 377904 190839
rect 377968 165170 377996 191791
rect 378046 187776 378102 187785
rect 378046 187711 378102 187720
rect 377956 165164 378008 165170
rect 377956 165106 378008 165112
rect 377956 156664 378008 156670
rect 377956 156606 378008 156612
rect 377968 81977 377996 156606
rect 377954 81968 378010 81977
rect 377954 81903 378010 81912
rect 377862 81016 377918 81025
rect 377862 80951 377918 80960
rect 378060 77897 378088 187711
rect 378046 77888 378102 77897
rect 378046 77823 378102 77832
rect 378520 42770 378548 262919
rect 378612 262070 378640 349522
rect 378704 262274 378732 369378
rect 378692 262268 378744 262274
rect 378692 262210 378744 262216
rect 378600 262064 378652 262070
rect 378600 262006 378652 262012
rect 378600 241460 378652 241466
rect 378600 241402 378652 241408
rect 378612 133890 378640 241402
rect 378692 241392 378744 241398
rect 378692 241334 378744 241340
rect 378704 240854 378732 241334
rect 378692 240848 378744 240854
rect 378692 240790 378744 240796
rect 378600 133884 378652 133890
rect 378600 133826 378652 133832
rect 378704 130626 378732 240790
rect 378692 130620 378744 130626
rect 378692 130562 378744 130568
rect 378692 130280 378744 130286
rect 378692 130222 378744 130228
rect 378600 130212 378652 130218
rect 378600 130154 378652 130160
rect 378612 44674 378640 130154
rect 378704 44742 378732 130222
rect 378692 44736 378744 44742
rect 378692 44678 378744 44684
rect 378600 44668 378652 44674
rect 378600 44610 378652 44616
rect 378508 42764 378560 42770
rect 378508 42706 378560 42712
rect 378796 42226 378824 476750
rect 378888 152318 378916 483618
rect 379060 481024 379112 481030
rect 379060 480966 379112 480972
rect 378968 468580 379020 468586
rect 378968 468522 379020 468528
rect 378980 152833 379008 468522
rect 379072 262818 379100 480966
rect 379520 479800 379572 479806
rect 379520 479742 379572 479748
rect 379244 475516 379296 475522
rect 379244 475458 379296 475464
rect 379152 458856 379204 458862
rect 379152 458798 379204 458804
rect 379060 262812 379112 262818
rect 379060 262754 379112 262760
rect 379060 240916 379112 240922
rect 379060 240858 379112 240864
rect 378966 152824 379022 152833
rect 378966 152759 379022 152768
rect 378876 152312 378928 152318
rect 378876 152254 378928 152260
rect 379072 130694 379100 240858
rect 379164 152697 379192 458798
rect 379256 263265 379284 475458
rect 379428 460896 379480 460902
rect 379428 460838 379480 460844
rect 379336 460760 379388 460766
rect 379336 460702 379388 460708
rect 379348 372026 379376 460702
rect 379440 373794 379468 460838
rect 379532 383654 379560 479742
rect 379532 383626 379744 383654
rect 379428 373788 379480 373794
rect 379428 373730 379480 373736
rect 379612 372360 379664 372366
rect 379612 372302 379664 372308
rect 379520 372156 379572 372162
rect 379520 372098 379572 372104
rect 379336 372020 379388 372026
rect 379336 371962 379388 371968
rect 379348 371362 379376 371962
rect 379532 371550 379560 372098
rect 379624 371754 379652 372302
rect 379612 371748 379664 371754
rect 379612 371690 379664 371696
rect 379520 371544 379572 371550
rect 379520 371486 379572 371492
rect 379348 371334 379560 371362
rect 379336 369368 379388 369374
rect 379336 369310 379388 369316
rect 379242 263256 379298 263265
rect 379242 263191 379298 263200
rect 379244 262064 379296 262070
rect 379244 262006 379296 262012
rect 379150 152688 379206 152697
rect 379150 152623 379206 152632
rect 379256 151706 379284 262006
rect 379348 261050 379376 369310
rect 379428 367940 379480 367946
rect 379428 367882 379480 367888
rect 379336 261044 379388 261050
rect 379336 260986 379388 260992
rect 379244 151700 379296 151706
rect 379244 151642 379296 151648
rect 379256 150482 379284 151642
rect 379348 151026 379376 260986
rect 379440 260794 379468 367882
rect 379532 364334 379560 371334
rect 379612 370660 379664 370666
rect 379612 370602 379664 370608
rect 379624 369889 379652 370602
rect 379610 369880 379666 369889
rect 379610 369815 379666 369824
rect 379716 368490 379744 383626
rect 379796 371748 379848 371754
rect 379796 371690 379848 371696
rect 379704 368484 379756 368490
rect 379704 368426 379756 368432
rect 379808 368370 379836 371690
rect 379888 371544 379940 371550
rect 379888 371486 379940 371492
rect 379716 368342 379836 368370
rect 379532 364306 379652 364334
rect 379624 262002 379652 364306
rect 379612 261996 379664 262002
rect 379612 261938 379664 261944
rect 379440 260766 379652 260794
rect 379518 260672 379574 260681
rect 379518 260607 379574 260616
rect 379428 241324 379480 241330
rect 379428 241266 379480 241272
rect 379440 240786 379468 241266
rect 379428 240780 379480 240786
rect 379428 240722 379480 240728
rect 379532 151366 379560 260607
rect 379624 260166 379652 260766
rect 379612 260160 379664 260166
rect 379612 260102 379664 260108
rect 379520 151360 379572 151366
rect 379520 151302 379572 151308
rect 379336 151020 379388 151026
rect 379336 150962 379388 150968
rect 379244 150476 379296 150482
rect 379244 150418 379296 150424
rect 379348 142154 379376 150962
rect 379428 150476 379480 150482
rect 379428 150418 379480 150424
rect 379256 142126 379376 142154
rect 379152 133884 379204 133890
rect 379152 133826 379204 133832
rect 379164 133754 379192 133826
rect 379152 133748 379204 133754
rect 379152 133690 379204 133696
rect 379060 130688 379112 130694
rect 379060 130630 379112 130636
rect 378876 130144 378928 130150
rect 378876 130086 378928 130092
rect 378888 43382 378916 130086
rect 379072 129878 379100 130630
rect 379060 129872 379112 129878
rect 379060 129814 379112 129820
rect 378968 129804 379020 129810
rect 378968 129746 379020 129752
rect 378876 43376 378928 43382
rect 378876 43318 378928 43324
rect 378784 42220 378836 42226
rect 378784 42162 378836 42168
rect 378980 42022 379008 129746
rect 378968 42016 379020 42022
rect 378968 41958 379020 41964
rect 379164 41206 379192 133690
rect 379256 43994 379284 142126
rect 379336 133816 379388 133822
rect 379336 133758 379388 133764
rect 379348 133550 379376 133758
rect 379336 133544 379388 133550
rect 379336 133486 379388 133492
rect 379336 130960 379388 130966
rect 379336 130902 379388 130908
rect 379348 130626 379376 130902
rect 379336 130620 379388 130626
rect 379336 130562 379388 130568
rect 379244 43988 379296 43994
rect 379244 43930 379296 43936
rect 379152 41200 379204 41206
rect 379152 41142 379204 41148
rect 377680 41132 377732 41138
rect 377680 41074 377732 41080
rect 377588 39704 377640 39710
rect 377588 39646 377640 39652
rect 379348 39642 379376 130562
rect 379440 41274 379468 150418
rect 379624 131073 379652 260102
rect 379716 241126 379744 368342
rect 379796 368280 379848 368286
rect 379796 368222 379848 368228
rect 379808 241262 379836 368222
rect 379900 241466 379928 371486
rect 379992 371414 380020 483686
rect 391952 469878 391980 535078
rect 396920 532302 396948 535078
rect 396908 532296 396960 532302
rect 396908 532238 396960 532244
rect 401612 531826 401640 535078
rect 405936 533254 405964 535078
rect 405924 533248 405976 533254
rect 405924 533190 405976 533196
rect 410536 532506 410564 535078
rect 414952 533322 414980 535078
rect 414940 533316 414992 533322
rect 414940 533258 414992 533264
rect 410524 532500 410576 532506
rect 410524 532442 410576 532448
rect 419552 531962 419580 535078
rect 419540 531956 419592 531962
rect 419540 531898 419592 531904
rect 423968 531894 423996 535078
rect 423956 531888 424008 531894
rect 423956 531830 424008 531836
rect 401600 531820 401652 531826
rect 401600 531762 401652 531768
rect 428384 531214 428412 573271
rect 428462 563816 428518 563825
rect 428462 563751 428518 563760
rect 428476 534750 428504 563751
rect 428554 535936 428610 535945
rect 428554 535871 428610 535880
rect 428464 534744 428516 534750
rect 428464 534686 428516 534692
rect 428372 531208 428424 531214
rect 428372 531150 428424 531156
rect 428568 529786 428596 535871
rect 428556 529780 428608 529786
rect 428556 529722 428608 529728
rect 429212 471986 429240 598295
rect 429304 545329 429332 650626
rect 430580 649324 430632 649330
rect 430580 649266 430632 649272
rect 429936 646604 429988 646610
rect 429936 646546 429988 646552
rect 429844 646400 429896 646406
rect 429844 646342 429896 646348
rect 429856 626550 429884 646342
rect 429948 636954 429976 646546
rect 430592 641209 430620 649266
rect 430672 648780 430724 648786
rect 430672 648722 430724 648728
rect 430578 641200 430634 641209
rect 430578 641135 430634 641144
rect 429936 636948 429988 636954
rect 429936 636890 429988 636896
rect 430684 631689 430712 648722
rect 430854 647320 430910 647329
rect 430854 647255 430910 647264
rect 430764 646264 430816 646270
rect 430764 646206 430816 646212
rect 430776 636449 430804 646206
rect 430762 636440 430818 636449
rect 430762 636375 430818 636384
rect 430670 631680 430726 631689
rect 430670 631615 430726 631624
rect 430868 626929 430896 647255
rect 432604 646536 432656 646542
rect 432604 646478 432656 646484
rect 432616 636886 432644 646478
rect 432604 636880 432656 636886
rect 432604 636822 432656 636828
rect 430854 626920 430910 626929
rect 430854 626855 430910 626864
rect 429844 626544 429896 626550
rect 429844 626486 429896 626492
rect 430578 617400 430634 617409
rect 430578 617335 430634 617344
rect 429382 593600 429438 593609
rect 429382 593535 429438 593544
rect 429290 545320 429346 545329
rect 429290 545255 429346 545264
rect 429396 529854 429424 593535
rect 429474 588160 429530 588169
rect 429474 588095 429530 588104
rect 429488 535022 429516 588095
rect 430592 542858 430620 617335
rect 430670 612640 430726 612649
rect 430670 612575 430726 612584
rect 430684 542994 430712 612575
rect 430762 603120 430818 603129
rect 430762 603055 430818 603064
rect 430776 543114 430804 603055
rect 430854 583400 430910 583409
rect 430854 583335 430910 583344
rect 430764 543108 430816 543114
rect 430764 543050 430816 543056
rect 430684 542966 430804 542994
rect 430592 542830 430712 542858
rect 430578 540560 430634 540569
rect 430578 540495 430634 540504
rect 429476 535016 429528 535022
rect 429476 534958 429528 534964
rect 430592 534954 430620 540495
rect 430684 535226 430712 542830
rect 430672 535220 430724 535226
rect 430672 535162 430724 535168
rect 430776 535158 430804 542966
rect 430764 535152 430816 535158
rect 430764 535094 430816 535100
rect 430580 534948 430632 534954
rect 430580 534890 430632 534896
rect 430868 533526 430896 583335
rect 430946 578640 431002 578649
rect 430946 578575 431002 578584
rect 430960 543250 430988 578575
rect 431038 569120 431094 569129
rect 431038 569055 431094 569064
rect 430948 543244 431000 543250
rect 430948 543186 431000 543192
rect 430948 543108 431000 543114
rect 430948 543050 431000 543056
rect 430856 533520 430908 533526
rect 430856 533462 430908 533468
rect 430960 533390 430988 543050
rect 431052 533594 431080 569055
rect 431130 559600 431186 559609
rect 431130 559535 431186 559544
rect 431144 534818 431172 559535
rect 431222 554840 431278 554849
rect 431222 554775 431278 554784
rect 431236 534886 431264 554775
rect 431314 550080 431370 550089
rect 431314 550015 431370 550024
rect 431328 535090 431356 550015
rect 431408 543244 431460 543250
rect 431408 543186 431460 543192
rect 431316 535084 431368 535090
rect 431316 535026 431368 535032
rect 431224 534880 431276 534886
rect 431224 534822 431276 534828
rect 431132 534812 431184 534818
rect 431132 534754 431184 534760
rect 431040 533588 431092 533594
rect 431040 533530 431092 533536
rect 431420 533458 431448 543186
rect 436756 534041 436784 699654
rect 498212 652050 498240 703582
rect 499224 703474 499252 703582
rect 499366 703520 499478 704960
rect 514730 703520 514842 704960
rect 530094 703520 530206 704960
rect 545458 703520 545570 704960
rect 560822 703520 560934 704960
rect 576186 703520 576298 704960
rect 499408 703474 499436 703520
rect 499224 703446 499436 703474
rect 530136 701010 530164 703520
rect 530124 701004 530176 701010
rect 530124 700946 530176 700952
rect 531228 701004 531280 701010
rect 531228 700946 531280 700952
rect 531240 700330 531268 700946
rect 531228 700324 531280 700330
rect 531228 700266 531280 700272
rect 545500 697610 545528 703520
rect 580264 700324 580316 700330
rect 580264 700266 580316 700272
rect 545488 697604 545540 697610
rect 545488 697546 545540 697552
rect 580276 671945 580304 700266
rect 580262 671936 580318 671945
rect 580262 671871 580318 671880
rect 580276 670721 580304 671871
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580906 670712 580962 670721
rect 580906 670647 580962 670656
rect 579894 659152 579950 659161
rect 579894 659087 579950 659096
rect 579908 658306 579936 659087
rect 579896 658300 579948 658306
rect 579896 658242 579948 658248
rect 498200 652044 498252 652050
rect 498200 651986 498252 651992
rect 457444 650072 457496 650078
rect 457444 650014 457496 650020
rect 456800 634772 456852 634778
rect 456800 634714 456852 634720
rect 456812 634681 456840 634714
rect 456798 634672 456854 634681
rect 456798 634607 456854 634616
rect 456800 626544 456852 626550
rect 456800 626486 456852 626492
rect 456812 626385 456840 626486
rect 456798 626376 456854 626385
rect 456798 626311 456854 626320
rect 457456 618225 457484 650014
rect 489920 648712 489972 648718
rect 489920 648654 489972 648660
rect 466736 646332 466788 646338
rect 466736 646274 466788 646280
rect 466748 634930 466776 646274
rect 474740 636948 474792 636954
rect 474740 636890 474792 636896
rect 474752 634930 474780 636890
rect 482928 636268 482980 636274
rect 482928 636210 482980 636216
rect 482940 634930 482968 636210
rect 466748 634902 467130 634930
rect 474752 634902 474858 634930
rect 482586 634902 482968 634930
rect 489932 634930 489960 648654
rect 580264 648644 580316 648650
rect 580264 648586 580316 648592
rect 497648 646196 497700 646202
rect 497648 646138 497700 646144
rect 497660 634930 497688 646138
rect 512000 646128 512052 646134
rect 512000 646070 512052 646076
rect 510620 646060 510672 646066
rect 510620 646002 510672 646008
rect 505468 636880 505520 636886
rect 505468 636822 505520 636828
rect 505480 634930 505508 636822
rect 489932 634902 490314 634930
rect 497660 634902 498042 634930
rect 505480 634902 505770 634930
rect 510632 623121 510660 646002
rect 511356 636268 511408 636274
rect 511356 636210 511408 636216
rect 510618 623112 510674 623121
rect 510618 623047 510674 623056
rect 457442 618216 457498 618225
rect 457442 618151 457498 618160
rect 457442 608968 457498 608977
rect 457442 608903 457498 608912
rect 436742 534032 436798 534041
rect 436742 533967 436798 533976
rect 457456 533662 457484 608903
rect 457534 600808 457590 600817
rect 457534 600743 457590 600752
rect 457548 533730 457576 600743
rect 511262 597680 511318 597689
rect 511262 597615 511318 597624
rect 457626 592648 457682 592657
rect 457626 592583 457682 592592
rect 457640 533866 457668 592583
rect 459572 585126 460046 585154
rect 466472 585126 467774 585154
rect 474752 585126 475502 585154
rect 483032 585126 483230 585154
rect 489932 585126 490958 585154
rect 498212 585126 498686 585154
rect 505112 585126 506414 585154
rect 457628 533860 457680 533866
rect 457628 533802 457680 533808
rect 459572 533798 459600 585126
rect 466472 535294 466500 585126
rect 466460 535288 466512 535294
rect 466460 535230 466512 535236
rect 459560 533792 459612 533798
rect 459560 533734 459612 533740
rect 457536 533724 457588 533730
rect 457536 533666 457588 533672
rect 457444 533656 457496 533662
rect 457444 533598 457496 533604
rect 431408 533452 431460 533458
rect 431408 533394 431460 533400
rect 430948 533384 431000 533390
rect 430948 533326 431000 533332
rect 474752 531282 474780 585126
rect 483032 533934 483060 585126
rect 489932 534002 489960 585126
rect 489920 533996 489972 534002
rect 489920 533938 489972 533944
rect 483020 533928 483072 533934
rect 483020 533870 483072 533876
rect 474740 531276 474792 531282
rect 474740 531218 474792 531224
rect 429384 529848 429436 529854
rect 429384 529790 429436 529796
rect 498212 494018 498240 585126
rect 505112 535362 505140 585126
rect 505100 535356 505152 535362
rect 505100 535298 505152 535304
rect 498200 494012 498252 494018
rect 498200 493954 498252 493960
rect 429200 471980 429252 471986
rect 429200 471922 429252 471928
rect 391940 469872 391992 469878
rect 391940 469814 391992 469820
rect 511276 462233 511304 597615
rect 511368 557530 511396 636210
rect 512012 630601 512040 646070
rect 511998 630592 512054 630601
rect 511998 630527 512054 630536
rect 511998 614136 512054 614145
rect 511998 614071 512054 614080
rect 511356 557524 511408 557530
rect 511356 557466 511408 557472
rect 512012 529922 512040 614071
rect 580276 608025 580304 648586
rect 580920 620809 580948 670647
rect 580906 620800 580962 620809
rect 580906 620735 580962 620744
rect 580262 608016 580318 608025
rect 580262 607951 580318 607960
rect 512090 605976 512146 605985
rect 512090 605911 512146 605920
rect 512104 534070 512132 605911
rect 512182 589384 512238 589393
rect 512182 589319 512238 589328
rect 512196 535430 512224 589319
rect 580920 569537 580948 620735
rect 580906 569528 580962 569537
rect 580906 569463 580962 569472
rect 580172 557524 580224 557530
rect 580172 557466 580224 557472
rect 580184 556753 580212 557466
rect 580170 556744 580226 556753
rect 580170 556679 580226 556688
rect 512184 535424 512236 535430
rect 512184 535366 512236 535372
rect 512092 534064 512144 534070
rect 512092 534006 512144 534012
rect 518164 530596 518216 530602
rect 518164 530538 518216 530544
rect 512000 529916 512052 529922
rect 512000 529858 512052 529864
rect 511262 462224 511318 462233
rect 511262 462159 511318 462168
rect 511276 461922 511304 462159
rect 511264 461916 511316 461922
rect 511264 461858 511316 461864
rect 517520 461916 517572 461922
rect 517520 461858 517572 461864
rect 499856 461100 499908 461106
rect 499856 461042 499908 461048
rect 500868 461100 500920 461106
rect 500868 461042 500920 461048
rect 498476 461032 498528 461038
rect 498474 461000 498476 461009
rect 499868 461009 499896 461042
rect 498528 461000 498530 461009
rect 498474 460935 498530 460944
rect 499854 461000 499910 461009
rect 500880 460970 500908 461042
rect 499854 460935 499910 460944
rect 500868 460964 500920 460970
rect 500868 460906 500920 460912
rect 516600 458312 516652 458318
rect 516600 458254 516652 458260
rect 516612 454753 516640 458254
rect 516598 454744 516654 454753
rect 516598 454679 516654 454688
rect 407762 375048 407818 375057
rect 407762 374983 407818 374992
rect 418250 375048 418306 375057
rect 418250 374983 418306 374992
rect 440330 375048 440386 375057
rect 440330 374983 440386 374992
rect 443090 375048 443146 375057
rect 443090 374983 443146 374992
rect 407776 374610 407804 374983
rect 418264 374678 418292 374983
rect 440344 374814 440372 374983
rect 440332 374808 440384 374814
rect 440332 374750 440384 374756
rect 418252 374672 418304 374678
rect 410706 374640 410762 374649
rect 407764 374604 407816 374610
rect 418252 374614 418304 374620
rect 410706 374575 410762 374584
rect 407764 374546 407816 374552
rect 410720 374542 410748 374575
rect 410708 374536 410760 374542
rect 410708 374478 410760 374484
rect 433338 374504 433394 374513
rect 433338 374439 433340 374448
rect 433392 374439 433394 374448
rect 433614 374504 433670 374513
rect 433614 374439 433670 374448
rect 433340 374410 433392 374416
rect 433628 374270 433656 374439
rect 443104 374406 443132 374983
rect 445942 374504 445998 374513
rect 445942 374439 445998 374448
rect 448242 374504 448298 374513
rect 448242 374439 448298 374448
rect 443092 374400 443144 374406
rect 443092 374342 443144 374348
rect 434812 374332 434864 374338
rect 434812 374274 434864 374280
rect 433616 374264 433668 374270
rect 415674 374232 415730 374241
rect 434824 374241 434852 374274
rect 433616 374206 433668 374212
rect 434810 374232 434866 374241
rect 415674 374167 415730 374176
rect 445956 374202 445984 374439
rect 434810 374167 434866 374176
rect 445944 374196 445996 374202
rect 404820 373992 404872 373998
rect 404820 373934 404872 373940
rect 404832 373833 404860 373934
rect 404818 373824 404874 373833
rect 404818 373759 404874 373768
rect 380900 373244 380952 373250
rect 380900 373186 380952 373192
rect 380912 372706 380940 373186
rect 380900 372700 380952 372706
rect 380900 372642 380952 372648
rect 380072 371680 380124 371686
rect 380072 371622 380124 371628
rect 379980 371408 380032 371414
rect 379980 371350 380032 371356
rect 380084 368286 380112 371622
rect 380072 368280 380124 368286
rect 380072 368222 380124 368228
rect 380912 349586 380940 372642
rect 405738 372192 405794 372201
rect 405738 372127 405794 372136
rect 396078 372056 396134 372065
rect 396078 371991 396080 372000
rect 396132 371991 396134 372000
rect 398838 372056 398894 372065
rect 398838 371991 398894 372000
rect 396080 371962 396132 371968
rect 398852 371958 398880 371991
rect 398840 371952 398892 371958
rect 397458 371920 397514 371929
rect 398840 371894 398892 371900
rect 405752 371890 405780 372127
rect 412822 371920 412878 371929
rect 397458 371855 397514 371864
rect 405740 371884 405792 371890
rect 397472 371822 397500 371855
rect 412822 371855 412878 371864
rect 405740 371826 405792 371832
rect 397460 371816 397512 371822
rect 397460 371758 397512 371764
rect 409878 371784 409934 371793
rect 409878 371719 409880 371728
rect 409932 371719 409934 371728
rect 411258 371784 411314 371793
rect 411258 371719 411314 371728
rect 409880 371690 409932 371696
rect 411272 371686 411300 371719
rect 411260 371680 411312 371686
rect 407118 371648 407174 371657
rect 411260 371622 411312 371628
rect 412638 371648 412694 371657
rect 407118 371583 407120 371592
rect 407172 371583 407174 371592
rect 412638 371583 412694 371592
rect 407120 371554 407172 371560
rect 412652 371550 412680 371583
rect 412640 371544 412692 371550
rect 411258 371512 411314 371521
rect 412640 371486 412692 371492
rect 411258 371447 411260 371456
rect 411312 371447 411314 371456
rect 411260 371418 411312 371424
rect 380992 371408 381044 371414
rect 380992 371350 381044 371356
rect 396078 371376 396134 371385
rect 381004 349761 381032 371350
rect 396078 371311 396134 371320
rect 402978 371376 403034 371385
rect 402978 371311 403034 371320
rect 403254 371376 403310 371385
rect 403254 371311 403310 371320
rect 408498 371376 408554 371385
rect 408498 371311 408554 371320
rect 396092 370598 396120 371311
rect 396080 370592 396132 370598
rect 396080 370534 396132 370540
rect 402992 370530 403020 371311
rect 402980 370524 403032 370530
rect 402980 370466 403032 370472
rect 403268 370394 403296 371311
rect 403256 370388 403308 370394
rect 403256 370330 403308 370336
rect 408512 368014 408540 371311
rect 412836 370802 412864 371855
rect 414018 371376 414074 371385
rect 414018 371311 414074 371320
rect 415398 371376 415454 371385
rect 415398 371311 415454 371320
rect 412824 370796 412876 370802
rect 412824 370738 412876 370744
rect 414032 370666 414060 371311
rect 415412 370870 415440 371311
rect 415400 370864 415452 370870
rect 415400 370806 415452 370812
rect 414020 370660 414072 370666
rect 414020 370602 414072 370608
rect 415688 369442 415716 374167
rect 445944 374138 445996 374144
rect 448256 374134 448284 374439
rect 448244 374128 448296 374134
rect 448244 374070 448296 374076
rect 421012 373924 421064 373930
rect 421012 373866 421064 373872
rect 421024 373833 421052 373866
rect 423036 373856 423088 373862
rect 421010 373824 421066 373833
rect 421010 373759 421066 373768
rect 423034 373824 423036 373833
rect 423088 373824 423090 373833
rect 423034 373759 423090 373768
rect 425426 373824 425482 373833
rect 425426 373759 425482 373768
rect 439410 373824 439466 373833
rect 439410 373759 439412 373768
rect 425440 373726 425468 373759
rect 439464 373759 439466 373768
rect 460938 373824 460994 373833
rect 460938 373759 460994 373768
rect 439412 373730 439464 373736
rect 425428 373720 425480 373726
rect 425428 373662 425480 373668
rect 438214 373144 438270 373153
rect 438214 373079 438270 373088
rect 426440 372700 426492 372706
rect 426440 372642 426492 372648
rect 425060 372632 425112 372638
rect 425058 372600 425060 372609
rect 426452 372609 426480 372642
rect 425112 372600 425114 372609
rect 425058 372535 425114 372544
rect 426438 372600 426494 372609
rect 426438 372535 426494 372544
rect 427818 372600 427874 372609
rect 438228 372570 438256 373079
rect 439424 372638 439452 373730
rect 450266 373688 450322 373697
rect 450266 373623 450268 373632
rect 450320 373623 450322 373632
rect 450268 373594 450320 373600
rect 460952 373590 460980 373759
rect 460940 373584 460992 373590
rect 452842 373552 452898 373561
rect 452842 373487 452844 373496
rect 452896 373487 452898 373496
rect 458178 373552 458234 373561
rect 460940 373526 460992 373532
rect 462778 373552 462834 373561
rect 458178 373487 458234 373496
rect 462778 373487 462834 373496
rect 452844 373458 452896 373464
rect 455418 373416 455474 373425
rect 455418 373351 455420 373360
rect 455472 373351 455474 373360
rect 455420 373322 455472 373328
rect 458192 373318 458220 373487
rect 462792 373454 462820 373487
rect 462780 373448 462832 373454
rect 462780 373390 462832 373396
rect 458180 373312 458232 373318
rect 458180 373254 458232 373260
rect 516692 372700 516744 372706
rect 516692 372642 516744 372648
rect 439412 372632 439464 372638
rect 439412 372574 439464 372580
rect 511908 372632 511960 372638
rect 511908 372574 511960 372580
rect 427818 372535 427874 372544
rect 438216 372564 438268 372570
rect 427832 372502 427860 372535
rect 438216 372506 438268 372512
rect 427820 372496 427872 372502
rect 427820 372438 427872 372444
rect 430578 371784 430634 371793
rect 430578 371719 430634 371728
rect 418250 371512 418306 371521
rect 418250 371447 418306 371456
rect 422298 371512 422354 371521
rect 422298 371447 422354 371456
rect 426438 371512 426494 371521
rect 426438 371447 426494 371456
rect 416778 371376 416834 371385
rect 416778 371311 416834 371320
rect 418158 371376 418214 371385
rect 418158 371311 418214 371320
rect 416792 370734 416820 371311
rect 416780 370728 416832 370734
rect 416780 370670 416832 370676
rect 418172 369510 418200 371311
rect 418160 369504 418212 369510
rect 418160 369446 418212 369452
rect 415676 369436 415728 369442
rect 415676 369378 415728 369384
rect 418264 369306 418292 371447
rect 422312 371414 422340 371447
rect 422300 371408 422352 371414
rect 419538 371376 419594 371385
rect 419538 371311 419594 371320
rect 420918 371376 420974 371385
rect 422300 371350 422352 371356
rect 423678 371376 423734 371385
rect 420918 371311 420974 371320
rect 423678 371311 423734 371320
rect 419552 369374 419580 371311
rect 419540 369368 419592 369374
rect 419540 369310 419592 369316
rect 418252 369300 418304 369306
rect 418252 369242 418304 369248
rect 420932 369073 420960 371311
rect 423692 369238 423720 371311
rect 423680 369232 423732 369238
rect 423680 369174 423732 369180
rect 420918 369064 420974 369073
rect 420918 368999 420974 369008
rect 408500 368008 408552 368014
rect 408500 367950 408552 367956
rect 426452 367946 426480 371447
rect 427818 371376 427874 371385
rect 427818 371311 427874 371320
rect 429198 371376 429254 371385
rect 429198 371311 429254 371320
rect 427832 369578 427860 371311
rect 427820 369572 427872 369578
rect 427820 369514 427872 369520
rect 426440 367940 426492 367946
rect 426440 367882 426492 367888
rect 429212 367878 429240 371311
rect 430592 369646 430620 371719
rect 438228 371414 438256 372506
rect 470598 372328 470654 372337
rect 470598 372263 470654 372272
rect 465078 371648 465134 371657
rect 465078 371583 465134 371592
rect 438216 371408 438268 371414
rect 430670 371376 430726 371385
rect 430670 371311 430726 371320
rect 431958 371376 432014 371385
rect 431958 371311 432014 371320
rect 436098 371376 436154 371385
rect 436098 371311 436154 371320
rect 437478 371376 437534 371385
rect 438216 371350 438268 371356
rect 437478 371311 437534 371320
rect 430580 369640 430632 369646
rect 430580 369582 430632 369588
rect 429200 367872 429252 367878
rect 429200 367814 429252 367820
rect 430684 367810 430712 371311
rect 431972 369170 432000 371311
rect 431960 369164 432012 369170
rect 431960 369106 432012 369112
rect 436112 368490 436140 371311
rect 437492 370938 437520 371311
rect 465092 371074 465120 371583
rect 467838 371376 467894 371385
rect 467838 371311 467894 371320
rect 465080 371068 465132 371074
rect 465080 371010 465132 371016
rect 467852 371006 467880 371311
rect 470612 371142 470640 372263
rect 503166 372192 503222 372201
rect 503166 372127 503222 372136
rect 483018 371920 483074 371929
rect 483018 371855 483074 371864
rect 473358 371376 473414 371385
rect 473358 371311 473414 371320
rect 480258 371376 480314 371385
rect 480258 371311 480314 371320
rect 473372 371210 473400 371311
rect 473360 371204 473412 371210
rect 473360 371146 473412 371152
rect 470600 371136 470652 371142
rect 470600 371078 470652 371084
rect 467840 371000 467892 371006
rect 467840 370942 467892 370948
rect 437480 370932 437532 370938
rect 437480 370874 437532 370880
rect 480272 369714 480300 371311
rect 483032 369782 483060 371855
rect 485778 371376 485834 371385
rect 485778 371311 485834 371320
rect 502338 371376 502394 371385
rect 503180 371346 503208 372127
rect 502338 371311 502394 371320
rect 503168 371340 503220 371346
rect 485792 369850 485820 371311
rect 502352 371278 502380 371311
rect 503168 371282 503220 371288
rect 502340 371272 502392 371278
rect 502260 371220 502340 371226
rect 502260 371214 502392 371220
rect 502260 371198 502380 371214
rect 485780 369844 485832 369850
rect 485780 369786 485832 369792
rect 483020 369776 483072 369782
rect 483020 369718 483072 369724
rect 480260 369708 480312 369714
rect 480260 369650 480312 369656
rect 436100 368484 436152 368490
rect 436100 368426 436152 368432
rect 430672 367804 430724 367810
rect 430672 367746 430724 367752
rect 500592 351348 500644 351354
rect 500592 351290 500644 351296
rect 499028 351280 499080 351286
rect 499028 351222 499080 351228
rect 499040 350577 499068 351222
rect 500604 350577 500632 351290
rect 499026 350568 499082 350577
rect 499026 350503 499082 350512
rect 500590 350568 500646 350577
rect 500590 350503 500646 350512
rect 502260 349858 502288 371198
rect 511920 350606 511948 372574
rect 516600 371408 516652 371414
rect 516600 371350 516652 371356
rect 510896 350600 510948 350606
rect 510894 350568 510896 350577
rect 511908 350600 511960 350606
rect 510948 350568 510950 350577
rect 511908 350542 511960 350548
rect 510894 350503 510950 350512
rect 502248 349852 502300 349858
rect 502248 349794 502300 349800
rect 380990 349752 381046 349761
rect 380990 349687 381046 349696
rect 380900 349580 380952 349586
rect 380900 349522 380952 349528
rect 425980 264920 426032 264926
rect 425980 264862 426032 264868
rect 473450 264888 473506 264897
rect 421104 264852 421156 264858
rect 421104 264794 421156 264800
rect 418436 264716 418488 264722
rect 418436 264658 418488 264664
rect 418448 264625 418476 264658
rect 421116 264625 421144 264794
rect 425992 264625 426020 264862
rect 473450 264823 473506 264832
rect 480902 264888 480958 264897
rect 480902 264823 480958 264832
rect 429752 264784 429804 264790
rect 429752 264726 429804 264732
rect 468482 264752 468538 264761
rect 429764 264625 429792 264726
rect 468482 264687 468538 264696
rect 470966 264752 471022 264761
rect 470966 264687 471022 264696
rect 468496 264654 468524 264687
rect 468484 264648 468536 264654
rect 418434 264616 418490 264625
rect 418434 264551 418490 264560
rect 421102 264616 421158 264625
rect 421102 264551 421158 264560
rect 423494 264616 423550 264625
rect 423494 264551 423550 264560
rect 425978 264616 426034 264625
rect 425978 264551 426034 264560
rect 429750 264616 429806 264625
rect 468484 264590 468536 264596
rect 429750 264551 429806 264560
rect 423508 264178 423536 264551
rect 470980 264450 471008 264687
rect 473464 264518 473492 264823
rect 475842 264616 475898 264625
rect 480916 264586 480944 264823
rect 483386 264752 483442 264761
rect 483386 264687 483442 264696
rect 485962 264752 486018 264761
rect 485962 264687 486018 264696
rect 475842 264551 475898 264560
rect 480904 264580 480956 264586
rect 473452 264512 473504 264518
rect 473452 264454 473504 264460
rect 470968 264444 471020 264450
rect 470968 264386 471020 264392
rect 475856 264246 475884 264551
rect 480904 264522 480956 264528
rect 483400 264382 483428 264687
rect 483388 264376 483440 264382
rect 483388 264318 483440 264324
rect 485976 264314 486004 264687
rect 485964 264308 486016 264314
rect 485964 264250 486016 264256
rect 475844 264240 475896 264246
rect 475844 264182 475896 264188
rect 423496 264172 423548 264178
rect 423496 264114 423548 264120
rect 433340 263696 433392 263702
rect 415858 263664 415914 263673
rect 433340 263638 433392 263644
rect 415858 263599 415914 263608
rect 432236 263628 432288 263634
rect 397458 263528 397514 263537
rect 397458 263463 397514 263472
rect 401598 263528 401654 263537
rect 401598 263463 401654 263472
rect 404358 263528 404414 263537
rect 404358 263463 404414 263472
rect 408314 263528 408370 263537
rect 408314 263463 408370 263472
rect 410706 263528 410762 263537
rect 410706 263463 410762 263472
rect 413650 263528 413706 263537
rect 413650 263463 413706 263472
rect 415766 263528 415822 263537
rect 415766 263463 415822 263472
rect 396078 262848 396134 262857
rect 396078 262783 396134 262792
rect 379980 262268 380032 262274
rect 379980 262210 380032 262216
rect 379888 241460 379940 241466
rect 379888 241402 379940 241408
rect 379796 241256 379848 241262
rect 379796 241198 379848 241204
rect 379704 241120 379756 241126
rect 379704 241062 379756 241068
rect 379888 240780 379940 240786
rect 379888 240722 379940 240728
rect 379900 240281 379928 240722
rect 379886 240272 379942 240281
rect 379886 240207 379942 240216
rect 379704 239896 379756 239902
rect 379704 239838 379756 239844
rect 379716 239601 379744 239838
rect 379702 239592 379758 239601
rect 379702 239527 379758 239536
rect 379796 151360 379848 151366
rect 379796 151302 379848 151308
rect 379704 151224 379756 151230
rect 379704 151166 379756 151172
rect 379716 150550 379744 151166
rect 379704 150544 379756 150550
rect 379704 150486 379756 150492
rect 379610 131064 379666 131073
rect 379610 130999 379666 131008
rect 379624 42090 379652 130999
rect 379716 44266 379744 150486
rect 379704 44260 379756 44266
rect 379704 44202 379756 44208
rect 379808 43858 379836 151302
rect 379900 130801 379928 240207
rect 379992 131102 380020 262210
rect 393412 261588 393464 261594
rect 393412 261530 393464 261536
rect 380348 261520 380400 261526
rect 380348 261462 380400 261468
rect 380360 260953 380388 261462
rect 389180 261044 389232 261050
rect 389180 260986 389232 260992
rect 388444 260976 388496 260982
rect 380346 260944 380402 260953
rect 388444 260918 388496 260924
rect 380346 260879 380402 260888
rect 388456 260778 388484 260918
rect 388444 260772 388496 260778
rect 388444 260714 388496 260720
rect 389192 260710 389220 260986
rect 390560 260908 390612 260914
rect 390560 260850 390612 260856
rect 389180 260704 389232 260710
rect 389180 260646 389232 260652
rect 390572 260642 390600 260850
rect 390560 260636 390612 260642
rect 390560 260578 390612 260584
rect 393424 260574 393452 261530
rect 393412 260568 393464 260574
rect 393412 260510 393464 260516
rect 393962 260128 394018 260137
rect 393962 260063 394018 260072
rect 393976 240825 394004 260063
rect 393962 240816 394018 240825
rect 393962 240751 394018 240760
rect 393976 239465 394004 240751
rect 396092 240514 396120 262783
rect 396170 262304 396226 262313
rect 396170 262239 396226 262248
rect 396184 262002 396212 262239
rect 396172 261996 396224 262002
rect 396172 261938 396224 261944
rect 396184 240650 396212 261938
rect 397472 240718 397500 263463
rect 398838 262304 398894 262313
rect 398838 262239 398894 262248
rect 400218 262304 400274 262313
rect 400218 262239 400274 262248
rect 398852 243710 398880 262239
rect 398840 243704 398892 243710
rect 398840 243646 398892 243652
rect 400232 243574 400260 262239
rect 401612 243642 401640 263463
rect 403070 262440 403126 262449
rect 403070 262375 403126 262384
rect 402978 262304 403034 262313
rect 402978 262239 403034 262248
rect 401600 243636 401652 243642
rect 401600 243578 401652 243584
rect 400220 243568 400272 243574
rect 400220 243510 400272 243516
rect 402992 241058 403020 262239
rect 402980 241052 403032 241058
rect 402980 240994 403032 241000
rect 403084 240990 403112 262375
rect 404372 241194 404400 263463
rect 408328 262750 408356 263463
rect 410720 262954 410748 263463
rect 410708 262948 410760 262954
rect 410708 262890 410760 262896
rect 413664 262886 413692 263463
rect 413652 262880 413704 262886
rect 412730 262848 412786 262857
rect 413652 262822 413704 262828
rect 415780 262818 415808 263463
rect 412730 262783 412786 262792
rect 415768 262812 415820 262818
rect 408316 262744 408368 262750
rect 408316 262686 408368 262692
rect 411258 262440 411314 262449
rect 411258 262375 411314 262384
rect 405738 262304 405794 262313
rect 405738 262239 405794 262248
rect 407210 262304 407266 262313
rect 407210 262239 407266 262248
rect 408498 262304 408554 262313
rect 408498 262239 408554 262248
rect 409878 262304 409934 262313
rect 409878 262239 409934 262248
rect 404360 241188 404412 241194
rect 404360 241130 404412 241136
rect 403072 240984 403124 240990
rect 403072 240926 403124 240932
rect 405752 240922 405780 262239
rect 407224 241330 407252 262239
rect 408512 241398 408540 262239
rect 408500 241392 408552 241398
rect 408500 241334 408552 241340
rect 407212 241324 407264 241330
rect 407212 241266 407264 241272
rect 409892 241126 409920 262239
rect 411272 241262 411300 262375
rect 411350 262304 411406 262313
rect 411350 262239 411406 262248
rect 411260 241256 411312 241262
rect 411260 241198 411312 241204
rect 409880 241120 409932 241126
rect 409880 241062 409932 241068
rect 405740 240916 405792 240922
rect 405740 240858 405792 240864
rect 411364 240854 411392 262239
rect 412744 241466 412772 262783
rect 415768 262754 415820 262760
rect 414018 262304 414074 262313
rect 415872 262274 415900 263599
rect 432236 263570 432288 263576
rect 432248 263537 432276 263570
rect 433352 263537 433380 263638
rect 453396 263560 453448 263566
rect 419354 263528 419410 263537
rect 419354 263463 419410 263472
rect 425242 263528 425298 263537
rect 425242 263463 425298 263472
rect 426438 263528 426494 263537
rect 426438 263463 426494 263472
rect 427450 263528 427506 263537
rect 427450 263463 427506 263472
rect 428186 263528 428242 263537
rect 428186 263463 428242 263472
rect 430946 263528 431002 263537
rect 430946 263463 431002 263472
rect 432234 263528 432290 263537
rect 432234 263463 432290 263472
rect 433338 263528 433394 263537
rect 433338 263463 433394 263472
rect 434626 263528 434682 263537
rect 435914 263528 435970 263537
rect 434682 263486 434760 263514
rect 434626 263463 434682 263472
rect 418158 262848 418214 262857
rect 418158 262783 418214 262792
rect 416778 262304 416834 262313
rect 414018 262239 414074 262248
rect 415860 262268 415912 262274
rect 412732 241460 412784 241466
rect 412732 241402 412784 241408
rect 411352 240848 411404 240854
rect 411352 240790 411404 240796
rect 414032 240786 414060 262239
rect 416778 262239 416834 262248
rect 415860 262210 415912 262216
rect 416792 240825 416820 262239
rect 418172 260574 418200 262783
rect 419368 260642 419396 263463
rect 419814 262984 419870 262993
rect 419814 262919 419870 262928
rect 421746 262984 421802 262993
rect 421746 262919 421802 262928
rect 419828 260710 419856 262919
rect 421760 260778 421788 262919
rect 423954 262576 424010 262585
rect 423954 262511 424010 262520
rect 423586 262304 423642 262313
rect 423642 262262 423720 262290
rect 423586 262239 423642 262248
rect 421748 260772 421800 260778
rect 421748 260714 421800 260720
rect 419816 260704 419868 260710
rect 419816 260646 419868 260652
rect 419356 260636 419408 260642
rect 419356 260578 419408 260584
rect 418160 260568 418212 260574
rect 418160 260510 418212 260516
rect 416778 240816 416834 240825
rect 414020 240780 414072 240786
rect 416778 240751 416834 240760
rect 414020 240722 414072 240728
rect 397460 240712 397512 240718
rect 397460 240654 397512 240660
rect 396172 240644 396224 240650
rect 396172 240586 396224 240592
rect 396080 240508 396132 240514
rect 396080 240450 396132 240456
rect 423692 239970 423720 262262
rect 423968 260234 423996 262511
rect 425256 261526 425284 263463
rect 425704 262268 425756 262274
rect 425704 262210 425756 262216
rect 425244 261520 425296 261526
rect 425244 261462 425296 261468
rect 423956 260228 424008 260234
rect 423956 260170 424008 260176
rect 423680 239964 423732 239970
rect 423680 239906 423732 239912
rect 425716 239902 425744 262210
rect 426452 262070 426480 263463
rect 426440 262064 426492 262070
rect 426440 262006 426492 262012
rect 427464 260166 427492 263463
rect 428200 262138 428228 263463
rect 428278 262304 428334 262313
rect 428278 262239 428280 262248
rect 428332 262239 428334 262248
rect 430670 262304 430726 262313
rect 430670 262239 430726 262248
rect 428280 262210 428332 262216
rect 428188 262132 428240 262138
rect 428188 262074 428240 262080
rect 427452 260160 427504 260166
rect 427452 260102 427504 260108
rect 425704 239896 425756 239902
rect 425704 239838 425756 239844
rect 393962 239456 394018 239465
rect 430684 239426 430712 262239
rect 430960 262206 430988 263463
rect 433524 263016 433576 263022
rect 433522 262984 433524 262993
rect 433576 262984 433578 262993
rect 433522 262919 433578 262928
rect 430948 262200 431000 262206
rect 430948 262142 431000 262148
rect 434732 240038 434760 263486
rect 435914 263463 435970 263472
rect 438766 263528 438822 263537
rect 438766 263463 438822 263472
rect 440882 263528 440938 263537
rect 440882 263463 440938 263472
rect 443458 263528 443514 263537
rect 443458 263463 443514 263472
rect 448242 263528 448298 263537
rect 448242 263463 448298 263472
rect 451002 263528 451058 263537
rect 451002 263463 451058 263472
rect 453394 263528 453396 263537
rect 453448 263528 453450 263537
rect 453394 263463 453450 263472
rect 455786 263528 455842 263537
rect 455786 263463 455788 263472
rect 435928 263158 435956 263463
rect 438400 263288 438452 263294
rect 438400 263230 438452 263236
rect 435916 263152 435968 263158
rect 435916 263094 435968 263100
rect 438412 262993 438440 263230
rect 435178 262984 435234 262993
rect 435178 262919 435234 262928
rect 438398 262984 438454 262993
rect 438398 262919 438454 262928
rect 435192 260846 435220 262919
rect 436098 262304 436154 262313
rect 436098 262239 436154 262248
rect 435180 260840 435232 260846
rect 435180 260782 435232 260788
rect 436112 240106 436140 262239
rect 438780 241466 438808 263463
rect 440896 263090 440924 263463
rect 443472 263362 443500 263463
rect 443460 263356 443512 263362
rect 443460 263298 443512 263304
rect 448256 263226 448284 263463
rect 451016 263430 451044 263463
rect 455840 263463 455842 263472
rect 503534 263528 503590 263537
rect 503534 263463 503590 263472
rect 455788 263434 455840 263440
rect 451004 263424 451056 263430
rect 451004 263366 451056 263372
rect 448244 263220 448296 263226
rect 448244 263162 448296 263168
rect 503548 263090 503576 263463
rect 440884 263084 440936 263090
rect 440884 263026 440936 263032
rect 503536 263084 503588 263090
rect 503536 263026 503588 263032
rect 503628 262948 503680 262954
rect 503628 262890 503680 262896
rect 503640 262313 503668 262890
rect 511908 262472 511960 262478
rect 511908 262414 511960 262420
rect 440146 262304 440202 262313
rect 440146 262239 440202 262248
rect 503626 262304 503682 262313
rect 503626 262239 503682 262248
rect 440160 244254 440188 262239
rect 440148 244248 440200 244254
rect 440148 244190 440200 244196
rect 438768 241460 438820 241466
rect 438768 241402 438820 241408
rect 503640 240990 503668 262239
rect 511920 241505 511948 262414
rect 511906 241496 511962 241505
rect 516612 241466 516640 371350
rect 516704 244254 516732 372642
rect 517532 372638 517560 461858
rect 517796 461032 517848 461038
rect 517796 460974 517848 460980
rect 517612 460964 517664 460970
rect 517612 460906 517664 460912
rect 517520 372632 517572 372638
rect 517520 372574 517572 372580
rect 517624 364334 517652 460906
rect 517624 364306 517744 364334
rect 517716 351354 517744 364306
rect 517704 351348 517756 351354
rect 517704 351290 517756 351296
rect 517520 350600 517572 350606
rect 517520 350542 517572 350548
rect 517532 262478 517560 350542
rect 517612 349852 517664 349858
rect 517612 349794 517664 349800
rect 517624 263090 517652 349794
rect 517612 263084 517664 263090
rect 517612 263026 517664 263032
rect 517520 262472 517572 262478
rect 517520 262414 517572 262420
rect 516692 244248 516744 244254
rect 516692 244190 516744 244196
rect 511906 241431 511962 241440
rect 516600 241460 516652 241466
rect 503628 240984 503680 240990
rect 503628 240926 503680 240932
rect 500776 240916 500828 240922
rect 500776 240858 500828 240864
rect 499028 240848 499080 240854
rect 499028 240790 499080 240796
rect 499040 240281 499068 240790
rect 500788 240281 500816 240858
rect 511920 240650 511948 241431
rect 516600 241402 516652 241408
rect 511908 240644 511960 240650
rect 511908 240586 511960 240592
rect 499026 240272 499082 240281
rect 499026 240207 499082 240216
rect 500774 240272 500830 240281
rect 500774 240207 500830 240216
rect 436100 240100 436152 240106
rect 436100 240042 436152 240048
rect 434720 240032 434772 240038
rect 434720 239974 434772 239980
rect 393962 239391 394018 239400
rect 430672 239420 430724 239426
rect 430672 239362 430724 239368
rect 418436 154556 418488 154562
rect 418436 154498 418488 154504
rect 418448 154465 418476 154498
rect 421012 154488 421064 154494
rect 418434 154456 418490 154465
rect 418434 154391 418490 154400
rect 421010 154456 421012 154465
rect 421064 154456 421066 154465
rect 421010 154391 421066 154400
rect 425978 154456 426034 154465
rect 443458 154456 443514 154465
rect 425978 154391 425980 154400
rect 426032 154391 426034 154400
rect 438860 154420 438912 154426
rect 425980 154362 426032 154368
rect 516612 154426 516640 241402
rect 443458 154391 443514 154400
rect 516600 154420 516652 154426
rect 438860 154362 438912 154368
rect 423402 153912 423458 153921
rect 423402 153847 423458 153856
rect 423416 153814 423444 153847
rect 423404 153808 423456 153814
rect 423404 153750 423456 153756
rect 431960 153264 432012 153270
rect 431960 153206 432012 153212
rect 431972 153105 432000 153206
rect 438872 153105 438900 154362
rect 443472 154358 443500 154391
rect 516600 154362 516652 154368
rect 443460 154352 443512 154358
rect 443460 154294 443512 154300
rect 475842 154320 475898 154329
rect 475842 154255 475844 154264
rect 475896 154255 475898 154264
rect 478418 154320 478474 154329
rect 478418 154255 478474 154264
rect 475844 154226 475896 154232
rect 478432 154222 478460 154255
rect 478420 154216 478472 154222
rect 473450 154184 473506 154193
rect 478420 154158 478472 154164
rect 480810 154184 480866 154193
rect 473450 154119 473452 154128
rect 473504 154119 473506 154128
rect 480810 154119 480866 154128
rect 473452 154090 473504 154096
rect 480824 154086 480852 154119
rect 480812 154080 480864 154086
rect 470874 154048 470930 154057
rect 480812 154022 480864 154028
rect 483202 154048 483258 154057
rect 470874 153983 470876 153992
rect 470928 153983 470930 153992
rect 483202 153983 483258 153992
rect 510528 154012 510580 154018
rect 470876 153954 470928 153960
rect 483216 153950 483244 153983
rect 510528 153954 510580 153960
rect 483204 153944 483256 153950
rect 483204 153886 483256 153892
rect 485962 153912 486018 153921
rect 485962 153847 485964 153856
rect 486016 153847 486018 153856
rect 485964 153818 486016 153824
rect 455420 153196 455472 153202
rect 455420 153138 455472 153144
rect 447140 153128 447192 153134
rect 396078 153096 396134 153105
rect 396078 153031 396134 153040
rect 397458 153096 397514 153105
rect 397458 153031 397514 153040
rect 398838 153096 398894 153105
rect 398838 153031 398894 153040
rect 400218 153096 400274 153105
rect 400218 153031 400274 153040
rect 401598 153096 401654 153105
rect 401598 153031 401654 153040
rect 403070 153096 403126 153105
rect 403070 153031 403126 153040
rect 404358 153096 404414 153105
rect 404358 153031 404414 153040
rect 405738 153096 405794 153105
rect 405738 153031 405794 153040
rect 407210 153096 407266 153105
rect 407210 153031 407266 153040
rect 408498 153096 408554 153105
rect 408498 153031 408554 153040
rect 409970 153096 410026 153105
rect 409970 153031 410026 153040
rect 411350 153096 411406 153105
rect 411350 153031 411406 153040
rect 412730 153096 412786 153105
rect 412730 153031 412786 153040
rect 414018 153096 414074 153105
rect 414018 153031 414074 153040
rect 415490 153096 415546 153105
rect 415490 153031 415546 153040
rect 415674 153096 415730 153105
rect 415674 153031 415730 153040
rect 416778 153096 416834 153105
rect 416778 153031 416834 153040
rect 418250 153096 418306 153105
rect 418250 153031 418306 153040
rect 419538 153096 419594 153105
rect 419538 153031 419594 153040
rect 420918 153096 420974 153105
rect 420918 153031 420974 153040
rect 422298 153096 422354 153105
rect 422298 153031 422354 153040
rect 423678 153096 423734 153105
rect 423678 153031 423734 153040
rect 425058 153096 425114 153105
rect 425058 153031 425114 153040
rect 426530 153096 426586 153105
rect 426530 153031 426586 153040
rect 427818 153096 427874 153105
rect 427818 153031 427874 153040
rect 429198 153096 429254 153105
rect 429198 153031 429254 153040
rect 430578 153096 430634 153105
rect 430578 153031 430634 153040
rect 431958 153096 432014 153105
rect 431958 153031 432014 153040
rect 433338 153096 433394 153105
rect 433338 153031 433394 153040
rect 433982 153096 434038 153105
rect 433982 153031 434038 153040
rect 434810 153096 434866 153105
rect 434810 153031 434866 153040
rect 436190 153096 436246 153105
rect 436190 153031 436246 153040
rect 438858 153096 438914 153105
rect 438858 153031 438914 153040
rect 440146 153096 440202 153105
rect 440146 153031 440202 153040
rect 440330 153096 440386 153105
rect 440330 153031 440386 153040
rect 445758 153096 445814 153105
rect 445758 153031 445814 153040
rect 447138 153096 447140 153105
rect 455432 153105 455460 153138
rect 447192 153096 447194 153105
rect 447138 153031 447194 153040
rect 449898 153096 449954 153105
rect 449898 153031 449954 153040
rect 452658 153096 452714 153105
rect 452658 153031 452714 153040
rect 455418 153096 455474 153105
rect 455418 153031 455474 153040
rect 458178 153096 458234 153105
rect 458178 153031 458180 153040
rect 380808 151632 380860 151638
rect 380808 151574 380860 151580
rect 380072 151564 380124 151570
rect 380072 151506 380124 151512
rect 380084 151298 380112 151506
rect 380164 151360 380216 151366
rect 380820 151337 380848 151574
rect 380164 151302 380216 151308
rect 380806 151328 380862 151337
rect 380072 151292 380124 151298
rect 380072 151234 380124 151240
rect 380176 150822 380204 151302
rect 380806 151263 380862 151272
rect 396092 150958 396120 153031
rect 396170 152552 396226 152561
rect 396170 152487 396226 152496
rect 396080 150952 396132 150958
rect 396080 150894 396132 150900
rect 380164 150816 380216 150822
rect 380164 150758 380216 150764
rect 379980 131096 380032 131102
rect 379980 131038 380032 131044
rect 379886 130792 379942 130801
rect 379886 130727 379942 130736
rect 379900 44538 379928 130727
rect 379992 129810 380020 131038
rect 380072 130824 380124 130830
rect 380072 130766 380124 130772
rect 380084 130558 380112 130766
rect 380256 130620 380308 130626
rect 380256 130562 380308 130568
rect 380072 130552 380124 130558
rect 380072 130494 380124 130500
rect 380164 130552 380216 130558
rect 380164 130494 380216 130500
rect 380176 130150 380204 130494
rect 380164 130144 380216 130150
rect 380164 130086 380216 130092
rect 380268 130082 380296 130562
rect 396092 130218 396120 150894
rect 396184 150890 396212 152487
rect 396172 150884 396224 150890
rect 396172 150826 396224 150832
rect 396184 130286 396212 150826
rect 397472 130354 397500 153031
rect 398852 133210 398880 153031
rect 400232 133618 400260 153031
rect 401612 133686 401640 153031
rect 402978 152552 403034 152561
rect 402978 152487 403034 152496
rect 401600 133680 401652 133686
rect 401600 133622 401652 133628
rect 400220 133612 400272 133618
rect 400220 133554 400272 133560
rect 398840 133204 398892 133210
rect 398840 133146 398892 133152
rect 402992 130762 403020 152487
rect 402980 130756 403032 130762
rect 402980 130698 403032 130704
rect 403084 130626 403112 153031
rect 403072 130620 403124 130626
rect 403072 130562 403124 130568
rect 404372 130490 404400 153031
rect 405752 130694 405780 153031
rect 407118 152416 407174 152425
rect 407118 152351 407174 152360
rect 407132 152318 407160 152351
rect 407120 152312 407172 152318
rect 407120 152254 407172 152260
rect 405740 130688 405792 130694
rect 405740 130630 405792 130636
rect 407224 130558 407252 153031
rect 408512 130830 408540 153031
rect 409878 152552 409934 152561
rect 409878 152487 409934 152496
rect 409892 152386 409920 152487
rect 409880 152380 409932 152386
rect 409880 152322 409932 152328
rect 409984 130898 410012 153031
rect 411258 152552 411314 152561
rect 411258 152487 411314 152496
rect 411272 131034 411300 152487
rect 411260 131028 411312 131034
rect 411260 130970 411312 130976
rect 411364 130966 411392 153031
rect 412744 133754 412772 153031
rect 413098 152552 413154 152561
rect 413098 152487 413154 152496
rect 413112 152454 413140 152487
rect 413100 152448 413152 152454
rect 413100 152390 413152 152396
rect 412732 133748 412784 133754
rect 412732 133690 412784 133696
rect 411352 130960 411404 130966
rect 411352 130902 411404 130908
rect 409972 130892 410024 130898
rect 409972 130834 410024 130840
rect 408500 130824 408552 130830
rect 414032 130801 414060 153031
rect 415504 142154 415532 153031
rect 415688 152522 415716 153031
rect 415676 152516 415728 152522
rect 415676 152458 415728 152464
rect 415412 142126 415532 142154
rect 415412 131102 415440 142126
rect 415400 131096 415452 131102
rect 415400 131038 415452 131044
rect 416792 130937 416820 153031
rect 418158 152552 418214 152561
rect 418158 152487 418214 152496
rect 418172 151298 418200 152487
rect 418264 151366 418292 153031
rect 418252 151360 418304 151366
rect 418252 151302 418304 151308
rect 418160 151292 418212 151298
rect 418160 151234 418212 151240
rect 419552 151026 419580 153031
rect 420932 151434 420960 153031
rect 422312 151570 422340 153031
rect 422300 151564 422352 151570
rect 422300 151506 422352 151512
rect 420920 151428 420972 151434
rect 420920 151370 420972 151376
rect 423692 151230 423720 153031
rect 425072 151502 425100 153031
rect 426438 152552 426494 152561
rect 426438 152487 426494 152496
rect 425060 151496 425112 151502
rect 425060 151438 425112 151444
rect 423680 151224 423732 151230
rect 423680 151166 423732 151172
rect 419540 151020 419592 151026
rect 419540 150962 419592 150968
rect 426452 131073 426480 152487
rect 426544 151706 426572 153031
rect 426532 151700 426584 151706
rect 426532 151642 426584 151648
rect 427832 151638 427860 153031
rect 427820 151632 427872 151638
rect 427820 151574 427872 151580
rect 426438 131064 426494 131073
rect 426438 130999 426494 131008
rect 416778 130928 416834 130937
rect 416778 130863 416834 130872
rect 408500 130766 408552 130772
rect 414018 130792 414074 130801
rect 414018 130727 414074 130736
rect 407212 130552 407264 130558
rect 407212 130494 407264 130500
rect 404360 130484 404412 130490
rect 404360 130426 404412 130432
rect 429212 130393 429240 153031
rect 430592 151162 430620 153031
rect 433352 152590 433380 153031
rect 433340 152584 433392 152590
rect 433340 152526 433392 152532
rect 430580 151156 430632 151162
rect 430580 151098 430632 151104
rect 433996 151094 434024 153031
rect 434824 152726 434852 153031
rect 434812 152720 434864 152726
rect 434812 152662 434864 152668
rect 434718 152552 434774 152561
rect 434718 152487 434774 152496
rect 436098 152552 436154 152561
rect 436098 152487 436154 152496
rect 433984 151088 434036 151094
rect 433984 151030 434036 151036
rect 434732 133822 434760 152487
rect 436112 133890 436140 152487
rect 436204 151774 436232 153031
rect 437480 152652 437532 152658
rect 437480 152594 437532 152600
rect 437492 152561 437520 152594
rect 437478 152552 437534 152561
rect 437478 152487 437534 152496
rect 436192 151768 436244 151774
rect 436192 151710 436244 151716
rect 436100 133884 436152 133890
rect 436100 133826 436152 133832
rect 434720 133816 434772 133822
rect 434720 133758 434772 133764
rect 438872 133113 438900 153031
rect 438858 133104 438914 133113
rect 438858 133039 438914 133048
rect 440160 130490 440188 153031
rect 440344 152862 440372 153031
rect 445772 152930 445800 153031
rect 445760 152924 445812 152930
rect 445760 152866 445812 152872
rect 440332 152856 440384 152862
rect 440332 152798 440384 152804
rect 449912 152794 449940 153031
rect 452672 152998 452700 153031
rect 458232 153031 458234 153040
rect 458180 153002 458232 153008
rect 452660 152992 452712 152998
rect 452660 152934 452712 152940
rect 449900 152788 449952 152794
rect 449900 152730 449952 152736
rect 503626 152688 503682 152697
rect 503626 152623 503628 152632
rect 503680 152623 503682 152632
rect 503628 152594 503680 152600
rect 503626 152552 503682 152561
rect 503626 152487 503628 152496
rect 503680 152487 503682 152496
rect 503628 152458 503680 152464
rect 500224 131028 500276 131034
rect 500224 130970 500276 130976
rect 498752 130960 498804 130966
rect 498752 130902 498804 130908
rect 440148 130484 440200 130490
rect 440148 130426 440200 130432
rect 466460 130484 466512 130490
rect 466460 130426 466512 130432
rect 429198 130384 429254 130393
rect 397460 130348 397512 130354
rect 429198 130319 429254 130328
rect 397460 130290 397512 130296
rect 396172 130280 396224 130286
rect 396172 130222 396224 130228
rect 396080 130212 396132 130218
rect 396080 130154 396132 130160
rect 380256 130076 380308 130082
rect 380256 130018 380308 130024
rect 379980 129804 380032 129810
rect 379980 129746 380032 129752
rect 466472 129742 466500 130426
rect 498764 129849 498792 130902
rect 500236 129849 500264 130970
rect 503640 130490 503668 152458
rect 510540 130506 510568 153954
rect 516704 132494 516732 244190
rect 517520 240644 517572 240650
rect 517520 240586 517572 240592
rect 517532 154018 517560 240586
rect 517520 154012 517572 154018
rect 517520 153954 517572 153960
rect 517624 152658 517652 263026
rect 517716 240922 517744 351290
rect 517808 351286 517836 460974
rect 518176 441590 518204 530538
rect 578884 529236 578936 529242
rect 578884 529178 578936 529184
rect 540244 502376 540296 502382
rect 540244 502318 540296 502324
rect 518898 454200 518954 454209
rect 518898 454135 518954 454144
rect 518164 441584 518216 441590
rect 518164 441526 518216 441532
rect 517888 371340 517940 371346
rect 517888 371282 517940 371288
rect 517796 351280 517848 351286
rect 517796 351222 517848 351228
rect 517704 240916 517756 240922
rect 517704 240858 517756 240864
rect 517612 152652 517664 152658
rect 517612 152594 517664 152600
rect 517624 142154 517652 152594
rect 516612 132466 516732 132494
rect 517532 142126 517652 142154
rect 503628 130484 503680 130490
rect 510540 130478 510660 130506
rect 503628 130426 503680 130432
rect 510632 130422 510660 130478
rect 510620 130416 510672 130422
rect 510618 130384 510620 130393
rect 510672 130384 510674 130393
rect 510618 130319 510674 130328
rect 498750 129840 498806 129849
rect 498750 129775 498806 129784
rect 500222 129840 500278 129849
rect 500222 129775 500278 129784
rect 516612 129742 516640 132466
rect 466460 129736 466512 129742
rect 466460 129678 466512 129684
rect 516600 129736 516652 129742
rect 516600 129678 516652 129684
rect 396078 44840 396134 44849
rect 396078 44775 396134 44784
rect 397090 44840 397146 44849
rect 397090 44775 397146 44784
rect 403070 44840 403126 44849
rect 403070 44775 403126 44784
rect 414570 44840 414626 44849
rect 414570 44775 414626 44784
rect 416962 44840 417018 44849
rect 416962 44775 417018 44784
rect 396092 44674 396120 44775
rect 397104 44742 397132 44775
rect 397092 44736 397144 44742
rect 397092 44678 397144 44684
rect 396080 44668 396132 44674
rect 396080 44610 396132 44616
rect 403084 44606 403112 44775
rect 410706 44704 410762 44713
rect 410706 44639 410762 44648
rect 403072 44600 403124 44606
rect 403072 44542 403124 44548
rect 404174 44568 404230 44577
rect 379888 44532 379940 44538
rect 404174 44503 404230 44512
rect 405462 44568 405518 44577
rect 405462 44503 405518 44512
rect 406474 44568 406530 44577
rect 406474 44503 406530 44512
rect 379888 44474 379940 44480
rect 379796 43852 379848 43858
rect 379796 43794 379848 43800
rect 404188 43314 404216 44503
rect 405476 44062 405504 44503
rect 406488 44130 406516 44503
rect 410720 44198 410748 44639
rect 414584 44538 414612 44775
rect 414572 44532 414624 44538
rect 414572 44474 414624 44480
rect 416976 44470 417004 44775
rect 419446 44704 419502 44713
rect 419446 44639 419502 44648
rect 423954 44704 424010 44713
rect 423954 44639 424010 44648
rect 418158 44568 418214 44577
rect 418158 44503 418214 44512
rect 416964 44464 417016 44470
rect 416964 44406 417016 44412
rect 418172 44334 418200 44503
rect 419460 44402 419488 44639
rect 420642 44568 420698 44577
rect 420642 44503 420698 44512
rect 421746 44568 421802 44577
rect 421746 44503 421802 44512
rect 422850 44568 422906 44577
rect 422850 44503 422906 44512
rect 419448 44396 419500 44402
rect 419448 44338 419500 44344
rect 418160 44328 418212 44334
rect 418160 44270 418212 44276
rect 410708 44192 410760 44198
rect 410708 44134 410760 44140
rect 406476 44124 406528 44130
rect 406476 44066 406528 44072
rect 405464 44056 405516 44062
rect 405464 43998 405516 44004
rect 420656 43994 420684 44503
rect 420644 43988 420696 43994
rect 420644 43930 420696 43936
rect 421760 43926 421788 44503
rect 421748 43920 421800 43926
rect 421748 43862 421800 43868
rect 422864 43790 422892 44503
rect 423968 44266 423996 44639
rect 425978 44568 426034 44577
rect 425978 44503 426034 44512
rect 439226 44568 439282 44577
rect 439226 44503 439282 44512
rect 455878 44568 455934 44577
rect 455878 44503 455934 44512
rect 458454 44568 458510 44577
rect 458454 44503 458510 44512
rect 425242 44432 425298 44441
rect 425242 44367 425298 44376
rect 423956 44260 424008 44266
rect 423956 44202 424008 44208
rect 425256 43858 425284 44367
rect 425244 43852 425296 43858
rect 425244 43794 425296 43800
rect 422852 43784 422904 43790
rect 422852 43726 422904 43732
rect 425992 43722 426020 44503
rect 425980 43716 426032 43722
rect 425980 43658 426032 43664
rect 421012 43580 421064 43586
rect 421012 43522 421064 43528
rect 421024 43489 421052 43522
rect 407578 43480 407634 43489
rect 407578 43415 407634 43424
rect 421010 43480 421066 43489
rect 421010 43415 421066 43424
rect 428186 43480 428242 43489
rect 439240 43450 439268 44503
rect 455892 43518 455920 44503
rect 458468 43654 458496 44503
rect 458456 43648 458508 43654
rect 458456 43590 458508 43596
rect 455880 43512 455932 43518
rect 455880 43454 455932 43460
rect 516612 43450 516640 129678
rect 428186 43415 428188 43424
rect 407592 43382 407620 43415
rect 428240 43415 428242 43424
rect 439228 43444 439280 43450
rect 428188 43386 428240 43392
rect 439228 43386 439280 43392
rect 516600 43444 516652 43450
rect 516600 43386 516652 43392
rect 407580 43376 407632 43382
rect 407580 43318 407632 43324
rect 404176 43308 404228 43314
rect 404176 43250 404228 43256
rect 398194 43208 398250 43217
rect 398194 43143 398250 43152
rect 401690 43208 401746 43217
rect 401690 43143 401746 43152
rect 379612 42084 379664 42090
rect 379612 42026 379664 42032
rect 379428 41268 379480 41274
rect 379428 41210 379480 41216
rect 398208 41002 398236 43143
rect 399390 42800 399446 42809
rect 399390 42735 399446 42744
rect 398196 40996 398248 41002
rect 398196 40938 398248 40944
rect 399404 40050 399432 42735
rect 400310 41848 400366 41857
rect 400310 41783 400366 41792
rect 399392 40044 399444 40050
rect 399392 39986 399444 39992
rect 379336 39636 379388 39642
rect 379336 39578 379388 39584
rect 376576 39568 376628 39574
rect 376576 39510 376628 39516
rect 400324 39506 400352 41783
rect 401704 41070 401732 43143
rect 408314 42800 408370 42809
rect 408314 42735 408370 42744
rect 408682 42800 408738 42809
rect 408682 42735 408738 42744
rect 409970 42800 410026 42809
rect 409970 42735 410026 42744
rect 411258 42800 411314 42809
rect 411258 42735 411314 42744
rect 411902 42800 411958 42809
rect 411902 42735 411958 42744
rect 413282 42800 413338 42809
rect 413282 42735 413338 42744
rect 413650 42800 413706 42809
rect 413650 42735 413706 42744
rect 415490 42800 415546 42809
rect 415490 42735 415546 42744
rect 426438 42800 426494 42809
rect 426438 42735 426494 42744
rect 427634 42800 427690 42809
rect 427634 42735 427690 42744
rect 428554 42800 428610 42809
rect 428554 42735 428610 42744
rect 429658 42800 429714 42809
rect 429658 42735 429714 42744
rect 430946 42800 431002 42809
rect 430946 42735 431002 42744
rect 432142 42800 432198 42809
rect 432142 42735 432198 42744
rect 433338 42800 433394 42809
rect 433338 42735 433394 42744
rect 434626 42800 434682 42809
rect 434626 42735 434682 42744
rect 435914 42800 435970 42809
rect 435914 42735 435970 42744
rect 436374 42800 436430 42809
rect 436374 42735 436430 42744
rect 438490 42800 438546 42809
rect 438490 42735 438546 42744
rect 440882 42800 440938 42809
rect 440882 42735 440938 42744
rect 443458 42800 443514 42809
rect 443458 42735 443514 42744
rect 445850 42800 445906 42809
rect 445850 42735 445906 42744
rect 448242 42800 448298 42809
rect 448242 42735 448298 42744
rect 453394 42800 453450 42809
rect 453394 42735 453450 42744
rect 485962 42800 486018 42809
rect 485962 42735 485964 42744
rect 408328 41410 408356 42735
rect 408316 41404 408368 41410
rect 408316 41346 408368 41352
rect 401692 41064 401744 41070
rect 401692 41006 401744 41012
rect 408696 39574 408724 42735
rect 409984 41138 410012 42735
rect 409972 41132 410024 41138
rect 409972 41074 410024 41080
rect 411272 39642 411300 42735
rect 411916 39710 411944 42735
rect 413296 41206 413324 42735
rect 413664 42158 413692 42735
rect 413652 42152 413704 42158
rect 413652 42094 413704 42100
rect 415504 42022 415532 42735
rect 415492 42016 415544 42022
rect 415492 41958 415544 41964
rect 426452 41274 426480 42735
rect 427648 42090 427676 42735
rect 427636 42084 427688 42090
rect 427636 42026 427688 42032
rect 426440 41268 426492 41274
rect 426440 41210 426492 41216
rect 413284 41200 413336 41206
rect 413284 41142 413336 41148
rect 428568 40905 428596 42735
rect 429672 41342 429700 42735
rect 430960 42226 430988 42735
rect 430948 42220 431000 42226
rect 430948 42162 431000 42168
rect 431130 41984 431186 41993
rect 431130 41919 431186 41928
rect 429660 41336 429712 41342
rect 429660 41278 429712 41284
rect 428554 40896 428610 40905
rect 428554 40831 428610 40840
rect 431144 39778 431172 41919
rect 432156 39846 432184 42735
rect 433352 41041 433380 42735
rect 433338 41032 433394 41041
rect 433338 40967 433394 40976
rect 434640 39914 434668 42735
rect 435928 42430 435956 42735
rect 435916 42424 435968 42430
rect 435916 42366 435968 42372
rect 435178 42120 435234 42129
rect 435178 42055 435234 42064
rect 434628 39908 434680 39914
rect 434628 39850 434680 39856
rect 432144 39840 432196 39846
rect 432144 39782 432196 39788
rect 431132 39772 431184 39778
rect 431132 39714 431184 39720
rect 411904 39704 411956 39710
rect 411904 39646 411956 39652
rect 411260 39636 411312 39642
rect 411260 39578 411312 39584
rect 408684 39568 408736 39574
rect 408684 39510 408736 39516
rect 400312 39500 400364 39506
rect 400312 39442 400364 39448
rect 435192 39438 435220 42055
rect 436388 39982 436416 42735
rect 438504 42294 438532 42735
rect 440896 42362 440924 42735
rect 443472 42498 443500 42735
rect 445864 42566 445892 42735
rect 448256 42634 448284 42735
rect 453408 42702 453436 42735
rect 486016 42735 486018 42744
rect 503258 42800 503314 42809
rect 503258 42735 503260 42744
rect 485964 42706 486016 42712
rect 503312 42735 503314 42744
rect 503534 42800 503590 42809
rect 503534 42735 503590 42744
rect 503260 42706 503312 42712
rect 503548 42702 503576 42735
rect 517532 42702 517560 142126
rect 517716 131034 517744 240858
rect 517808 240854 517836 351222
rect 517900 262954 517928 371282
rect 518912 354674 518940 454135
rect 519174 393816 519230 393825
rect 519174 393751 519230 393760
rect 518990 390824 519046 390833
rect 518990 390759 519046 390768
rect 519004 356794 519032 390759
rect 519082 389328 519138 389337
rect 519082 389263 519138 389272
rect 519096 360874 519124 389263
rect 519084 360868 519136 360874
rect 519084 360810 519136 360816
rect 519188 359582 519216 393751
rect 519358 392184 519414 392193
rect 519358 392119 519414 392128
rect 519266 388104 519322 388113
rect 519266 388039 519322 388048
rect 519176 359576 519228 359582
rect 519176 359518 519228 359524
rect 519280 358086 519308 388039
rect 519372 366382 519400 392119
rect 519360 366376 519412 366382
rect 519360 366318 519412 366324
rect 519372 364334 519400 366318
rect 519372 364306 519492 364334
rect 519360 359576 519412 359582
rect 519360 359518 519412 359524
rect 519268 358080 519320 358086
rect 519268 358022 519320 358028
rect 518992 356788 519044 356794
rect 518992 356730 519044 356736
rect 518912 354646 519032 354674
rect 519004 343777 519032 354646
rect 518990 343768 519046 343777
rect 518990 343703 519046 343712
rect 518898 284744 518954 284753
rect 518898 284679 518954 284688
rect 517888 262948 517940 262954
rect 517888 262890 517940 262896
rect 517888 240984 517940 240990
rect 517888 240926 517940 240932
rect 517796 240848 517848 240854
rect 517796 240790 517848 240796
rect 517704 131028 517756 131034
rect 517704 130970 517756 130976
rect 517808 130966 517836 240790
rect 517900 152522 517928 240926
rect 518912 174321 518940 284679
rect 519004 234569 519032 343703
rect 519082 281480 519138 281489
rect 519082 281415 519138 281424
rect 518990 234560 519046 234569
rect 518990 234495 519046 234504
rect 518898 174312 518954 174321
rect 518898 174247 518954 174256
rect 517888 152516 517940 152522
rect 517888 152458 517940 152464
rect 517796 130960 517848 130966
rect 517796 130902 517848 130908
rect 517612 130484 517664 130490
rect 517612 130426 517664 130432
rect 517624 42770 517652 130426
rect 518912 64841 518940 174247
rect 519096 171329 519124 281415
rect 519174 279848 519230 279857
rect 519174 279783 519230 279792
rect 519082 171320 519138 171329
rect 519082 171255 519138 171264
rect 519096 171134 519124 171255
rect 519004 171106 519124 171134
rect 518898 64832 518954 64841
rect 518898 64767 518954 64776
rect 519004 61985 519032 171106
rect 519082 169824 519138 169833
rect 519188 169810 519216 279783
rect 519280 278633 519308 358022
rect 519372 284753 519400 359518
rect 519358 284744 519414 284753
rect 519358 284679 519414 284688
rect 519464 282713 519492 364306
rect 519636 360868 519688 360874
rect 519636 360810 519688 360816
rect 519544 356788 519596 356794
rect 519544 356730 519596 356736
rect 519450 282704 519506 282713
rect 519450 282639 519506 282648
rect 519266 278624 519322 278633
rect 519266 278559 519322 278568
rect 519138 169782 519216 169810
rect 519082 169759 519138 169768
rect 518990 61976 519046 61985
rect 518990 61911 519046 61920
rect 519096 60489 519124 169759
rect 519280 169017 519308 278559
rect 519358 234560 519414 234569
rect 519358 234495 519414 234504
rect 519266 169008 519322 169017
rect 519266 168943 519322 168952
rect 519082 60480 519138 60489
rect 519082 60415 519138 60424
rect 519280 59265 519308 168943
rect 519372 124137 519400 234495
rect 519464 172689 519492 282639
rect 519556 281489 519584 356730
rect 519542 281480 519598 281489
rect 519542 281415 519598 281424
rect 519648 279857 519676 360810
rect 540256 339454 540284 502318
rect 578896 390425 578924 529178
rect 580920 518401 580948 569463
rect 580906 518392 580962 518401
rect 580906 518327 580962 518336
rect 580172 494012 580224 494018
rect 580172 493954 580224 493960
rect 580184 492833 580212 493954
rect 580170 492824 580226 492833
rect 580170 492759 580226 492768
rect 580920 467129 580948 518327
rect 580906 467120 580962 467129
rect 580906 467055 580962 467064
rect 579896 441584 579948 441590
rect 579894 441552 579896 441561
rect 579948 441552 579950 441561
rect 579894 441487 579950 441496
rect 580920 415993 580948 467055
rect 580906 415984 580962 415993
rect 580906 415919 580962 415928
rect 578882 390416 578938 390425
rect 578882 390351 578938 390360
rect 580920 364857 580948 415919
rect 580906 364848 580962 364857
rect 580906 364783 580962 364792
rect 540244 339448 540296 339454
rect 540244 339390 540296 339396
rect 580172 339448 580224 339454
rect 580172 339390 580224 339396
rect 580184 339153 580212 339390
rect 580170 339144 580226 339153
rect 580170 339079 580226 339088
rect 580920 313585 580948 364783
rect 580906 313576 580962 313585
rect 580906 313511 580962 313520
rect 519634 279848 519690 279857
rect 519634 279783 519690 279792
rect 580920 262449 580948 313511
rect 580906 262440 580962 262449
rect 580906 262375 580962 262384
rect 580920 223961 580948 262375
rect 580906 223952 580962 223961
rect 580906 223887 580962 223896
rect 580920 185609 580948 223887
rect 580906 185600 580962 185609
rect 580906 185535 580962 185544
rect 519450 172680 519506 172689
rect 519450 172615 519506 172624
rect 519358 124128 519414 124137
rect 519358 124063 519414 124072
rect 519464 63345 519492 172615
rect 580920 147257 580948 185535
rect 580906 147248 580962 147257
rect 580906 147183 580962 147192
rect 580906 108760 580962 108769
rect 580906 108695 580962 108704
rect 580920 70417 580948 108695
rect 580906 70408 580962 70417
rect 580906 70343 580962 70352
rect 519450 63336 519506 63345
rect 519450 63271 519506 63280
rect 519266 59256 519322 59265
rect 519266 59191 519322 59200
rect 517612 42764 517664 42770
rect 517612 42706 517664 42712
rect 453396 42696 453448 42702
rect 453396 42638 453448 42644
rect 503536 42696 503588 42702
rect 503536 42638 503588 42644
rect 517520 42696 517572 42702
rect 517520 42638 517572 42644
rect 448244 42628 448296 42634
rect 448244 42570 448296 42576
rect 445852 42560 445904 42566
rect 445852 42502 445904 42508
rect 443460 42492 443512 42498
rect 443460 42434 443512 42440
rect 440884 42356 440936 42362
rect 440884 42298 440936 42304
rect 438492 42288 438544 42294
rect 438492 42230 438544 42236
rect 436376 39976 436428 39982
rect 436376 39918 436428 39924
rect 375012 39432 375064 39438
rect 375012 39374 375064 39380
rect 435180 39432 435232 39438
rect 435180 39374 435232 39380
rect 274732 39364 274784 39370
rect 274732 39306 274784 39312
rect 212356 39296 212408 39302
rect 212356 39238 212408 39244
rect 273536 39296 273588 39302
rect 273536 39238 273588 39244
rect 580920 32065 580948 70343
rect 580446 32056 580502 32065
rect 580446 31991 580502 32000
rect 580906 32056 580962 32065
rect 580906 31991 580962 32000
rect 580460 31754 580488 31991
rect 580448 31748 580500 31754
rect 580448 31690 580500 31696
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6338 -960 6450 480
rect 7534 -960 7646 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12226 -960 12338 480
rect 13422 -960 13534 480
rect 14618 -960 14730 480
rect 15814 -960 15926 480
rect 17010 -960 17122 480
rect 18114 -960 18226 480
rect 19310 -960 19422 480
rect 20506 -960 20618 480
rect 21702 -960 21814 480
rect 22898 -960 23010 480
rect 24002 -960 24114 480
rect 25198 -960 25310 480
rect 26394 -960 26506 480
rect 27590 -960 27702 480
rect 28786 -960 28898 480
rect 29890 -960 30002 480
rect 31086 -960 31198 480
rect 32282 -960 32394 480
rect 33478 -960 33590 480
rect 34674 -960 34786 480
rect 35778 -960 35890 480
rect 36974 -960 37086 480
rect 38170 -960 38282 480
rect 39366 -960 39478 480
rect 40562 -960 40674 480
rect 41666 -960 41778 480
rect 42862 -960 42974 480
rect 44058 -960 44170 480
rect 45254 -960 45366 480
rect 46450 -960 46562 480
rect 47554 -960 47666 480
rect 48750 -960 48862 480
rect 49946 -960 50058 480
rect 51142 -960 51254 480
rect 52338 -960 52450 480
rect 53442 -960 53554 480
rect 54638 -960 54750 480
rect 55834 -960 55946 480
rect 57030 -960 57142 480
rect 58226 -960 58338 480
rect 59330 -960 59442 480
rect 60526 -960 60638 480
rect 61722 -960 61834 480
rect 62918 -960 63030 480
rect 64114 -960 64226 480
rect 65218 -960 65330 480
rect 66414 -960 66526 480
rect 67610 -960 67722 480
rect 68806 -960 68918 480
rect 70002 -960 70114 480
rect 71106 -960 71218 480
rect 72302 -960 72414 480
rect 73498 -960 73610 480
rect 74694 -960 74806 480
rect 75890 -960 76002 480
rect 76994 -960 77106 480
rect 78190 -960 78302 480
rect 79386 -960 79498 480
rect 80582 -960 80694 480
rect 81778 -960 81890 480
rect 82882 -960 82994 480
rect 84078 -960 84190 480
rect 85274 -960 85386 480
rect 86470 -960 86582 480
rect 87666 -960 87778 480
rect 88770 -960 88882 480
rect 89966 -960 90078 480
rect 91162 -960 91274 480
rect 92358 -960 92470 480
rect 93554 -960 93666 480
rect 94658 -960 94770 480
rect 95854 -960 95966 480
rect 97050 -960 97162 480
rect 98246 -960 98358 480
rect 99442 -960 99554 480
rect 100546 -960 100658 480
rect 101742 -960 101854 480
rect 102938 -960 103050 480
rect 104134 -960 104246 480
rect 105330 -960 105442 480
rect 106434 -960 106546 480
rect 107630 -960 107742 480
rect 108826 -960 108938 480
rect 110022 -960 110134 480
rect 111218 -960 111330 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124098 -960 124210 480
rect 125294 -960 125406 480
rect 126490 -960 126602 480
rect 127686 -960 127798 480
rect 128882 -960 128994 480
rect 129986 -960 130098 480
rect 131182 -960 131294 480
rect 132378 -960 132490 480
rect 133574 -960 133686 480
rect 134770 -960 134882 480
rect 135874 -960 135986 480
rect 137070 -960 137182 480
rect 138266 -960 138378 480
rect 139462 -960 139574 480
rect 140658 -960 140770 480
rect 141762 -960 141874 480
rect 142958 -960 143070 480
rect 144154 -960 144266 480
rect 145350 -960 145462 480
rect 146546 -960 146658 480
rect 147650 -960 147762 480
rect 148846 -960 148958 480
rect 150042 -960 150154 480
rect 151238 -960 151350 480
rect 152342 -960 152454 480
rect 153538 -960 153650 480
rect 154734 -960 154846 480
rect 155930 -960 156042 480
rect 157126 -960 157238 480
rect 158230 -960 158342 480
rect 159426 -960 159538 480
rect 160622 -960 160734 480
rect 161818 -960 161930 480
rect 163014 -960 163126 480
rect 164118 -960 164230 480
rect 165314 -960 165426 480
rect 166510 -960 166622 480
rect 167706 -960 167818 480
rect 168902 -960 169014 480
rect 170006 -960 170118 480
rect 171202 -960 171314 480
rect 172398 -960 172510 480
rect 173594 -960 173706 480
rect 174790 -960 174902 480
rect 175894 -960 176006 480
rect 177090 -960 177202 480
rect 178286 -960 178398 480
rect 179482 -960 179594 480
rect 180678 -960 180790 480
rect 181782 -960 181894 480
rect 182978 -960 183090 480
rect 184174 -960 184286 480
rect 185370 -960 185482 480
rect 186566 -960 186678 480
rect 187670 -960 187782 480
rect 188866 -960 188978 480
rect 190062 -960 190174 480
rect 191258 -960 191370 480
rect 192454 -960 192566 480
rect 193558 -960 193670 480
rect 194754 -960 194866 480
rect 195950 -960 196062 480
rect 197146 -960 197258 480
rect 198342 -960 198454 480
rect 199446 -960 199558 480
rect 200642 -960 200754 480
rect 201838 -960 201950 480
rect 203034 -960 203146 480
rect 204230 -960 204342 480
rect 205334 -960 205446 480
rect 206530 -960 206642 480
rect 207726 -960 207838 480
rect 208922 -960 209034 480
rect 210118 -960 210230 480
rect 211222 -960 211334 480
rect 212418 -960 212530 480
rect 213614 -960 213726 480
rect 214810 -960 214922 480
rect 216006 -960 216118 480
rect 217110 -960 217222 480
rect 218306 -960 218418 480
rect 219502 -960 219614 480
rect 220698 -960 220810 480
rect 221894 -960 222006 480
rect 222998 -960 223110 480
rect 224194 -960 224306 480
rect 225390 -960 225502 480
rect 226586 -960 226698 480
rect 227782 -960 227894 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240662 -960 240774 480
rect 241858 -960 241970 480
rect 243054 -960 243166 480
rect 244250 -960 244362 480
rect 245446 -960 245558 480
rect 246550 -960 246662 480
rect 247746 -960 247858 480
rect 248942 -960 249054 480
rect 250138 -960 250250 480
rect 251334 -960 251446 480
rect 252438 -960 252550 480
rect 253634 -960 253746 480
rect 254830 -960 254942 480
rect 256026 -960 256138 480
rect 257222 -960 257334 480
rect 258326 -960 258438 480
rect 259522 -960 259634 480
rect 260718 -960 260830 480
rect 261914 -960 262026 480
rect 263110 -960 263222 480
rect 264214 -960 264326 480
rect 265410 -960 265522 480
rect 266606 -960 266718 480
rect 267802 -960 267914 480
rect 268998 -960 269110 480
rect 270102 -960 270214 480
rect 271298 -960 271410 480
rect 272494 -960 272606 480
rect 273690 -960 273802 480
rect 274886 -960 274998 480
rect 275990 -960 276102 480
rect 277186 -960 277298 480
rect 278382 -960 278494 480
rect 279578 -960 279690 480
rect 280774 -960 280886 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285466 -960 285578 480
rect 286662 -960 286774 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298346 -960 298458 480
rect 299542 -960 299654 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304234 -960 304346 480
rect 305430 -960 305542 480
rect 306626 -960 306738 480
rect 307822 -960 307934 480
rect 309018 -960 309130 480
rect 310122 -960 310234 480
rect 311318 -960 311430 480
rect 312514 -960 312626 480
rect 313710 -960 313822 480
rect 314906 -960 315018 480
rect 316010 -960 316122 480
rect 317206 -960 317318 480
rect 318402 -960 318514 480
rect 319598 -960 319710 480
rect 320794 -960 320906 480
rect 321898 -960 322010 480
rect 323094 -960 323206 480
rect 324290 -960 324402 480
rect 325486 -960 325598 480
rect 326682 -960 326794 480
rect 327786 -960 327898 480
rect 328982 -960 329094 480
rect 330178 -960 330290 480
rect 331374 -960 331486 480
rect 332570 -960 332682 480
rect 333674 -960 333786 480
rect 334870 -960 334982 480
rect 336066 -960 336178 480
rect 337262 -960 337374 480
rect 338458 -960 338570 480
rect 339562 -960 339674 480
rect 340758 -960 340870 480
rect 341954 -960 342066 480
rect 343150 -960 343262 480
rect 344346 -960 344458 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357226 -960 357338 480
rect 358422 -960 358534 480
rect 359618 -960 359730 480
rect 360814 -960 360926 480
rect 362010 -960 362122 480
rect 363114 -960 363226 480
rect 364310 -960 364422 480
rect 365506 -960 365618 480
rect 366702 -960 366814 480
rect 367898 -960 368010 480
rect 369002 -960 369114 480
rect 370198 -960 370310 480
rect 371394 -960 371506 480
rect 372590 -960 372702 480
rect 373786 -960 373898 480
rect 374890 -960 375002 480
rect 376086 -960 376198 480
rect 377282 -960 377394 480
rect 378478 -960 378590 480
rect 379674 -960 379786 480
rect 380778 -960 380890 480
rect 381974 -960 382086 480
rect 383170 -960 383282 480
rect 384366 -960 384478 480
rect 385562 -960 385674 480
rect 386666 -960 386778 480
rect 387862 -960 387974 480
rect 389058 -960 389170 480
rect 390254 -960 390366 480
rect 391450 -960 391562 480
rect 392554 -960 392666 480
rect 393750 -960 393862 480
rect 394946 -960 395058 480
rect 396142 -960 396254 480
rect 397338 -960 397450 480
rect 398442 -960 398554 480
rect 399638 -960 399750 480
rect 400834 -960 400946 480
rect 402030 -960 402142 480
rect 403226 -960 403338 480
rect 404330 -960 404442 480
rect 405526 -960 405638 480
rect 406722 -960 406834 480
rect 407918 -960 408030 480
rect 409114 -960 409226 480
rect 410218 -960 410330 480
rect 411414 -960 411526 480
rect 412610 -960 412722 480
rect 413806 -960 413918 480
rect 415002 -960 415114 480
rect 416106 -960 416218 480
rect 417302 -960 417414 480
rect 418498 -960 418610 480
rect 419694 -960 419806 480
rect 420890 -960 421002 480
rect 421994 -960 422106 480
rect 423190 -960 423302 480
rect 424386 -960 424498 480
rect 425582 -960 425694 480
rect 426778 -960 426890 480
rect 427882 -960 427994 480
rect 429078 -960 429190 480
rect 430274 -960 430386 480
rect 431470 -960 431582 480
rect 432666 -960 432778 480
rect 433770 -960 433882 480
rect 434966 -960 435078 480
rect 436162 -960 436274 480
rect 437358 -960 437470 480
rect 438554 -960 438666 480
rect 439658 -960 439770 480
rect 440854 -960 440966 480
rect 442050 -960 442162 480
rect 443246 -960 443358 480
rect 444350 -960 444462 480
rect 445546 -960 445658 480
rect 446742 -960 446854 480
rect 447938 -960 448050 480
rect 449134 -960 449246 480
rect 450238 -960 450350 480
rect 451434 -960 451546 480
rect 452630 -960 452742 480
rect 453826 -960 453938 480
rect 455022 -960 455134 480
rect 456126 -960 456238 480
rect 457322 -960 457434 480
rect 458518 -960 458630 480
rect 459714 -960 459826 480
rect 460910 -960 461022 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473790 -960 473902 480
rect 474986 -960 475098 480
rect 476182 -960 476294 480
rect 477378 -960 477490 480
rect 478574 -960 478686 480
rect 479678 -960 479790 480
rect 480874 -960 480986 480
rect 482070 -960 482182 480
rect 483266 -960 483378 480
rect 484462 -960 484574 480
rect 485566 -960 485678 480
rect 486762 -960 486874 480
rect 487958 -960 488070 480
rect 489154 -960 489266 480
rect 490350 -960 490462 480
rect 491454 -960 491566 480
rect 492650 -960 492762 480
rect 493846 -960 493958 480
rect 495042 -960 495154 480
rect 496238 -960 496350 480
rect 497342 -960 497454 480
rect 498538 -960 498650 480
rect 499734 -960 499846 480
rect 500930 -960 501042 480
rect 502126 -960 502238 480
rect 503230 -960 503342 480
rect 504426 -960 504538 480
rect 505622 -960 505734 480
rect 506818 -960 506930 480
rect 508014 -960 508126 480
rect 509118 -960 509230 480
rect 510314 -960 510426 480
rect 511510 -960 511622 480
rect 512706 -960 512818 480
rect 513902 -960 514014 480
rect 515006 -960 515118 480
rect 516202 -960 516314 480
rect 517398 -960 517510 480
rect 518594 -960 518706 480
rect 519790 -960 519902 480
rect 520894 -960 521006 480
rect 522090 -960 522202 480
rect 523286 -960 523398 480
rect 524482 -960 524594 480
rect 525678 -960 525790 480
rect 526782 -960 526894 480
rect 527978 -960 528090 480
rect 529174 -960 529286 480
rect 530370 -960 530482 480
rect 531566 -960 531678 480
rect 532670 -960 532782 480
rect 533866 -960 533978 480
rect 535062 -960 535174 480
rect 536258 -960 536370 480
rect 537454 -960 537566 480
rect 538558 -960 538670 480
rect 539754 -960 539866 480
rect 540950 -960 541062 480
rect 542146 -960 542258 480
rect 543342 -960 543454 480
rect 544446 -960 544558 480
rect 545642 -960 545754 480
rect 546838 -960 546950 480
rect 548034 -960 548146 480
rect 549230 -960 549342 480
rect 550334 -960 550446 480
rect 551530 -960 551642 480
rect 552726 -960 552838 480
rect 553922 -960 554034 480
rect 555118 -960 555230 480
rect 556222 -960 556334 480
rect 557418 -960 557530 480
rect 558614 -960 558726 480
rect 559810 -960 559922 480
rect 561006 -960 561118 480
rect 562110 -960 562222 480
rect 563306 -960 563418 480
rect 564502 -960 564614 480
rect 565698 -960 565810 480
rect 566894 -960 567006 480
rect 567998 -960 568110 480
rect 569194 -960 569306 480
rect 570390 -960 570502 480
rect 571586 -960 571698 480
rect 572782 -960 572894 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577474 -960 577586 480
rect 578670 -960 578782 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 685072 3478 685128
rect 2778 659912 2834 659968
rect 3422 634752 3478 634808
rect 2778 609592 2834 609648
rect 3514 584432 3570 584488
rect 2778 559272 2834 559328
rect 3422 554784 3478 554840
rect 3422 521600 3478 521656
rect 2778 509088 2834 509144
rect 3514 471280 3570 471336
rect 2778 458768 2834 458824
rect 3146 421096 3202 421152
rect 2778 408448 2834 408504
rect 2778 358264 2834 358320
rect 2778 307944 2834 308000
rect 2778 257624 2834 257680
rect 2778 207304 2834 207360
rect 2870 169668 2872 169688
rect 2872 169668 2924 169688
rect 2924 169668 2926 169688
rect 2870 169632 2926 169668
rect 2778 157120 2834 157176
rect 2962 119312 3018 119368
rect 2778 106800 2834 106856
rect 3514 370776 3570 370832
rect 3422 81640 3478 81696
rect 2778 69128 2834 69184
rect 57426 635568 57482 635624
rect 57242 602248 57298 602304
rect 57150 586608 57206 586664
rect 57058 580488 57114 580544
rect 57702 629448 57758 629504
rect 57610 626728 57666 626784
rect 57518 608368 57574 608424
rect 57334 598848 57390 598904
rect 57426 596128 57482 596184
rect 59082 632848 59138 632904
rect 58898 623328 58954 623384
rect 58530 617208 58586 617264
rect 57886 611088 57942 611144
rect 58438 590008 58494 590064
rect 58806 604968 58862 605024
rect 58714 583888 58770 583944
rect 58990 620608 59046 620664
rect 59266 614488 59322 614544
rect 59266 592728 59322 592784
rect 59542 577732 59598 577788
rect 120998 597624 121054 597680
rect 121090 579808 121146 579864
rect 121182 577088 121238 577144
rect 121550 589328 121606 589384
rect 122194 628768 122250 628824
rect 121826 626048 121882 626104
rect 121734 622648 121790 622704
rect 121918 619928 121974 619984
rect 122010 613808 122066 613864
rect 122102 595448 122158 595504
rect 122286 585928 122342 585984
rect 122930 634888 122986 634944
rect 123022 632168 123078 632224
rect 123206 616528 123262 616584
rect 123114 610408 123170 610464
rect 123298 607688 123354 607744
rect 124126 604288 124182 604344
rect 123390 601568 123446 601624
rect 123482 592048 123538 592104
rect 123574 583208 123630 583264
rect 137282 635568 137338 635624
rect 136638 623328 136694 623384
rect 137098 620608 137154 620664
rect 137006 617208 137062 617264
rect 136638 592728 136694 592784
rect 136638 590008 136694 590064
rect 137558 614488 137614 614544
rect 137282 611088 137338 611144
rect 137374 604968 137430 605024
rect 137374 602248 137430 602304
rect 137466 596128 137522 596184
rect 137742 629448 137798 629504
rect 137926 611088 137982 611144
rect 137926 583888 137982 583944
rect 138570 580488 138626 580544
rect 138478 577768 138534 577824
rect 139122 632848 139178 632904
rect 139030 626728 139086 626784
rect 138938 608368 138994 608424
rect 138846 598848 138902 598904
rect 139306 586608 139362 586664
rect 200762 613264 200818 613320
rect 201038 592048 201094 592104
rect 201130 583208 201186 583264
rect 201222 577088 201278 577144
rect 201590 634888 201646 634944
rect 201774 632168 201830 632224
rect 201682 628768 201738 628824
rect 201958 626048 202014 626104
rect 201866 619928 201922 619984
rect 202970 622648 203026 622704
rect 202878 607688 202934 607744
rect 202142 601568 202198 601624
rect 202050 595448 202106 595504
rect 202234 585928 202290 585984
rect 203154 616528 203210 616584
rect 203062 610408 203118 610464
rect 203890 604288 203946 604344
rect 203246 598168 203302 598224
rect 203338 589328 203394 589384
rect 203430 579808 203486 579864
rect 216678 635568 216734 635624
rect 216678 632848 216734 632904
rect 216678 626728 216734 626784
rect 216678 623328 216734 623384
rect 216678 604968 216734 605024
rect 216678 602248 216734 602304
rect 216678 592728 216734 592784
rect 216678 590008 216734 590064
rect 216678 586608 216734 586664
rect 216678 577768 216734 577824
rect 217046 598848 217102 598904
rect 217690 629448 217746 629504
rect 217598 617208 217654 617264
rect 217414 608368 217470 608424
rect 217782 614488 217838 614544
rect 217782 596128 217838 596184
rect 217598 557504 217654 557560
rect 218702 611088 218758 611144
rect 218150 580488 218206 580544
rect 217966 557504 218022 557560
rect 219254 620608 219310 620664
rect 219162 583888 219218 583944
rect 241518 556144 241574 556200
rect 248694 556688 248750 556744
rect 255134 556416 255190 556472
rect 258722 556552 258778 556608
rect 280894 610000 280950 610056
rect 281078 647264 281134 647320
rect 281630 634888 281686 634944
rect 281170 589328 281226 589384
rect 282090 632168 282146 632224
rect 281722 626048 281778 626104
rect 281630 583208 281686 583264
rect 281262 579808 281318 579864
rect 281538 577088 281594 577144
rect 281906 601568 281962 601624
rect 281814 595448 281870 595504
rect 281998 598168 282054 598224
rect 283470 628768 283526 628824
rect 283010 622648 283066 622704
rect 282918 592048 282974 592104
rect 283378 619928 283434 619984
rect 283286 616528 283342 616584
rect 283102 613808 283158 613864
rect 283194 607688 283250 607744
rect 283654 604288 283710 604344
rect 283562 585928 283618 585984
rect 290922 556280 290978 556336
rect 300674 556688 300730 556744
rect 300490 556416 300546 556472
rect 302330 532480 302386 532536
rect 303158 556552 303214 556608
rect 303250 547440 303306 547496
rect 303158 535472 303214 535528
rect 57702 525036 57704 525056
rect 57704 525036 57756 525056
rect 57756 525036 57758 525056
rect 42338 486376 42394 486432
rect 3422 44004 3424 44024
rect 3424 44004 3476 44024
rect 3476 44004 3478 44024
rect 3422 43968 3478 44004
rect 57702 525000 57758 525036
rect 309782 647400 309838 647456
rect 302974 517520 303030 517576
rect 302882 502560 302938 502616
rect 43718 486784 43774 486840
rect 43810 486648 43866 486704
rect 46846 489096 46902 489152
rect 46570 263200 46626 263256
rect 46478 260344 46534 260400
rect 46386 260072 46442 260128
rect 46754 486512 46810 486568
rect 48226 263064 48282 263120
rect 49054 489232 49110 489288
rect 48962 263336 49018 263392
rect 49054 262792 49110 262848
rect 50526 491272 50582 491328
rect 49422 462984 49478 463040
rect 49330 462848 49386 462904
rect 49238 459584 49294 459640
rect 49606 380976 49662 381032
rect 49422 152904 49478 152960
rect 49330 152632 49386 152688
rect 50526 489504 50582 489560
rect 50434 260752 50490 260808
rect 50618 489368 50674 489424
rect 50434 260208 50490 260264
rect 50434 130600 50490 130656
rect 50802 373904 50858 373960
rect 50986 459584 51042 459640
rect 50986 375264 51042 375320
rect 51078 374992 51134 375048
rect 51446 263608 51502 263664
rect 52366 491272 52422 491328
rect 51630 132368 51686 132424
rect 52182 465976 52238 466032
rect 52274 459584 52330 459640
rect 52274 372680 52330 372736
rect 52918 319912 52974 319968
rect 53562 466248 53618 466304
rect 53470 459584 53526 459640
rect 53010 130872 53066 130928
rect 53654 466112 53710 466168
rect 54390 129648 54446 129704
rect 54298 129512 54354 129568
rect 55494 459584 55550 459640
rect 56230 372680 56286 372736
rect 56046 131008 56102 131064
rect 56138 130872 56194 130928
rect 56138 130464 56194 130520
rect 56874 383016 56930 383072
rect 57242 412392 57298 412448
rect 57242 411204 57244 411224
rect 57244 411204 57296 411224
rect 57296 411204 57298 411224
rect 57242 411168 57298 411204
rect 57242 408584 57298 408640
rect 57242 407224 57298 407280
rect 57242 405748 57298 405784
rect 57242 405728 57244 405748
rect 57244 405728 57296 405748
rect 57296 405728 57298 405748
rect 57242 404388 57298 404424
rect 57242 404368 57244 404388
rect 57244 404368 57296 404388
rect 57296 404368 57298 404388
rect 57242 403028 57298 403064
rect 57242 403008 57244 403028
rect 57244 403008 57296 403028
rect 57296 403008 57298 403028
rect 57242 384956 57244 384976
rect 57244 384956 57296 384976
rect 57296 384956 57298 384976
rect 57242 384920 57298 384956
rect 56782 301688 56838 301744
rect 56598 300872 56654 300928
rect 56690 293936 56746 293992
rect 56598 191664 56654 191720
rect 56874 264152 56930 264208
rect 56782 193160 56838 193216
rect 56782 191664 56838 191720
rect 56782 190848 56838 190904
rect 56690 185408 56746 185464
rect 56874 187856 56930 187912
rect 56782 81368 56838 81424
rect 57518 383288 57574 383344
rect 57426 297744 57482 297800
rect 57334 294888 57390 294944
rect 57334 293936 57390 293992
rect 57334 292576 57390 292632
rect 57242 273264 57298 273320
rect 57150 237360 57206 237416
rect 57150 185680 57206 185736
rect 57058 183504 57114 183560
rect 56966 133764 56968 133784
rect 56968 133764 57020 133784
rect 57020 133764 57022 133784
rect 56966 133728 57022 133764
rect 56874 78376 56930 78432
rect 57610 301688 57666 301744
rect 57702 300872 57758 300928
rect 57702 299376 57758 299432
rect 57518 295976 57574 296032
rect 57426 187856 57482 187912
rect 57334 187720 57390 187776
rect 57610 275576 57666 275632
rect 57610 193160 57666 193216
rect 57610 191800 57666 191856
rect 57518 185680 57574 185736
rect 57426 183504 57482 183560
rect 57334 79328 57390 79384
rect 57150 76608 57206 76664
rect 57886 299376 57942 299432
rect 57886 273264 57942 273320
rect 57702 188672 57758 188728
rect 57702 187720 57758 187776
rect 57702 185408 57758 185464
rect 57610 82456 57666 82512
rect 58622 264832 58678 264888
rect 58990 272992 59046 273048
rect 57886 163240 57942 163296
rect 57794 150456 57850 150512
rect 57702 75520 57758 75576
rect 57426 73752 57482 73808
rect 2778 31320 2834 31376
rect 58622 237360 58678 237416
rect 58898 238584 58954 238640
rect 58898 237360 58954 237416
rect 57978 131008 58034 131064
rect 57886 53352 57942 53408
rect 59082 165552 59138 165608
rect 60002 465840 60058 465896
rect 59818 262656 59874 262712
rect 58990 130600 59046 130656
rect 66166 492224 66222 492280
rect 68926 492260 68928 492280
rect 68928 492260 68980 492280
rect 68980 492260 68982 492280
rect 68926 492224 68982 492260
rect 68650 491680 68706 491736
rect 69018 460808 69074 460864
rect 69202 463392 69258 463448
rect 69110 460536 69166 460592
rect 70490 463256 70546 463312
rect 71778 460672 71834 460728
rect 72882 492496 72938 492552
rect 71962 492360 72018 492416
rect 74262 491544 74318 491600
rect 73158 461488 73214 461544
rect 74630 460400 74686 460456
rect 76010 492088 76066 492144
rect 77758 492360 77814 492416
rect 77298 491952 77354 492008
rect 78586 492224 78642 492280
rect 76010 460264 76066 460320
rect 74722 460128 74778 460184
rect 67730 459992 67786 460048
rect 80794 491816 80850 491872
rect 81530 465704 81586 465760
rect 84382 466248 84438 466304
rect 84290 465976 84346 466032
rect 80150 463120 80206 463176
rect 85762 466112 85818 466168
rect 80058 459040 80114 459096
rect 89902 458904 89958 458960
rect 92662 465840 92718 465896
rect 93858 462984 93914 463040
rect 93950 462848 94006 462904
rect 107658 462848 107714 462904
rect 115662 489504 115718 489560
rect 120354 489640 120410 489696
rect 120262 489368 120318 489424
rect 120170 489232 120226 489288
rect 121458 486920 121514 486976
rect 121642 486784 121698 486840
rect 123022 486648 123078 486704
rect 122838 483928 122894 483984
rect 125782 489096 125838 489152
rect 125690 483792 125746 483848
rect 127070 486512 127126 486568
rect 127162 486376 127218 486432
rect 126978 483656 127034 483712
rect 129646 487736 129702 487792
rect 145102 491816 145158 491872
rect 143722 486376 143778 486432
rect 143538 478080 143594 478136
rect 145010 483656 145066 483712
rect 146574 491952 146630 492008
rect 147770 492224 147826 492280
rect 146298 475360 146354 475416
rect 144918 472504 144974 472560
rect 149150 492088 149206 492144
rect 150254 492360 150310 492416
rect 147770 486512 147826 486568
rect 147678 465704 147734 465760
rect 153750 490456 153806 490512
rect 150530 479440 150586 479496
rect 151818 476720 151874 476776
rect 153198 475496 153254 475552
rect 156050 469784 156106 469840
rect 155958 468424 156014 468480
rect 154578 460264 154634 460320
rect 157430 474000 157486 474056
rect 160282 465840 160338 465896
rect 158718 463120 158774 463176
rect 157338 460128 157394 460184
rect 161570 461488 161626 461544
rect 161478 459040 161534 459096
rect 164330 469920 164386 469976
rect 166998 460400 167054 460456
rect 169850 465976 169906 466032
rect 169758 463256 169814 463312
rect 169942 462984 169998 463040
rect 171414 489096 171470 489152
rect 171322 461624 171378 461680
rect 172702 467064 172758 467120
rect 172518 459312 172574 459368
rect 171138 459176 171194 459232
rect 178314 461352 178370 461408
rect 179602 478216 179658 478272
rect 180062 462168 180118 462224
rect 185766 492496 185822 492552
rect 183650 463392 183706 463448
rect 187054 491680 187110 491736
rect 186318 459448 186374 459504
rect 162858 458904 162914 458960
rect 91282 458768 91338 458824
rect 150438 458768 150494 458824
rect 191194 492224 191250 492280
rect 191194 491408 191250 491464
rect 190918 460964 190974 461000
rect 190918 460944 190920 460964
rect 190920 460944 190972 460964
rect 190972 460944 190974 460964
rect 105450 374992 105506 375048
rect 140962 374856 141018 374912
rect 163410 374584 163466 374640
rect 165986 374604 166042 374640
rect 165986 374584 165988 374604
rect 165988 374584 166040 374604
rect 166040 374584 166042 374604
rect 179326 374584 179382 374640
rect 143538 374448 143594 374504
rect 153474 374448 153530 374504
rect 158534 374468 158590 374504
rect 158534 374448 158536 374468
rect 158536 374448 158588 374468
rect 158588 374448 158590 374468
rect 148966 374312 149022 374368
rect 160926 374448 160982 374504
rect 146206 374196 146262 374232
rect 146206 374176 146208 374196
rect 146208 374176 146260 374196
rect 146260 374176 146262 374196
rect 98366 373768 98422 373824
rect 103518 373804 103520 373824
rect 103520 373804 103572 373824
rect 103572 373804 103574 373824
rect 103518 373768 103574 373804
rect 110418 373768 110474 373824
rect 95054 373632 95110 373688
rect 96158 373632 96214 373688
rect 90178 373360 90234 373416
rect 96066 373380 96122 373416
rect 98274 373496 98330 373552
rect 113546 373632 113602 373688
rect 116122 373632 116178 373688
rect 118330 373668 118332 373688
rect 118332 373668 118384 373688
rect 118384 373668 118386 373688
rect 118330 373632 118386 373668
rect 121366 373632 121422 373688
rect 124126 373632 124182 373688
rect 125690 373652 125746 373688
rect 125690 373632 125692 373652
rect 125692 373632 125744 373652
rect 125744 373632 125746 373652
rect 107842 373516 107898 373552
rect 128910 373668 128912 373688
rect 128912 373668 128964 373688
rect 128964 373668 128966 373688
rect 128910 373632 128966 373668
rect 131026 373632 131082 373688
rect 133694 373652 133750 373688
rect 133694 373632 133696 373652
rect 133696 373632 133748 373652
rect 133748 373632 133750 373652
rect 136454 373632 136510 373688
rect 139214 373632 139270 373688
rect 151726 373632 151782 373688
rect 107842 373496 107844 373516
rect 107844 373496 107896 373516
rect 107896 373496 107898 373516
rect 96066 373360 96068 373380
rect 96068 373360 96120 373380
rect 96120 373360 96122 373380
rect 88338 373224 88394 373280
rect 100850 373244 100906 373280
rect 156510 373496 156566 373552
rect 100850 373224 100852 373244
rect 100852 373224 100904 373244
rect 100904 373224 100906 373244
rect 92386 373088 92442 373144
rect 93674 373108 93730 373144
rect 93674 373088 93676 373108
rect 93676 373088 93728 373108
rect 93728 373088 93730 373108
rect 84750 372564 84806 372600
rect 84750 372544 84752 372564
rect 84752 372544 84804 372564
rect 84804 372544 84806 372564
rect 86774 372544 86830 372600
rect 88062 372544 88118 372600
rect 89350 372544 89406 372600
rect 90914 372544 90970 372600
rect 91558 372544 91614 372600
rect 79506 372408 79562 372464
rect 84566 372408 84622 372464
rect 78310 372272 78366 372328
rect 76838 371728 76894 371784
rect 77206 371728 77262 371784
rect 81438 372000 81494 372056
rect 80058 371356 80060 371376
rect 80060 371356 80112 371376
rect 80112 371356 80114 371376
rect 80058 371320 80114 371356
rect 83830 371456 83886 371512
rect 93398 372544 93454 372600
rect 100022 372544 100078 372600
rect 104622 372544 104678 372600
rect 112994 372544 113050 372600
rect 114466 372544 114522 372600
rect 102046 371592 102102 371648
rect 101678 371320 101734 371376
rect 102782 371320 102838 371376
rect 110142 372272 110198 372328
rect 107014 371592 107070 371648
rect 108854 371592 108910 371648
rect 105634 371320 105690 371376
rect 111614 371592 111670 371648
rect 110142 370504 110198 370560
rect 107014 369008 107070 369064
rect 182730 372408 182786 372464
rect 183282 371864 183338 371920
rect 179326 351908 179328 351928
rect 179328 351908 179380 351928
rect 179380 351908 179382 351928
rect 179326 351872 179382 351908
rect 179694 350548 179696 350568
rect 179696 350548 179748 350568
rect 179748 350548 179750 350568
rect 179694 350512 179750 350548
rect 191286 350512 191342 350568
rect 196622 350548 196624 350568
rect 196624 350548 196676 350568
rect 196676 350548 196678 350568
rect 196622 350512 196678 350548
rect 110970 264868 110972 264888
rect 110972 264868 111024 264888
rect 111024 264868 111026 264888
rect 110970 264832 111026 264868
rect 125966 264852 126022 264888
rect 125966 264832 125968 264852
rect 125968 264832 126020 264852
rect 126020 264832 126022 264852
rect 128358 264832 128414 264888
rect 130934 264832 130990 264888
rect 133418 264832 133474 264888
rect 135902 264832 135958 264888
rect 138478 264832 138534 264888
rect 140870 264696 140926 264752
rect 143538 264696 143594 264752
rect 145930 264696 145986 264752
rect 148506 264696 148562 264752
rect 60738 264152 60794 264208
rect 80058 263472 80114 263528
rect 88338 263472 88394 263528
rect 89994 263472 90050 263528
rect 90730 263472 90786 263528
rect 91282 263472 91338 263528
rect 92386 263472 92442 263528
rect 93582 263472 93638 263528
rect 96066 263472 96122 263528
rect 98090 263472 98146 263528
rect 101034 263472 101090 263528
rect 103518 263472 103574 263528
rect 105634 263472 105690 263528
rect 108210 263472 108266 263528
rect 109314 263472 109370 263528
rect 113362 263472 113418 263528
rect 115938 263472 115994 263528
rect 116214 263472 116270 263528
rect 118054 263472 118110 263528
rect 120906 263508 120908 263528
rect 120908 263508 120960 263528
rect 120960 263508 120962 263528
rect 120906 263472 120962 263508
rect 123482 263492 123538 263528
rect 123482 263472 123484 263492
rect 123484 263472 123536 263492
rect 123536 263472 123538 263492
rect 66258 262792 66314 262848
rect 78678 262792 78734 262848
rect 77298 262248 77354 262304
rect 81438 263200 81494 263256
rect 84750 263200 84806 263256
rect 80150 262792 80206 262848
rect 80150 260344 80206 260400
rect 82082 263064 82138 263120
rect 84198 262928 84254 262984
rect 87602 262928 87658 262984
rect 85946 262520 86002 262576
rect 88614 262928 88670 262984
rect 96526 263200 96582 263256
rect 96526 260208 96582 260264
rect 99470 263200 99526 263256
rect 97906 262248 97962 262304
rect 99286 262248 99342 262304
rect 100758 262928 100814 262984
rect 101770 262676 101826 262712
rect 101770 262656 101772 262676
rect 101772 262656 101824 262676
rect 101824 262656 101826 262676
rect 102322 262656 102378 262712
rect 105082 262656 105138 262712
rect 108026 262656 108082 262712
rect 107566 262384 107622 262440
rect 107566 262248 107622 262304
rect 114374 263336 114430 263392
rect 114650 262520 114706 262576
rect 110418 262248 110474 262304
rect 113178 262248 113234 262304
rect 150990 263472 151046 263528
rect 155958 263508 155960 263528
rect 155960 263508 156012 263528
rect 156012 263508 156014 263528
rect 155958 263472 156014 263508
rect 158534 263492 158590 263528
rect 158534 263472 158536 263492
rect 158536 263472 158588 263492
rect 158588 263472 158590 263492
rect 161110 263472 161166 263528
rect 163502 263472 163558 263528
rect 166078 263472 166134 263528
rect 118698 262928 118754 262984
rect 183466 262384 183522 262440
rect 183374 262248 183430 262304
rect 114650 260072 114706 260128
rect 197358 491544 197414 491600
rect 197634 491680 197690 491736
rect 197726 491272 197782 491328
rect 179326 240216 179382 240272
rect 180154 240216 180210 240272
rect 190918 240236 190974 240272
rect 190918 240216 190920 240236
rect 190920 240216 190972 240236
rect 190972 240216 190974 240236
rect 96066 154672 96122 154728
rect 113362 154672 113418 154728
rect 163318 154692 163374 154728
rect 163318 154672 163320 154692
rect 163320 154672 163372 154692
rect 163372 154672 163374 154692
rect 98458 154128 98514 154184
rect 101034 154128 101090 154184
rect 105818 154128 105874 154184
rect 108210 154148 108266 154184
rect 165894 154672 165950 154728
rect 138386 154264 138442 154320
rect 108210 154128 108212 154148
rect 108212 154128 108264 154148
rect 108264 154128 108266 154148
rect 143538 154128 143594 154184
rect 145930 154012 145986 154048
rect 145930 153992 145932 154012
rect 145932 153992 145984 154012
rect 145984 153992 145986 154012
rect 150898 153992 150954 154048
rect 153290 153876 153346 153912
rect 153290 153856 153292 153876
rect 153292 153856 153344 153876
rect 153344 153856 153346 153876
rect 75918 153040 75974 153096
rect 77298 153040 77354 153096
rect 78678 153040 78734 153096
rect 81438 153040 81494 153096
rect 82818 153040 82874 153096
rect 84198 153040 84254 153096
rect 85578 153040 85634 153096
rect 86958 153040 87014 153096
rect 88430 153040 88486 153096
rect 89810 153040 89866 153096
rect 91098 153040 91154 153096
rect 92478 153040 92534 153096
rect 93858 153040 93914 153096
rect 95238 153040 95294 153096
rect 96618 153040 96674 153096
rect 97998 153040 98054 153096
rect 99378 153040 99434 153096
rect 100850 153040 100906 153096
rect 102138 153040 102194 153096
rect 103610 153040 103666 153096
rect 106370 153040 106426 153096
rect 109038 153040 109094 153096
rect 110418 153040 110474 153096
rect 111154 153040 111210 153096
rect 111798 153040 111854 153096
rect 114558 153040 114614 153096
rect 76010 152496 76066 152552
rect 80058 151952 80114 152008
rect 84290 151952 84346 152008
rect 88338 152360 88394 152416
rect 88890 152768 88946 152824
rect 88890 152496 88946 152552
rect 89718 152380 89774 152416
rect 89718 152360 89720 152380
rect 89720 152360 89772 152380
rect 89772 152360 89774 152380
rect 91190 152768 91246 152824
rect 98642 133048 98698 133104
rect 97262 130600 97318 130656
rect 95238 130464 95294 130520
rect 100758 152768 100814 152824
rect 103518 152768 103574 152824
rect 106278 152768 106334 152824
rect 104898 152088 104954 152144
rect 109130 152768 109186 152824
rect 113178 152768 113234 152824
rect 114742 153040 114798 153096
rect 117318 153040 117374 153096
rect 117502 153040 117558 153096
rect 118698 153040 118754 153096
rect 125598 153040 125654 153096
rect 128358 153040 128414 153096
rect 129738 153040 129794 153096
rect 132774 153060 132830 153096
rect 132774 153040 132776 153060
rect 132776 153040 132828 153060
rect 132828 153040 132830 153060
rect 115938 152516 115994 152552
rect 115938 152496 115940 152516
rect 115940 152496 115992 152516
rect 115992 152496 115994 152516
rect 117410 152768 117466 152824
rect 135258 153076 135260 153096
rect 135260 153076 135312 153096
rect 135312 153076 135314 153096
rect 135258 153040 135314 153076
rect 155958 153040 156014 153096
rect 120078 152768 120134 152824
rect 122838 152788 122894 152824
rect 122838 152768 122840 152788
rect 122840 152768 122892 152788
rect 122892 152768 122894 152788
rect 183466 152768 183522 152824
rect 183466 152516 183522 152552
rect 183466 152496 183468 152516
rect 183468 152496 183520 152516
rect 183520 152496 183522 152516
rect 102138 131008 102194 131064
rect 99378 130328 99434 130384
rect 191746 130328 191802 130384
rect 179050 129784 179106 129840
rect 179786 129784 179842 129840
rect 77114 44784 77170 44840
rect 83094 44784 83150 44840
rect 84198 44784 84254 44840
rect 94502 44784 94558 44840
rect 96986 44784 97042 44840
rect 98090 44784 98146 44840
rect 100758 44648 100814 44704
rect 101770 44648 101826 44704
rect 102782 44648 102838 44704
rect 103886 44648 103942 44704
rect 143538 44648 143594 44704
rect 145930 44648 145986 44704
rect 113270 44512 113326 44568
rect 158442 44104 158498 44160
rect 160834 44104 160890 44160
rect 115938 43696 115994 43752
rect 85394 43152 85450 43208
rect 92386 43152 92442 43208
rect 95882 43152 95938 43208
rect 128358 43152 128414 43208
rect 76010 42744 76066 42800
rect 78218 42744 78274 42800
rect 80426 42744 80482 42800
rect 78770 41792 78826 41848
rect 81806 41792 81862 41848
rect 86498 42744 86554 42800
rect 87602 42744 87658 42800
rect 88338 42744 88394 42800
rect 88614 42744 88670 42800
rect 90730 42744 90786 42800
rect 91282 42744 91338 42800
rect 89994 41792 90050 41848
rect 93306 42744 93362 42800
rect 93674 42744 93730 42800
rect 96250 42744 96306 42800
rect 106370 42744 106426 42800
rect 107014 42744 107070 42800
rect 108578 42744 108634 42800
rect 111890 42744 111946 42800
rect 113178 42744 113234 42800
rect 114190 42744 114246 42800
rect 115754 42744 115810 42800
rect 116306 42744 116362 42800
rect 118238 42744 118294 42800
rect 119066 42744 119122 42800
rect 109314 42200 109370 42256
rect 111154 42200 111210 42256
rect 133418 42744 133474 42800
rect 135902 42744 135958 42800
rect 155958 42764 156014 42800
rect 155958 42744 155960 42764
rect 155960 42744 156012 42764
rect 156012 42744 156014 42764
rect 183466 42764 183522 42800
rect 183466 42744 183468 42764
rect 183468 42744 183520 42764
rect 183520 42744 183522 42764
rect 198646 375264 198702 375320
rect 198186 264560 198242 264616
rect 200210 491952 200266 492008
rect 200210 491680 200266 491736
rect 200670 492088 200726 492144
rect 200854 492224 200910 492280
rect 199014 454688 199070 454744
rect 199198 394576 199254 394632
rect 199382 391312 199438 391368
rect 199566 461352 199622 461408
rect 199750 394576 199806 394632
rect 199566 392672 199622 392728
rect 199474 389816 199530 389872
rect 199474 389136 199530 389192
rect 199382 366288 199438 366344
rect 198830 344120 198886 344176
rect 198738 284280 198794 284336
rect 198922 280064 198978 280120
rect 198830 233960 198886 234016
rect 198738 174936 198794 174992
rect 199290 282648 199346 282704
rect 199106 281288 199162 281344
rect 199014 278568 199070 278624
rect 198830 169768 198886 169824
rect 198738 168408 198794 168464
rect 199198 233960 199254 234016
rect 199106 171264 199162 171320
rect 199014 168408 199070 168464
rect 199658 389136 199714 389192
rect 200578 374584 200634 374640
rect 199474 281288 199530 281344
rect 199842 284280 199898 284336
rect 199750 282648 199806 282704
rect 199658 280064 199714 280120
rect 199382 174936 199438 174992
rect 199290 172624 199346 172680
rect 199198 124072 199254 124128
rect 201774 492260 201776 492280
rect 201776 492260 201828 492280
rect 201828 492260 201830 492280
rect 201774 492224 201830 492260
rect 203062 373224 203118 373280
rect 202326 264424 202382 264480
rect 205730 492088 205786 492144
rect 204902 465840 204958 465896
rect 205270 262656 205326 262712
rect 206466 459040 206522 459096
rect 207662 465976 207718 466032
rect 208122 373360 208178 373416
rect 207662 152768 207718 152824
rect 209226 463256 209282 463312
rect 209686 372544 209742 372600
rect 209502 372000 209558 372056
rect 209594 371184 209650 371240
rect 199382 64640 199438 64696
rect 199290 63280 199346 63336
rect 199106 61920 199162 61976
rect 198830 60424 198886 60480
rect 198738 59200 198794 59256
rect 183190 42644 183192 42664
rect 183192 42644 183244 42664
rect 183244 42644 183246 42664
rect 183190 42608 183246 42644
rect 165802 42472 165858 42528
rect 211158 491544 211214 491600
rect 211066 369144 211122 369200
rect 210882 130464 210938 130520
rect 211618 372136 211674 372192
rect 211434 264288 211490 264344
rect 211710 370504 211766 370560
rect 212814 492496 212870 492552
rect 212814 373632 212870 373688
rect 212446 369144 212502 369200
rect 165802 39888 165858 39944
rect 212998 373632 213054 373688
rect 213090 373224 213146 373280
rect 213458 459448 213514 459504
rect 213274 263200 213330 263256
rect 213826 373768 213882 373824
rect 213458 263336 213514 263392
rect 213734 369144 213790 369200
rect 213918 372408 213974 372464
rect 213918 371728 213974 371784
rect 214286 372408 214342 372464
rect 215114 369144 215170 369200
rect 214378 131008 214434 131064
rect 214838 130464 214894 130520
rect 217230 492360 217286 492416
rect 217782 492496 217838 492552
rect 215758 262928 215814 262984
rect 216770 410896 216826 410952
rect 216770 408720 216826 408776
rect 216678 384956 216680 384976
rect 216680 384956 216732 384976
rect 216732 384956 216734 384976
rect 216678 384920 216734 384956
rect 216678 383288 216734 383344
rect 216310 372272 216366 372328
rect 215850 130328 215906 130384
rect 217230 407768 217286 407824
rect 216862 404948 216864 404968
rect 216864 404948 216916 404968
rect 216916 404948 216918 404968
rect 216862 404912 216918 404948
rect 217046 383016 217102 383072
rect 217046 375264 217102 375320
rect 217046 374992 217102 375048
rect 217322 404232 217378 404288
rect 216862 373904 216918 373960
rect 216678 372680 216734 372736
rect 216586 369824 216642 369880
rect 216494 262928 216550 262984
rect 216678 298016 216734 298072
rect 216954 295976 217010 296032
rect 216954 295296 217010 295352
rect 216862 294888 216918 294944
rect 216862 293936 216918 293992
rect 217138 301824 217194 301880
rect 217046 293120 217102 293176
rect 216678 274896 216734 274952
rect 216678 273264 216734 273320
rect 216678 272992 216734 273048
rect 216770 193160 216826 193216
rect 216770 191800 216826 191856
rect 216678 187720 216734 187776
rect 216678 165008 216734 165064
rect 216678 163376 216734 163432
rect 216862 191664 216918 191720
rect 216770 81912 216826 81968
rect 216954 185000 217010 185056
rect 216862 80960 216918 81016
rect 217874 411848 217930 411904
rect 217690 410896 217746 410952
rect 217598 406000 217654 406056
rect 217690 300872 217746 300928
rect 217322 298016 217378 298072
rect 217506 295296 217562 295352
rect 217414 293936 217470 293992
rect 217138 193160 217194 193216
rect 217046 163104 217102 163160
rect 216954 74976 217010 75032
rect 216678 53216 216734 53272
rect 217506 185952 217562 186008
rect 217414 185000 217470 185056
rect 217414 183232 217470 183288
rect 217966 407768 218022 407824
rect 217966 404232 218022 404288
rect 217966 403144 218022 403200
rect 217966 375264 218022 375320
rect 217874 301824 217930 301880
rect 217782 298696 217838 298752
rect 217690 191664 217746 191720
rect 217690 190984 217746 191040
rect 217874 293120 217930 293176
rect 217782 188672 217838 188728
rect 217506 76064 217562 76120
rect 217414 73208 217470 73264
rect 218150 372816 218206 372872
rect 218702 465704 218758 465760
rect 218518 371048 218574 371104
rect 218334 350376 218390 350432
rect 218610 369008 218666 369064
rect 218426 263608 218482 263664
rect 217966 187720 218022 187776
rect 217874 183232 217930 183288
rect 217782 78784 217838 78840
rect 218242 153040 218298 153096
rect 217966 77832 218022 77888
rect 219438 374040 219494 374096
rect 219346 372816 219402 372872
rect 219530 372136 219586 372192
rect 219622 369008 219678 369064
rect 218978 44784 219034 44840
rect 219254 44784 219310 44840
rect 224406 492496 224462 492552
rect 224866 491816 224922 491872
rect 223578 475360 223634 475416
rect 226430 467200 226486 467256
rect 229190 483656 229246 483712
rect 232318 491952 232374 492008
rect 233238 492088 233294 492144
rect 231950 479440 232006 479496
rect 231858 478080 231914 478136
rect 234158 491816 234214 491872
rect 235906 492496 235962 492552
rect 235814 492360 235870 492416
rect 235262 492224 235318 492280
rect 236550 487736 236606 487792
rect 233330 472504 233386 472560
rect 233238 467064 233294 467120
rect 221002 459584 221058 459640
rect 258170 462848 258226 462904
rect 265070 465704 265126 465760
rect 278962 474000 279018 474056
rect 278870 471144 278926 471200
rect 292578 476720 292634 476776
rect 296718 462984 296774 463040
rect 316682 582664 316738 582720
rect 317602 645224 317658 645280
rect 317694 640464 317750 640520
rect 317970 635704 318026 635760
rect 317418 630944 317474 631000
rect 317970 626184 318026 626240
rect 317970 621424 318026 621480
rect 317418 616664 317474 616720
rect 317970 611904 318026 611960
rect 317970 602384 318026 602440
rect 317970 597624 318026 597680
rect 317970 592864 318026 592920
rect 317418 586508 317420 586528
rect 317420 586508 317472 586528
rect 317472 586508 317474 586528
rect 317418 586472 317474 586508
rect 317510 577904 317566 577960
rect 317970 573144 318026 573200
rect 317970 568384 318026 568440
rect 317970 563624 318026 563680
rect 319534 647536 319590 647592
rect 318798 607144 318854 607200
rect 317970 558864 318026 558920
rect 317970 554104 318026 554160
rect 317418 549344 317474 549400
rect 317970 544584 318026 544640
rect 318338 556280 318394 556336
rect 318522 554784 318578 554840
rect 318706 539824 318762 539880
rect 328090 646176 328146 646232
rect 346582 646040 346638 646096
rect 391938 647536 391994 647592
rect 418802 647400 418858 647456
rect 405370 645904 405426 645960
rect 429198 598304 429254 598360
rect 428370 573280 428426 573336
rect 319902 556144 319958 556200
rect 319902 535336 319958 535392
rect 319718 532616 319774 532672
rect 324870 533976 324926 534032
rect 337658 532616 337714 532672
rect 339682 461216 339738 461272
rect 338302 460980 338304 461000
rect 338304 460980 338356 461000
rect 338356 460980 338358 461000
rect 338302 460944 338358 460980
rect 350998 460964 351054 461000
rect 350998 460944 351000 460964
rect 351000 460944 351052 460964
rect 351052 460944 351054 460964
rect 298098 460128 298154 460184
rect 263690 374992 263746 375048
rect 311806 374992 311862 375048
rect 244278 374468 244334 374504
rect 244278 374448 244280 374468
rect 244280 374448 244332 374468
rect 244332 374448 244334 374468
rect 248694 374448 248750 374504
rect 250074 374448 250130 374504
rect 220726 371048 220782 371104
rect 220910 371456 220966 371512
rect 236458 373632 236514 373688
rect 222106 372000 222162 372056
rect 238114 372544 238170 372600
rect 239126 372544 239182 372600
rect 222106 371456 222162 371512
rect 271142 374448 271198 374504
rect 275834 374448 275890 374504
rect 258078 373904 258134 373960
rect 242898 373632 242954 373688
rect 253938 373244 253994 373280
rect 253938 373224 253940 373244
rect 253940 373224 253992 373244
rect 253992 373224 253994 373244
rect 255410 373224 255466 373280
rect 256698 373224 256754 373280
rect 247130 373088 247186 373144
rect 244278 372544 244334 372600
rect 245658 371864 245714 371920
rect 246026 371864 246082 371920
rect 269210 373360 269266 373416
rect 261298 373088 261354 373144
rect 264978 373088 265034 373144
rect 251178 372544 251234 372600
rect 252558 372544 252614 372600
rect 259458 372544 259514 372600
rect 259642 372544 259698 372600
rect 262218 372580 262220 372600
rect 262220 372580 262272 372600
rect 262272 372580 262274 372600
rect 262218 372544 262274 372580
rect 266358 372544 266414 372600
rect 246026 371592 246082 371648
rect 251178 371628 251180 371648
rect 251180 371628 251232 371648
rect 251232 371628 251234 371648
rect 251178 371592 251234 371628
rect 258170 371592 258226 371648
rect 247038 371456 247094 371512
rect 249798 371456 249854 371512
rect 252650 371456 252706 371512
rect 255318 371456 255374 371512
rect 222014 371320 222070 371376
rect 260838 371456 260894 371512
rect 263598 371456 263654 371512
rect 264978 371456 265034 371512
rect 267738 371456 267794 371512
rect 271878 372544 271934 372600
rect 273258 372564 273314 372600
rect 314566 374720 314622 374776
rect 320914 374448 320970 374504
rect 300858 373088 300914 373144
rect 273258 372544 273260 372564
rect 273260 372544 273312 372564
rect 273312 372544 273314 372564
rect 280066 372408 280122 372464
rect 276018 371728 276074 371784
rect 270314 371320 270370 371376
rect 270498 371320 270554 371376
rect 273258 371320 273314 371376
rect 292578 372136 292634 372192
rect 277306 371456 277362 371512
rect 276018 371320 276074 371376
rect 277398 371320 277454 371376
rect 280158 371320 280214 371376
rect 282918 371320 282974 371376
rect 285678 371320 285734 371376
rect 287242 371320 287298 371376
rect 289818 371320 289874 371376
rect 295338 371320 295394 371376
rect 298098 371320 298154 371376
rect 326066 372564 326122 372600
rect 326066 372544 326068 372564
rect 326068 372544 326120 372564
rect 326120 372544 326122 372564
rect 343178 372136 343234 372192
rect 343454 372136 343510 372192
rect 302238 371728 302294 371784
rect 304998 371320 305054 371376
rect 307758 371320 307814 371376
rect 310518 371320 310574 371376
rect 313278 371320 313334 371376
rect 322938 371320 322994 371376
rect 338486 350512 338542 350568
rect 340510 350512 340566 350568
rect 351642 350512 351698 350568
rect 250442 264968 250498 265024
rect 274178 264968 274234 265024
rect 220082 240216 220138 240272
rect 291842 264560 291898 264616
rect 293406 264560 293462 264616
rect 280802 264288 280858 264344
rect 283378 264288 283434 264344
rect 285954 264288 286010 264344
rect 288162 264308 288218 264344
rect 288162 264288 288164 264308
rect 288164 264288 288216 264308
rect 288216 264288 288218 264308
rect 290922 264324 290924 264344
rect 290924 264324 290976 264344
rect 290976 264324 290978 264344
rect 290922 264288 290978 264324
rect 291842 264288 291898 264344
rect 235998 263472 236054 263528
rect 238758 263472 238814 263528
rect 243082 263472 243138 263528
rect 247130 263472 247186 263528
rect 247682 263472 247738 263528
rect 253570 263472 253626 263528
rect 256146 263472 256202 263528
rect 258170 263472 258226 263528
rect 260838 263472 260894 263528
rect 262218 263472 262274 263528
rect 263598 263472 263654 263528
rect 264978 263472 265034 263528
rect 265898 263472 265954 263528
rect 268290 263472 268346 263528
rect 269762 263472 269818 263528
rect 270866 263472 270922 263528
rect 271234 263472 271290 263528
rect 272062 263472 272118 263528
rect 273258 263472 273314 263528
rect 275926 263472 275982 263528
rect 276110 263472 276166 263528
rect 279238 263472 279294 263528
rect 305826 263492 305882 263528
rect 305826 263472 305828 263492
rect 305828 263472 305880 263492
rect 305880 263472 305882 263492
rect 237378 262248 237434 262304
rect 240138 262248 240194 262304
rect 241518 262248 241574 262304
rect 244370 262928 244426 262984
rect 244278 262248 244334 262304
rect 245658 262248 245714 262304
rect 251178 262384 251234 262440
rect 248418 262248 248474 262304
rect 249798 262248 249854 262304
rect 251270 262248 251326 262304
rect 252650 262248 252706 262304
rect 253938 262248 253994 262304
rect 255318 262248 255374 262304
rect 256698 262248 256754 262304
rect 258354 262928 258410 262984
rect 259550 262384 259606 262440
rect 259458 262248 259514 262304
rect 260930 262928 260986 262984
rect 263598 262248 263654 262304
rect 266358 262384 266414 262440
rect 266450 262248 266506 262304
rect 267738 262248 267794 262304
rect 273350 262964 273352 262984
rect 273352 262964 273404 262984
rect 273404 262964 273406 262984
rect 273350 262928 273406 262964
rect 308402 263508 308404 263528
rect 308404 263508 308456 263528
rect 308456 263508 308458 263528
rect 308402 263472 308458 263508
rect 323030 263472 323086 263528
rect 325790 263472 325846 263528
rect 343454 263472 343510 263528
rect 277306 262248 277362 262304
rect 278686 262248 278742 262304
rect 343546 263064 343602 263120
rect 339406 240216 339462 240272
rect 340050 240216 340106 240272
rect 351550 240216 351606 240272
rect 261022 154536 261078 154592
rect 273534 154536 273590 154592
rect 287978 154128 288034 154184
rect 288162 154128 288218 154184
rect 293314 154148 293370 154184
rect 293314 154128 293316 154148
rect 293316 154128 293368 154148
rect 293368 154128 293370 154148
rect 298466 154012 298522 154048
rect 298466 153992 298468 154012
rect 298468 153992 298520 154012
rect 298520 153992 298522 154012
rect 303434 153992 303490 154048
rect 287978 153856 288034 153912
rect 308402 153876 308458 153912
rect 308402 153856 308404 153876
rect 308404 153856 308456 153876
rect 308456 153856 308458 153876
rect 236090 153040 236146 153096
rect 237378 153040 237434 153096
rect 240138 153040 240194 153096
rect 241518 153040 241574 153096
rect 242898 153040 242954 153096
rect 244278 153040 244334 153096
rect 245658 153040 245714 153096
rect 247038 153040 247094 153096
rect 248418 153040 248474 153096
rect 249798 153040 249854 153096
rect 250258 153040 250314 153096
rect 251178 153040 251234 153096
rect 252558 153040 252614 153096
rect 253570 153040 253626 153096
rect 253938 153040 253994 153096
rect 255318 153040 255374 153096
rect 255962 153040 256018 153096
rect 256698 153040 256754 153096
rect 258078 153040 258134 153096
rect 259550 153040 259606 153096
rect 261206 153040 261262 153096
rect 262218 153040 262274 153096
rect 263598 153040 263654 153096
rect 264978 153040 265034 153096
rect 266358 153040 266414 153096
rect 267738 153040 267794 153096
rect 269118 153040 269174 153096
rect 270498 153040 270554 153096
rect 271878 153040 271934 153096
rect 273258 153040 273314 153096
rect 274730 153040 274786 153096
rect 277950 153040 278006 153096
rect 280066 153040 280122 153096
rect 280250 153040 280306 153096
rect 282918 153040 282974 153096
rect 285678 153076 285680 153096
rect 285680 153076 285732 153096
rect 285732 153076 285734 153096
rect 285678 153040 285734 153076
rect 289818 153060 289874 153096
rect 289818 153040 289820 153060
rect 289820 153040 289872 153060
rect 289872 153040 289874 153060
rect 235998 152360 236054 152416
rect 238758 151952 238814 152008
rect 237378 130464 237434 130520
rect 244370 152360 244426 152416
rect 247130 152380 247186 152416
rect 247130 152360 247132 152380
rect 247132 152360 247184 152380
rect 247184 152360 247186 152380
rect 249798 130872 249854 130928
rect 251270 152360 251326 152416
rect 259458 152632 259514 152688
rect 258262 152516 258318 152552
rect 258262 152496 258264 152516
rect 258264 152496 258316 152516
rect 258316 152496 258318 152516
rect 265070 152652 265126 152688
rect 265070 152632 265072 152652
rect 265072 152632 265124 152652
rect 265124 152632 265126 152652
rect 266450 152632 266506 152688
rect 268014 152632 268070 152688
rect 274638 152632 274694 152688
rect 277398 151952 277454 152008
rect 278686 151816 278742 151872
rect 274638 131008 274694 131064
rect 300858 153040 300914 153096
rect 320178 153040 320234 153096
rect 343546 152768 343602 152824
rect 343546 152516 343602 152552
rect 343546 152496 343548 152516
rect 343548 152496 343600 152516
rect 343600 152496 343602 152516
rect 269118 130328 269174 130384
rect 338486 129784 338542 129840
rect 340602 129784 340658 129840
rect 351734 129784 351790 129840
rect 235998 44784 236054 44840
rect 237102 44784 237158 44840
rect 243082 44784 243138 44840
rect 244278 44784 244334 44840
rect 255870 44648 255926 44704
rect 256974 44648 257030 44704
rect 258078 44648 258134 44704
rect 262862 44648 262918 44704
rect 315854 44648 315910 44704
rect 259458 44512 259514 44568
rect 260654 44512 260710 44568
rect 261758 44512 261814 44568
rect 263874 44512 263930 44568
rect 308494 44512 308550 44568
rect 300858 44104 300914 44160
rect 279238 43832 279294 43888
rect 265162 43152 265218 43208
rect 272154 43152 272210 43208
rect 325882 43152 325938 43208
rect 238114 42744 238170 42800
rect 239126 42744 239182 42800
rect 240506 42744 240562 42800
rect 241610 42744 241666 42800
rect 245290 42744 245346 42800
rect 246394 42744 246450 42800
rect 250074 42744 250130 42800
rect 251178 42744 251234 42800
rect 253386 42744 253442 42800
rect 260930 42744 260986 42800
rect 248602 41928 248658 41984
rect 247682 41792 247738 41848
rect 251730 41928 251786 41984
rect 250074 39888 250130 39944
rect 254122 42064 254178 42120
rect 268198 42744 268254 42800
rect 268474 42744 268530 42800
rect 271234 42744 271290 42800
rect 266358 42336 266414 42392
rect 266634 42336 266690 42392
rect 269762 42336 269818 42392
rect 273258 42744 273314 42800
rect 276110 42744 276166 42800
rect 276938 42744 276994 42800
rect 278318 42744 278374 42800
rect 293314 42744 293370 42800
rect 298466 42744 298522 42800
rect 302514 42744 302570 42800
rect 310978 42744 311034 42800
rect 313370 42744 313426 42800
rect 318338 42744 318394 42800
rect 320914 42764 320970 42800
rect 320914 42744 320916 42764
rect 320916 42744 320968 42764
rect 320968 42744 320970 42764
rect 273534 42200 273590 42256
rect 274730 42200 274786 42256
rect 343178 42764 343234 42800
rect 343178 42744 343180 42764
rect 343180 42744 343232 42764
rect 343232 42744 343234 42764
rect 343454 42744 343510 42800
rect 358818 454688 358874 454744
rect 358910 393760 358966 393816
rect 359002 390768 359058 390824
rect 359094 388048 359150 388104
rect 359094 366288 359150 366344
rect 358910 344120 358966 344176
rect 358818 284280 358874 284336
rect 359186 282376 359242 282432
rect 359002 280064 359058 280120
rect 359094 278704 359150 278760
rect 358910 233960 358966 234016
rect 358818 174936 358874 174992
rect 358818 172352 358874 172408
rect 358818 171264 358874 171320
rect 358542 151680 358598 151736
rect 359922 392128 359978 392184
rect 359830 389272 359886 389328
rect 359370 280064 359426 280120
rect 359278 233960 359334 234016
rect 359186 172624 359242 172680
rect 358910 169768 358966 169824
rect 358818 61920 358874 61976
rect 359002 168544 359058 168600
rect 358910 60424 358966 60480
rect 359646 284280 359702 284336
rect 359554 281424 359610 281480
rect 359462 278704 359518 278760
rect 359370 169768 359426 169824
rect 359554 174936 359610 174992
rect 359278 124072 359334 124128
rect 359646 172352 359702 172408
rect 359554 64640 359610 64696
rect 359186 63280 359242 63336
rect 359002 59200 359058 59256
rect 361210 151544 361266 151600
rect 362222 44376 362278 44432
rect 366730 262656 366786 262712
rect 368386 372000 368442 372056
rect 367926 152224 367982 152280
rect 370594 152904 370650 152960
rect 372434 371864 372490 371920
rect 372986 369008 373042 369064
rect 373446 263336 373502 263392
rect 374366 133728 374422 133784
rect 375194 373904 375250 373960
rect 375286 372680 375342 372736
rect 375838 239808 375894 239864
rect 377034 407768 377090 407824
rect 376942 384956 376944 384976
rect 376944 384956 376996 384976
rect 376996 384956 376998 384976
rect 376942 384920 376998 384956
rect 376942 383288 376998 383344
rect 376850 383016 376906 383072
rect 376390 263064 376446 263120
rect 376022 53080 376078 53136
rect 377126 370368 377182 370424
rect 377310 409944 377366 410000
rect 377402 407768 377458 407824
rect 377402 406000 377458 406056
rect 377586 411848 377642 411904
rect 377218 301824 377274 301880
rect 376850 300872 376906 300928
rect 376758 295296 376814 295352
rect 376942 298696 376998 298752
rect 377126 293936 377182 293992
rect 376850 274896 376906 274952
rect 376758 273264 376814 273320
rect 376758 272992 376814 273048
rect 376850 191664 376906 191720
rect 376942 188672 376998 188728
rect 376942 187856 376998 187912
rect 376942 185952 376998 186008
rect 376758 163104 376814 163160
rect 376942 165008 376998 165064
rect 376942 163376 376998 163432
rect 376574 130328 376630 130384
rect 377402 300872 377458 300928
rect 377310 297744 377366 297800
rect 377218 193160 377274 193216
rect 377218 187856 377274 187912
rect 377126 185000 377182 185056
rect 376942 76064 376998 76120
rect 377770 410896 377826 410952
rect 377770 409944 377826 410000
rect 377862 408720 377918 408776
rect 377678 404948 377680 404968
rect 377680 404948 377732 404968
rect 377732 404948 377734 404968
rect 377678 404912 377734 404948
rect 377586 301824 377642 301880
rect 377770 403144 377826 403200
rect 377678 294888 377734 294944
rect 377678 293936 377734 293992
rect 377954 406000 378010 406056
rect 377862 298696 377918 298752
rect 378046 372680 378102 372736
rect 377954 295976 378010 296032
rect 377954 295296 378010 295352
rect 377770 293120 377826 293176
rect 377310 187720 377366 187776
rect 377494 183504 377550 183560
rect 377218 129784 377274 129840
rect 377126 74976 377182 75032
rect 376942 54984 376998 55040
rect 376942 53216 376998 53272
rect 377310 78784 377366 78840
rect 378506 262928 378562 262984
rect 378046 239808 378102 239864
rect 377954 193160 378010 193216
rect 377954 191800 378010 191856
rect 377862 191664 377918 191720
rect 377862 190848 377918 190904
rect 377770 183504 377826 183560
rect 377678 133728 377734 133784
rect 377494 73208 377550 73264
rect 378046 187720 378102 187776
rect 377954 81912 378010 81968
rect 377862 80960 377918 81016
rect 378046 77832 378102 77888
rect 378966 152768 379022 152824
rect 379242 263200 379298 263256
rect 379150 152632 379206 152688
rect 379610 369824 379666 369880
rect 379518 260616 379574 260672
rect 428462 563760 428518 563816
rect 428554 535880 428610 535936
rect 430578 641144 430634 641200
rect 430854 647264 430910 647320
rect 430762 636384 430818 636440
rect 430670 631624 430726 631680
rect 430854 626864 430910 626920
rect 430578 617344 430634 617400
rect 429382 593544 429438 593600
rect 429290 545264 429346 545320
rect 429474 588104 429530 588160
rect 430670 612584 430726 612640
rect 430762 603064 430818 603120
rect 430854 583344 430910 583400
rect 430578 540504 430634 540560
rect 430946 578584 431002 578640
rect 431038 569064 431094 569120
rect 431130 559544 431186 559600
rect 431222 554784 431278 554840
rect 431314 550024 431370 550080
rect 580262 671880 580318 671936
rect 580262 670656 580318 670712
rect 580906 670656 580962 670712
rect 579894 659096 579950 659152
rect 456798 634616 456854 634672
rect 456798 626320 456854 626376
rect 510618 623056 510674 623112
rect 457442 618160 457498 618216
rect 457442 608912 457498 608968
rect 436742 533976 436798 534032
rect 457534 600752 457590 600808
rect 511262 597624 511318 597680
rect 457626 592592 457682 592648
rect 511998 630536 512054 630592
rect 511998 614080 512054 614136
rect 580906 620744 580962 620800
rect 580262 607960 580318 608016
rect 512090 605920 512146 605976
rect 512182 589328 512238 589384
rect 580906 569472 580962 569528
rect 580170 556688 580226 556744
rect 511262 462168 511318 462224
rect 498474 460980 498476 461000
rect 498476 460980 498528 461000
rect 498528 460980 498530 461000
rect 498474 460944 498530 460980
rect 499854 460944 499910 461000
rect 516598 454688 516654 454744
rect 407762 374992 407818 375048
rect 418250 374992 418306 375048
rect 440330 374992 440386 375048
rect 443090 374992 443146 375048
rect 410706 374584 410762 374640
rect 433338 374468 433394 374504
rect 433338 374448 433340 374468
rect 433340 374448 433392 374468
rect 433392 374448 433394 374468
rect 433614 374448 433670 374504
rect 445942 374448 445998 374504
rect 448242 374448 448298 374504
rect 415674 374176 415730 374232
rect 434810 374176 434866 374232
rect 404818 373768 404874 373824
rect 405738 372136 405794 372192
rect 396078 372020 396134 372056
rect 396078 372000 396080 372020
rect 396080 372000 396132 372020
rect 396132 372000 396134 372020
rect 398838 372000 398894 372056
rect 397458 371864 397514 371920
rect 412822 371864 412878 371920
rect 409878 371748 409934 371784
rect 409878 371728 409880 371748
rect 409880 371728 409932 371748
rect 409932 371728 409934 371748
rect 411258 371728 411314 371784
rect 407118 371612 407174 371648
rect 407118 371592 407120 371612
rect 407120 371592 407172 371612
rect 407172 371592 407174 371612
rect 412638 371592 412694 371648
rect 411258 371476 411314 371512
rect 411258 371456 411260 371476
rect 411260 371456 411312 371476
rect 411312 371456 411314 371476
rect 396078 371320 396134 371376
rect 402978 371320 403034 371376
rect 403254 371320 403310 371376
rect 408498 371320 408554 371376
rect 414018 371320 414074 371376
rect 415398 371320 415454 371376
rect 421010 373768 421066 373824
rect 423034 373804 423036 373824
rect 423036 373804 423088 373824
rect 423088 373804 423090 373824
rect 423034 373768 423090 373804
rect 425426 373768 425482 373824
rect 439410 373788 439466 373824
rect 439410 373768 439412 373788
rect 439412 373768 439464 373788
rect 439464 373768 439466 373788
rect 460938 373768 460994 373824
rect 438214 373088 438270 373144
rect 425058 372580 425060 372600
rect 425060 372580 425112 372600
rect 425112 372580 425114 372600
rect 425058 372544 425114 372580
rect 426438 372544 426494 372600
rect 427818 372544 427874 372600
rect 450266 373652 450322 373688
rect 450266 373632 450268 373652
rect 450268 373632 450320 373652
rect 450320 373632 450322 373652
rect 452842 373516 452898 373552
rect 452842 373496 452844 373516
rect 452844 373496 452896 373516
rect 452896 373496 452898 373516
rect 458178 373496 458234 373552
rect 462778 373496 462834 373552
rect 455418 373380 455474 373416
rect 455418 373360 455420 373380
rect 455420 373360 455472 373380
rect 455472 373360 455474 373380
rect 430578 371728 430634 371784
rect 418250 371456 418306 371512
rect 422298 371456 422354 371512
rect 426438 371456 426494 371512
rect 416778 371320 416834 371376
rect 418158 371320 418214 371376
rect 419538 371320 419594 371376
rect 420918 371320 420974 371376
rect 423678 371320 423734 371376
rect 420918 369008 420974 369064
rect 427818 371320 427874 371376
rect 429198 371320 429254 371376
rect 470598 372272 470654 372328
rect 465078 371592 465134 371648
rect 430670 371320 430726 371376
rect 431958 371320 432014 371376
rect 436098 371320 436154 371376
rect 437478 371320 437534 371376
rect 467838 371320 467894 371376
rect 503166 372136 503222 372192
rect 483018 371864 483074 371920
rect 473358 371320 473414 371376
rect 480258 371320 480314 371376
rect 485778 371320 485834 371376
rect 502338 371320 502394 371376
rect 499026 350512 499082 350568
rect 500590 350512 500646 350568
rect 510894 350548 510896 350568
rect 510896 350548 510948 350568
rect 510948 350548 510950 350568
rect 510894 350512 510950 350548
rect 380990 349696 381046 349752
rect 473450 264832 473506 264888
rect 480902 264832 480958 264888
rect 468482 264696 468538 264752
rect 470966 264696 471022 264752
rect 418434 264560 418490 264616
rect 421102 264560 421158 264616
rect 423494 264560 423550 264616
rect 425978 264560 426034 264616
rect 429750 264560 429806 264616
rect 475842 264560 475898 264616
rect 483386 264696 483442 264752
rect 485962 264696 486018 264752
rect 415858 263608 415914 263664
rect 397458 263472 397514 263528
rect 401598 263472 401654 263528
rect 404358 263472 404414 263528
rect 408314 263472 408370 263528
rect 410706 263472 410762 263528
rect 413650 263472 413706 263528
rect 415766 263472 415822 263528
rect 396078 262792 396134 262848
rect 379886 240216 379942 240272
rect 379702 239536 379758 239592
rect 379610 131008 379666 131064
rect 380346 260888 380402 260944
rect 393962 260072 394018 260128
rect 393962 240760 394018 240816
rect 396170 262248 396226 262304
rect 398838 262248 398894 262304
rect 400218 262248 400274 262304
rect 403070 262384 403126 262440
rect 402978 262248 403034 262304
rect 412730 262792 412786 262848
rect 411258 262384 411314 262440
rect 405738 262248 405794 262304
rect 407210 262248 407266 262304
rect 408498 262248 408554 262304
rect 409878 262248 409934 262304
rect 411350 262248 411406 262304
rect 414018 262248 414074 262304
rect 419354 263472 419410 263528
rect 425242 263472 425298 263528
rect 426438 263472 426494 263528
rect 427450 263472 427506 263528
rect 428186 263472 428242 263528
rect 430946 263472 431002 263528
rect 432234 263472 432290 263528
rect 433338 263472 433394 263528
rect 434626 263472 434682 263528
rect 418158 262792 418214 262848
rect 416778 262248 416834 262304
rect 419814 262928 419870 262984
rect 421746 262928 421802 262984
rect 423954 262520 424010 262576
rect 423586 262248 423642 262304
rect 416778 240760 416834 240816
rect 428278 262268 428334 262304
rect 428278 262248 428280 262268
rect 428280 262248 428332 262268
rect 428332 262248 428334 262268
rect 430670 262248 430726 262304
rect 393962 239400 394018 239456
rect 433522 262964 433524 262984
rect 433524 262964 433576 262984
rect 433576 262964 433578 262984
rect 433522 262928 433578 262964
rect 435914 263472 435970 263528
rect 438766 263472 438822 263528
rect 440882 263472 440938 263528
rect 443458 263472 443514 263528
rect 448242 263472 448298 263528
rect 451002 263472 451058 263528
rect 453394 263508 453396 263528
rect 453396 263508 453448 263528
rect 453448 263508 453450 263528
rect 453394 263472 453450 263508
rect 455786 263492 455842 263528
rect 455786 263472 455788 263492
rect 455788 263472 455840 263492
rect 455840 263472 455842 263492
rect 435178 262928 435234 262984
rect 438398 262928 438454 262984
rect 436098 262248 436154 262304
rect 503534 263472 503590 263528
rect 440146 262248 440202 262304
rect 503626 262248 503682 262304
rect 511906 241440 511962 241496
rect 499026 240216 499082 240272
rect 500774 240216 500830 240272
rect 418434 154400 418490 154456
rect 421010 154436 421012 154456
rect 421012 154436 421064 154456
rect 421064 154436 421066 154456
rect 421010 154400 421066 154436
rect 425978 154420 426034 154456
rect 425978 154400 425980 154420
rect 425980 154400 426032 154420
rect 426032 154400 426034 154420
rect 443458 154400 443514 154456
rect 423402 153856 423458 153912
rect 475842 154284 475898 154320
rect 475842 154264 475844 154284
rect 475844 154264 475896 154284
rect 475896 154264 475898 154284
rect 478418 154264 478474 154320
rect 473450 154148 473506 154184
rect 473450 154128 473452 154148
rect 473452 154128 473504 154148
rect 473504 154128 473506 154148
rect 480810 154128 480866 154184
rect 470874 154012 470930 154048
rect 470874 153992 470876 154012
rect 470876 153992 470928 154012
rect 470928 153992 470930 154012
rect 483202 153992 483258 154048
rect 485962 153876 486018 153912
rect 485962 153856 485964 153876
rect 485964 153856 486016 153876
rect 486016 153856 486018 153876
rect 396078 153040 396134 153096
rect 397458 153040 397514 153096
rect 398838 153040 398894 153096
rect 400218 153040 400274 153096
rect 401598 153040 401654 153096
rect 403070 153040 403126 153096
rect 404358 153040 404414 153096
rect 405738 153040 405794 153096
rect 407210 153040 407266 153096
rect 408498 153040 408554 153096
rect 409970 153040 410026 153096
rect 411350 153040 411406 153096
rect 412730 153040 412786 153096
rect 414018 153040 414074 153096
rect 415490 153040 415546 153096
rect 415674 153040 415730 153096
rect 416778 153040 416834 153096
rect 418250 153040 418306 153096
rect 419538 153040 419594 153096
rect 420918 153040 420974 153096
rect 422298 153040 422354 153096
rect 423678 153040 423734 153096
rect 425058 153040 425114 153096
rect 426530 153040 426586 153096
rect 427818 153040 427874 153096
rect 429198 153040 429254 153096
rect 430578 153040 430634 153096
rect 431958 153040 432014 153096
rect 433338 153040 433394 153096
rect 433982 153040 434038 153096
rect 434810 153040 434866 153096
rect 436190 153040 436246 153096
rect 438858 153040 438914 153096
rect 440146 153040 440202 153096
rect 440330 153040 440386 153096
rect 445758 153040 445814 153096
rect 447138 153076 447140 153096
rect 447140 153076 447192 153096
rect 447192 153076 447194 153096
rect 447138 153040 447194 153076
rect 449898 153040 449954 153096
rect 452658 153040 452714 153096
rect 455418 153040 455474 153096
rect 458178 153060 458234 153096
rect 458178 153040 458180 153060
rect 458180 153040 458232 153060
rect 458232 153040 458234 153060
rect 380806 151272 380862 151328
rect 396170 152496 396226 152552
rect 379886 130736 379942 130792
rect 402978 152496 403034 152552
rect 407118 152360 407174 152416
rect 409878 152496 409934 152552
rect 411258 152496 411314 152552
rect 413098 152496 413154 152552
rect 418158 152496 418214 152552
rect 426438 152496 426494 152552
rect 426438 131008 426494 131064
rect 416778 130872 416834 130928
rect 414018 130736 414074 130792
rect 434718 152496 434774 152552
rect 436098 152496 436154 152552
rect 437478 152496 437534 152552
rect 438858 133048 438914 133104
rect 503626 152652 503682 152688
rect 503626 152632 503628 152652
rect 503628 152632 503680 152652
rect 503680 152632 503682 152652
rect 503626 152516 503682 152552
rect 503626 152496 503628 152516
rect 503628 152496 503680 152516
rect 503680 152496 503682 152516
rect 429198 130328 429254 130384
rect 518898 454144 518954 454200
rect 510618 130364 510620 130384
rect 510620 130364 510672 130384
rect 510672 130364 510674 130384
rect 510618 130328 510674 130364
rect 498750 129784 498806 129840
rect 500222 129784 500278 129840
rect 396078 44784 396134 44840
rect 397090 44784 397146 44840
rect 403070 44784 403126 44840
rect 414570 44784 414626 44840
rect 416962 44784 417018 44840
rect 410706 44648 410762 44704
rect 404174 44512 404230 44568
rect 405462 44512 405518 44568
rect 406474 44512 406530 44568
rect 419446 44648 419502 44704
rect 423954 44648 424010 44704
rect 418158 44512 418214 44568
rect 420642 44512 420698 44568
rect 421746 44512 421802 44568
rect 422850 44512 422906 44568
rect 425978 44512 426034 44568
rect 439226 44512 439282 44568
rect 455878 44512 455934 44568
rect 458454 44512 458510 44568
rect 425242 44376 425298 44432
rect 407578 43424 407634 43480
rect 421010 43424 421066 43480
rect 428186 43444 428242 43480
rect 428186 43424 428188 43444
rect 428188 43424 428240 43444
rect 428240 43424 428242 43444
rect 398194 43152 398250 43208
rect 401690 43152 401746 43208
rect 399390 42744 399446 42800
rect 400310 41792 400366 41848
rect 408314 42744 408370 42800
rect 408682 42744 408738 42800
rect 409970 42744 410026 42800
rect 411258 42744 411314 42800
rect 411902 42744 411958 42800
rect 413282 42744 413338 42800
rect 413650 42744 413706 42800
rect 415490 42744 415546 42800
rect 426438 42744 426494 42800
rect 427634 42744 427690 42800
rect 428554 42744 428610 42800
rect 429658 42744 429714 42800
rect 430946 42744 431002 42800
rect 432142 42744 432198 42800
rect 433338 42744 433394 42800
rect 434626 42744 434682 42800
rect 435914 42744 435970 42800
rect 436374 42744 436430 42800
rect 438490 42744 438546 42800
rect 440882 42744 440938 42800
rect 443458 42744 443514 42800
rect 445850 42744 445906 42800
rect 448242 42744 448298 42800
rect 453394 42744 453450 42800
rect 485962 42764 486018 42800
rect 485962 42744 485964 42764
rect 485964 42744 486016 42764
rect 486016 42744 486018 42764
rect 431130 41928 431186 41984
rect 428554 40840 428610 40896
rect 433338 40976 433394 41032
rect 435178 42064 435234 42120
rect 503258 42764 503314 42800
rect 503258 42744 503260 42764
rect 503260 42744 503312 42764
rect 503312 42744 503314 42764
rect 503534 42744 503590 42800
rect 519174 393760 519230 393816
rect 518990 390768 519046 390824
rect 519082 389272 519138 389328
rect 519358 392128 519414 392184
rect 519266 388048 519322 388104
rect 518990 343712 519046 343768
rect 518898 284688 518954 284744
rect 519082 281424 519138 281480
rect 518990 234504 519046 234560
rect 518898 174256 518954 174312
rect 519174 279792 519230 279848
rect 519082 171264 519138 171320
rect 518898 64776 518954 64832
rect 519082 169768 519138 169824
rect 519358 284688 519414 284744
rect 519450 282648 519506 282704
rect 519266 278568 519322 278624
rect 518990 61920 519046 61976
rect 519358 234504 519414 234560
rect 519266 168952 519322 169008
rect 519082 60424 519138 60480
rect 519542 281424 519598 281480
rect 580906 518336 580962 518392
rect 580170 492768 580226 492824
rect 580906 467064 580962 467120
rect 579894 441532 579896 441552
rect 579896 441532 579948 441552
rect 579948 441532 579950 441552
rect 579894 441496 579950 441532
rect 580906 415928 580962 415984
rect 578882 390360 578938 390416
rect 580906 364792 580962 364848
rect 580170 339088 580226 339144
rect 580906 313520 580962 313576
rect 519634 279792 519690 279848
rect 580906 262384 580962 262440
rect 580906 223896 580962 223952
rect 580906 185544 580962 185600
rect 519450 172624 519506 172680
rect 519358 124072 519414 124128
rect 580906 147192 580962 147248
rect 580906 108704 580962 108760
rect 580906 70352 580962 70408
rect 519450 63280 519506 63336
rect 519266 59200 519322 59256
rect 580446 32000 580502 32056
rect 580906 32000 580962 32056
<< metal3 >>
rect -960 697492 480 697732
rect 583520 697356 584960 697596
rect -960 685130 480 685220
rect 3417 685130 3483 685133
rect -960 685128 3483 685130
rect -960 685072 3422 685128
rect 3478 685072 3483 685128
rect -960 685070 3483 685072
rect -960 684980 480 685070
rect 3417 685067 3483 685070
rect 583520 684572 584960 684812
rect -960 672332 480 672572
rect 580257 671938 580323 671941
rect 583520 671938 584960 672028
rect 580257 671936 584960 671938
rect 580257 671880 580262 671936
rect 580318 671880 584960 671936
rect 580257 671878 584960 671880
rect 580257 671875 580323 671878
rect 583520 671788 584960 671878
rect 580257 670714 580323 670717
rect 580901 670714 580967 670717
rect 580257 670712 580967 670714
rect 580257 670656 580262 670712
rect 580318 670656 580906 670712
rect 580962 670656 580967 670712
rect 580257 670654 580967 670656
rect 580257 670651 580323 670654
rect 580901 670651 580967 670654
rect -960 659970 480 660060
rect 2773 659970 2839 659973
rect -960 659968 2839 659970
rect -960 659912 2778 659968
rect 2834 659912 2839 659968
rect -960 659910 2839 659912
rect -960 659820 480 659910
rect 2773 659907 2839 659910
rect 579889 659154 579955 659157
rect 583520 659154 584960 659244
rect 579889 659152 584960 659154
rect 579889 659096 579894 659152
rect 579950 659096 584960 659152
rect 579889 659094 584960 659096
rect 579889 659091 579955 659094
rect 583520 659004 584960 659094
rect 319529 647594 319595 647597
rect 391933 647594 391999 647597
rect 319529 647592 391999 647594
rect 319529 647536 319534 647592
rect 319590 647536 391938 647592
rect 391994 647536 391999 647592
rect 319529 647534 391999 647536
rect 319529 647531 319595 647534
rect 391933 647531 391999 647534
rect 309777 647458 309843 647461
rect 418797 647458 418863 647461
rect 309777 647456 418863 647458
rect -960 647172 480 647412
rect 309777 647400 309782 647456
rect 309838 647400 418802 647456
rect 418858 647400 418863 647456
rect 309777 647398 418863 647400
rect 309777 647395 309843 647398
rect 418797 647395 418863 647398
rect 281073 647322 281139 647325
rect 430849 647322 430915 647325
rect 281073 647320 430915 647322
rect 281073 647264 281078 647320
rect 281134 647264 430854 647320
rect 430910 647264 430915 647320
rect 281073 647262 430915 647264
rect 281073 647259 281139 647262
rect 430849 647259 430915 647262
rect 53046 646172 53052 646236
rect 53116 646234 53122 646236
rect 328085 646234 328151 646237
rect 53116 646232 328151 646234
rect 53116 646176 328090 646232
rect 328146 646176 328151 646232
rect 583520 646220 584960 646460
rect 53116 646174 328151 646176
rect 53116 646172 53122 646174
rect 328085 646171 328151 646174
rect 51574 646036 51580 646100
rect 51644 646098 51650 646100
rect 346577 646098 346643 646101
rect 51644 646096 346643 646098
rect 51644 646040 346582 646096
rect 346638 646040 346643 646096
rect 51644 646038 346643 646040
rect 51644 646036 51650 646038
rect 346577 646035 346643 646038
rect 54334 645900 54340 645964
rect 54404 645962 54410 645964
rect 405365 645962 405431 645965
rect 54404 645960 405431 645962
rect 54404 645904 405370 645960
rect 405426 645904 405431 645960
rect 54404 645902 405431 645904
rect 54404 645900 54410 645902
rect 405365 645899 405431 645902
rect 317597 645282 317663 645285
rect 317597 645280 320068 645282
rect 317597 645224 317602 645280
rect 317658 645224 320068 645280
rect 317597 645222 320068 645224
rect 317597 645219 317663 645222
rect 430573 641202 430639 641205
rect 428812 641200 430639 641202
rect 428812 641144 430578 641200
rect 430634 641144 430639 641200
rect 428812 641142 430639 641144
rect 430573 641139 430639 641142
rect 317689 640522 317755 640525
rect 317689 640520 320068 640522
rect 317689 640464 317694 640520
rect 317750 640464 320068 640520
rect 317689 640462 320068 640464
rect 317689 640459 317755 640462
rect 430757 636442 430823 636445
rect 428812 636440 430823 636442
rect 428812 636384 430762 636440
rect 430818 636384 430823 636440
rect 428812 636382 430823 636384
rect 430757 636379 430823 636382
rect 317965 635762 318031 635765
rect 317965 635760 320068 635762
rect 317965 635704 317970 635760
rect 318026 635704 320068 635760
rect 317965 635702 320068 635704
rect 317965 635699 318031 635702
rect 57421 635626 57487 635629
rect 137277 635626 137343 635629
rect 216673 635626 216739 635629
rect 57421 635624 60076 635626
rect 57421 635568 57426 635624
rect 57482 635568 60076 635624
rect 57421 635566 60076 635568
rect 137277 635624 140116 635626
rect 137277 635568 137282 635624
rect 137338 635568 140116 635624
rect 137277 635566 140116 635568
rect 216673 635624 220156 635626
rect 216673 635568 216678 635624
rect 216734 635568 220156 635624
rect 216673 635566 220156 635568
rect 57421 635563 57487 635566
rect 137277 635563 137343 635566
rect 216673 635563 216739 635566
rect 122925 634946 122991 634949
rect 201585 634946 201651 634949
rect 281625 634946 281691 634949
rect 120796 634944 122991 634946
rect -960 634810 480 634900
rect 120796 634888 122930 634944
rect 122986 634888 122991 634944
rect 120796 634886 122991 634888
rect 200836 634944 201651 634946
rect 200836 634888 201590 634944
rect 201646 634888 201651 634944
rect 200836 634886 201651 634888
rect 280876 634944 281691 634946
rect 280876 634888 281630 634944
rect 281686 634888 281691 634944
rect 280876 634886 281691 634888
rect 122925 634883 122991 634886
rect 201585 634883 201651 634886
rect 281625 634883 281691 634886
rect 3417 634810 3483 634813
rect -960 634808 3483 634810
rect -960 634752 3422 634808
rect 3478 634752 3483 634808
rect -960 634750 3483 634752
rect -960 634660 480 634750
rect 3417 634747 3483 634750
rect 456793 634674 456859 634677
rect 456793 634672 460122 634674
rect 456793 634616 456798 634672
rect 456854 634616 460122 634672
rect 456793 634614 460122 634616
rect 456793 634611 456859 634614
rect 460062 634032 460122 634614
rect 583520 633436 584960 633676
rect 59077 632906 59143 632909
rect 139117 632906 139183 632909
rect 216673 632906 216739 632909
rect 59077 632904 60076 632906
rect 59077 632848 59082 632904
rect 59138 632848 60076 632904
rect 59077 632846 60076 632848
rect 139117 632904 140032 632906
rect 139117 632848 139122 632904
rect 139178 632848 140032 632904
rect 139117 632846 140032 632848
rect 216673 632904 220064 632906
rect 216673 632848 216678 632904
rect 216734 632848 220064 632904
rect 216673 632846 220064 632848
rect 59077 632843 59143 632846
rect 139117 632843 139183 632846
rect 216673 632843 216739 632846
rect 123017 632226 123083 632229
rect 201769 632226 201835 632229
rect 282085 632226 282151 632229
rect 120796 632224 123083 632226
rect 120796 632168 123022 632224
rect 123078 632168 123083 632224
rect 120796 632166 123083 632168
rect 200836 632224 201835 632226
rect 200836 632168 201774 632224
rect 201830 632168 201835 632224
rect 200836 632166 201835 632168
rect 280876 632224 282151 632226
rect 280876 632168 282090 632224
rect 282146 632168 282151 632224
rect 280876 632166 282151 632168
rect 123017 632163 123083 632166
rect 201769 632163 201835 632166
rect 282085 632163 282151 632166
rect 430665 631682 430731 631685
rect 428812 631680 430731 631682
rect 428812 631624 430670 631680
rect 430726 631624 430731 631680
rect 428812 631622 430731 631624
rect 430665 631619 430731 631622
rect 317413 631002 317479 631005
rect 317413 631000 320068 631002
rect 317413 630944 317418 631000
rect 317474 630944 320068 631000
rect 317413 630942 320068 630944
rect 317413 630939 317479 630942
rect 509926 630594 509986 630632
rect 511993 630594 512059 630597
rect 509926 630592 512059 630594
rect 509926 630536 511998 630592
rect 512054 630536 512059 630592
rect 509926 630534 512059 630536
rect 511993 630531 512059 630534
rect 57697 629506 57763 629509
rect 137737 629506 137803 629509
rect 217685 629506 217751 629509
rect 57697 629504 60076 629506
rect 57697 629448 57702 629504
rect 57758 629448 60076 629504
rect 57697 629446 60076 629448
rect 137737 629504 140032 629506
rect 137737 629448 137742 629504
rect 137798 629448 140032 629504
rect 137737 629446 140032 629448
rect 217685 629504 220064 629506
rect 217685 629448 217690 629504
rect 217746 629448 220064 629504
rect 217685 629446 220064 629448
rect 57697 629443 57763 629446
rect 137737 629443 137803 629446
rect 217685 629443 217751 629446
rect 122189 628826 122255 628829
rect 201677 628826 201743 628829
rect 283465 628826 283531 628829
rect 120796 628824 122255 628826
rect 120796 628768 122194 628824
rect 122250 628768 122255 628824
rect 120796 628766 122255 628768
rect 200836 628824 201743 628826
rect 200836 628768 201682 628824
rect 201738 628768 201743 628824
rect 200836 628766 201743 628768
rect 280876 628824 283531 628826
rect 280876 628768 283470 628824
rect 283526 628768 283531 628824
rect 280876 628766 283531 628768
rect 122189 628763 122255 628766
rect 201677 628763 201743 628766
rect 283465 628763 283531 628766
rect 430849 626922 430915 626925
rect 428812 626920 430915 626922
rect 428812 626864 430854 626920
rect 430910 626864 430915 626920
rect 428812 626862 430915 626864
rect 430849 626859 430915 626862
rect 57605 626786 57671 626789
rect 139025 626786 139091 626789
rect 216673 626786 216739 626789
rect 57605 626784 60076 626786
rect 57605 626728 57610 626784
rect 57666 626728 60076 626784
rect 57605 626726 60076 626728
rect 139025 626784 140032 626786
rect 139025 626728 139030 626784
rect 139086 626728 140032 626784
rect 139025 626726 140032 626728
rect 216673 626784 220064 626786
rect 216673 626728 216678 626784
rect 216734 626728 220064 626784
rect 216673 626726 220064 626728
rect 57605 626723 57671 626726
rect 139025 626723 139091 626726
rect 216673 626723 216739 626726
rect 456793 626378 456859 626381
rect 456793 626376 460122 626378
rect 456793 626320 456798 626376
rect 456854 626320 460122 626376
rect 456793 626318 460122 626320
rect 456793 626315 456859 626318
rect 317965 626242 318031 626245
rect 317965 626240 320068 626242
rect 317965 626184 317970 626240
rect 318026 626184 320068 626240
rect 317965 626182 320068 626184
rect 317965 626179 318031 626182
rect 121821 626106 121887 626109
rect 201953 626106 202019 626109
rect 281717 626106 281783 626109
rect 120796 626104 121887 626106
rect 120796 626048 121826 626104
rect 121882 626048 121887 626104
rect 120796 626046 121887 626048
rect 200836 626104 202019 626106
rect 200836 626048 201958 626104
rect 202014 626048 202019 626104
rect 200836 626046 202019 626048
rect 280876 626104 281783 626106
rect 280876 626048 281722 626104
rect 281778 626048 281783 626104
rect 280876 626046 281783 626048
rect 121821 626043 121887 626046
rect 201953 626043 202019 626046
rect 281717 626043 281783 626046
rect 460062 625872 460122 626318
rect 58893 623386 58959 623389
rect 136633 623386 136699 623389
rect 216673 623386 216739 623389
rect 58893 623384 60076 623386
rect 58893 623328 58898 623384
rect 58954 623328 60076 623384
rect 58893 623326 60076 623328
rect 136633 623384 140032 623386
rect 136633 623328 136638 623384
rect 136694 623328 140032 623384
rect 136633 623326 140032 623328
rect 216673 623384 220064 623386
rect 216673 623328 216678 623384
rect 216734 623328 220064 623384
rect 216673 623326 220064 623328
rect 58893 623323 58959 623326
rect 136633 623323 136699 623326
rect 216673 623323 216739 623326
rect 510613 623114 510679 623117
rect 509926 623112 510679 623114
rect 509926 623056 510618 623112
rect 510674 623056 510679 623112
rect 509926 623054 510679 623056
rect 121729 622706 121795 622709
rect 202965 622706 203031 622709
rect 283005 622706 283071 622709
rect 120796 622704 121795 622706
rect 120796 622648 121734 622704
rect 121790 622648 121795 622704
rect 120796 622646 121795 622648
rect 200836 622704 203031 622706
rect 200836 622648 202970 622704
rect 203026 622648 203031 622704
rect 200836 622646 203031 622648
rect 280876 622704 283071 622706
rect 280876 622648 283010 622704
rect 283066 622648 283071 622704
rect 280876 622646 283071 622648
rect 121729 622643 121795 622646
rect 202965 622643 203031 622646
rect 283005 622643 283071 622646
rect 509926 622472 509986 623054
rect 510613 623051 510679 623054
rect -960 622148 480 622388
rect 430614 622162 430620 622164
rect 428812 622102 430620 622162
rect 430614 622100 430620 622102
rect 430684 622100 430690 622164
rect 317965 621482 318031 621485
rect 317965 621480 320068 621482
rect 317965 621424 317970 621480
rect 318026 621424 320068 621480
rect 317965 621422 320068 621424
rect 317965 621419 318031 621422
rect 580901 620802 580967 620805
rect 583520 620802 584960 620892
rect 580901 620800 584960 620802
rect 580901 620744 580906 620800
rect 580962 620744 584960 620800
rect 580901 620742 584960 620744
rect 580901 620739 580967 620742
rect 58985 620666 59051 620669
rect 137093 620666 137159 620669
rect 219249 620666 219315 620669
rect 58985 620664 60076 620666
rect 58985 620608 58990 620664
rect 59046 620608 60076 620664
rect 58985 620606 60076 620608
rect 137093 620664 140032 620666
rect 137093 620608 137098 620664
rect 137154 620608 140032 620664
rect 137093 620606 140032 620608
rect 219249 620664 220064 620666
rect 219249 620608 219254 620664
rect 219310 620608 220064 620664
rect 583520 620652 584960 620742
rect 219249 620606 220064 620608
rect 58985 620603 59051 620606
rect 137093 620603 137159 620606
rect 219249 620603 219315 620606
rect 121913 619986 121979 619989
rect 201861 619986 201927 619989
rect 283373 619986 283439 619989
rect 120796 619984 121979 619986
rect 120796 619928 121918 619984
rect 121974 619928 121979 619984
rect 120796 619926 121979 619928
rect 200836 619984 201927 619986
rect 200836 619928 201866 619984
rect 201922 619928 201927 619984
rect 200836 619926 201927 619928
rect 280876 619984 283439 619986
rect 280876 619928 283378 619984
rect 283434 619928 283439 619984
rect 280876 619926 283439 619928
rect 121913 619923 121979 619926
rect 201861 619923 201927 619926
rect 283373 619923 283439 619926
rect 457437 618218 457503 618221
rect 457437 618216 460122 618218
rect 457437 618160 457442 618216
rect 457498 618160 460122 618216
rect 457437 618158 460122 618160
rect 457437 618155 457503 618158
rect 460062 617712 460122 618158
rect 430573 617402 430639 617405
rect 428812 617400 430639 617402
rect 428812 617344 430578 617400
rect 430634 617344 430639 617400
rect 428812 617342 430639 617344
rect 430573 617339 430639 617342
rect 58525 617266 58591 617269
rect 137001 617266 137067 617269
rect 217593 617266 217659 617269
rect 58525 617264 60076 617266
rect 58525 617208 58530 617264
rect 58586 617208 60076 617264
rect 58525 617206 60076 617208
rect 137001 617264 140032 617266
rect 137001 617208 137006 617264
rect 137062 617208 140032 617264
rect 137001 617206 140032 617208
rect 217593 617264 220064 617266
rect 217593 617208 217598 617264
rect 217654 617208 220064 617264
rect 217593 617206 220064 617208
rect 58525 617203 58591 617206
rect 137001 617203 137067 617206
rect 217593 617203 217659 617206
rect 317413 616722 317479 616725
rect 317413 616720 320068 616722
rect 317413 616664 317418 616720
rect 317474 616664 320068 616720
rect 317413 616662 320068 616664
rect 317413 616659 317479 616662
rect 123201 616586 123267 616589
rect 203149 616586 203215 616589
rect 283281 616586 283347 616589
rect 120796 616584 123267 616586
rect 120796 616528 123206 616584
rect 123262 616528 123267 616584
rect 120796 616526 123267 616528
rect 200836 616584 203215 616586
rect 200836 616528 203154 616584
rect 203210 616528 203215 616584
rect 200836 616526 203215 616528
rect 280876 616584 283347 616586
rect 280876 616528 283286 616584
rect 283342 616528 283347 616584
rect 280876 616526 283347 616528
rect 123201 616523 123267 616526
rect 203149 616523 203215 616526
rect 283281 616523 283347 616526
rect 59261 614546 59327 614549
rect 137553 614546 137619 614549
rect 217777 614546 217843 614549
rect 59261 614544 60076 614546
rect 59261 614488 59266 614544
rect 59322 614488 60076 614544
rect 59261 614486 60076 614488
rect 137553 614544 140032 614546
rect 137553 614488 137558 614544
rect 137614 614488 140032 614544
rect 137553 614486 140032 614488
rect 217777 614544 220064 614546
rect 217777 614488 217782 614544
rect 217838 614488 220064 614544
rect 217777 614486 220064 614488
rect 59261 614483 59327 614486
rect 137553 614483 137619 614486
rect 217777 614483 217843 614486
rect 509926 614138 509986 614312
rect 511993 614138 512059 614141
rect 509926 614136 512059 614138
rect 509926 614080 511998 614136
rect 512054 614080 512059 614136
rect 509926 614078 512059 614080
rect 511993 614075 512059 614078
rect 122005 613866 122071 613869
rect 283097 613866 283163 613869
rect 120796 613864 122071 613866
rect 120796 613808 122010 613864
rect 122066 613808 122071 613864
rect 280876 613864 283163 613866
rect 120796 613806 122071 613808
rect 122005 613803 122071 613806
rect 200806 613325 200866 613836
rect 280876 613808 283102 613864
rect 283158 613808 283163 613864
rect 280876 613806 283163 613808
rect 283097 613803 283163 613806
rect 200757 613320 200866 613325
rect 200757 613264 200762 613320
rect 200818 613264 200866 613320
rect 200757 613262 200866 613264
rect 200757 613259 200823 613262
rect 430665 612642 430731 612645
rect 428812 612640 430731 612642
rect 428812 612584 430670 612640
rect 430726 612584 430731 612640
rect 428812 612582 430731 612584
rect 430665 612579 430731 612582
rect 317965 611962 318031 611965
rect 317965 611960 320068 611962
rect 317965 611904 317970 611960
rect 318026 611904 320068 611960
rect 317965 611902 320068 611904
rect 317965 611899 318031 611902
rect 57881 611146 57947 611149
rect 137277 611146 137343 611149
rect 137921 611146 137987 611149
rect 218697 611146 218763 611149
rect 57881 611144 60076 611146
rect 57881 611088 57886 611144
rect 57942 611088 60076 611144
rect 57881 611086 60076 611088
rect 137277 611144 140032 611146
rect 137277 611088 137282 611144
rect 137338 611088 137926 611144
rect 137982 611088 140032 611144
rect 137277 611086 140032 611088
rect 218697 611144 220064 611146
rect 218697 611088 218702 611144
rect 218758 611088 220064 611144
rect 218697 611086 220064 611088
rect 57881 611083 57947 611086
rect 137277 611083 137343 611086
rect 137921 611083 137987 611086
rect 218697 611083 218763 611086
rect 123109 610466 123175 610469
rect 203057 610466 203123 610469
rect 120796 610464 123175 610466
rect 120796 610408 123114 610464
rect 123170 610408 123175 610464
rect 120796 610406 123175 610408
rect 200836 610464 203123 610466
rect 200836 610408 203062 610464
rect 203118 610408 203123 610464
rect 200836 610406 203123 610408
rect 123109 610403 123175 610406
rect 203057 610403 203123 610406
rect 280846 610061 280906 610436
rect 280846 610056 280955 610061
rect 280846 610000 280894 610056
rect 280950 610000 280955 610056
rect 280846 609998 280955 610000
rect 280889 609995 280955 609998
rect -960 609650 480 609740
rect 2773 609650 2839 609653
rect -960 609648 2839 609650
rect -960 609592 2778 609648
rect 2834 609592 2839 609648
rect -960 609590 2839 609592
rect -960 609500 480 609590
rect 2773 609587 2839 609590
rect 457437 608970 457503 608973
rect 460062 608970 460122 609552
rect 457437 608968 460122 608970
rect 457437 608912 457442 608968
rect 457498 608912 460122 608968
rect 457437 608910 460122 608912
rect 457437 608907 457503 608910
rect 57513 608426 57579 608429
rect 138933 608426 138999 608429
rect 217409 608426 217475 608429
rect 57513 608424 60076 608426
rect 57513 608368 57518 608424
rect 57574 608368 60076 608424
rect 57513 608366 60076 608368
rect 138933 608424 140032 608426
rect 138933 608368 138938 608424
rect 138994 608368 140032 608424
rect 138933 608366 140032 608368
rect 217409 608424 220064 608426
rect 217409 608368 217414 608424
rect 217470 608368 220064 608424
rect 217409 608366 220064 608368
rect 57513 608363 57579 608366
rect 138933 608363 138999 608366
rect 217409 608363 217475 608366
rect 580257 608018 580323 608021
rect 583520 608018 584960 608108
rect 580257 608016 584960 608018
rect 580257 607960 580262 608016
rect 580318 607960 584960 608016
rect 580257 607958 584960 607960
rect 580257 607955 580323 607958
rect 430798 607882 430804 607884
rect 428812 607822 430804 607882
rect 430798 607820 430804 607822
rect 430868 607820 430874 607884
rect 583520 607868 584960 607958
rect 123293 607746 123359 607749
rect 202873 607746 202939 607749
rect 283189 607746 283255 607749
rect 120796 607744 123359 607746
rect 120796 607688 123298 607744
rect 123354 607688 123359 607744
rect 120796 607686 123359 607688
rect 200836 607744 202939 607746
rect 200836 607688 202878 607744
rect 202934 607688 202939 607744
rect 200836 607686 202939 607688
rect 280876 607744 283255 607746
rect 280876 607688 283194 607744
rect 283250 607688 283255 607744
rect 280876 607686 283255 607688
rect 123293 607683 123359 607686
rect 202873 607683 202939 607686
rect 283189 607683 283255 607686
rect 318793 607202 318859 607205
rect 318793 607200 320068 607202
rect 318793 607144 318798 607200
rect 318854 607144 320068 607200
rect 318793 607142 320068 607144
rect 318793 607139 318859 607142
rect 509926 605978 509986 606152
rect 512085 605978 512151 605981
rect 509926 605976 512151 605978
rect 509926 605920 512090 605976
rect 512146 605920 512151 605976
rect 509926 605918 512151 605920
rect 512085 605915 512151 605918
rect 58801 605026 58867 605029
rect 137369 605026 137435 605029
rect 216673 605026 216739 605029
rect 58801 605024 60076 605026
rect 58801 604968 58806 605024
rect 58862 604968 60076 605024
rect 58801 604966 60076 604968
rect 137369 605024 140032 605026
rect 137369 604968 137374 605024
rect 137430 604968 140032 605024
rect 137369 604966 140032 604968
rect 216673 605024 220064 605026
rect 216673 604968 216678 605024
rect 216734 604968 220064 605024
rect 216673 604966 220064 604968
rect 58801 604963 58867 604966
rect 137369 604963 137435 604966
rect 216673 604963 216739 604966
rect 124121 604346 124187 604349
rect 203885 604346 203951 604349
rect 283649 604346 283715 604349
rect 120796 604344 124187 604346
rect 120796 604288 124126 604344
rect 124182 604288 124187 604344
rect 120796 604286 124187 604288
rect 200836 604344 203951 604346
rect 200836 604288 203890 604344
rect 203946 604288 203951 604344
rect 200836 604286 203951 604288
rect 280876 604344 283715 604346
rect 280876 604288 283654 604344
rect 283710 604288 283715 604344
rect 280876 604286 283715 604288
rect 124121 604283 124187 604286
rect 203885 604283 203951 604286
rect 283649 604283 283715 604286
rect 430757 603122 430823 603125
rect 428812 603120 430823 603122
rect 428812 603064 430762 603120
rect 430818 603064 430823 603120
rect 428812 603062 430823 603064
rect 430757 603059 430823 603062
rect 317965 602442 318031 602445
rect 317965 602440 320068 602442
rect 317965 602384 317970 602440
rect 318026 602384 320068 602440
rect 317965 602382 320068 602384
rect 317965 602379 318031 602382
rect 57237 602306 57303 602309
rect 137369 602306 137435 602309
rect 216673 602306 216739 602309
rect 57237 602304 60076 602306
rect 57237 602248 57242 602304
rect 57298 602248 60076 602304
rect 57237 602246 60076 602248
rect 137369 602304 140032 602306
rect 137369 602248 137374 602304
rect 137430 602248 140032 602304
rect 137369 602246 140032 602248
rect 216673 602304 220064 602306
rect 216673 602248 216678 602304
rect 216734 602248 220064 602304
rect 216673 602246 220064 602248
rect 57237 602243 57303 602246
rect 137369 602243 137435 602246
rect 216673 602243 216739 602246
rect 123385 601626 123451 601629
rect 202137 601626 202203 601629
rect 281901 601626 281967 601629
rect 120796 601624 123451 601626
rect 120796 601568 123390 601624
rect 123446 601568 123451 601624
rect 120796 601566 123451 601568
rect 200836 601624 202203 601626
rect 200836 601568 202142 601624
rect 202198 601568 202203 601624
rect 200836 601566 202203 601568
rect 280876 601624 281967 601626
rect 280876 601568 281906 601624
rect 281962 601568 281967 601624
rect 280876 601566 281967 601568
rect 123385 601563 123451 601566
rect 202137 601563 202203 601566
rect 281901 601563 281967 601566
rect 457529 600810 457595 600813
rect 460062 600810 460122 601392
rect 457529 600808 460122 600810
rect 457529 600752 457534 600808
rect 457590 600752 460122 600808
rect 457529 600750 460122 600752
rect 457529 600747 457595 600750
rect 57329 598906 57395 598909
rect 138841 598906 138907 598909
rect 217041 598906 217107 598909
rect 57329 598904 60076 598906
rect 57329 598848 57334 598904
rect 57390 598848 60076 598904
rect 57329 598846 60076 598848
rect 138841 598904 140032 598906
rect 138841 598848 138846 598904
rect 138902 598848 140032 598904
rect 138841 598846 140032 598848
rect 217041 598904 220064 598906
rect 217041 598848 217046 598904
rect 217102 598848 220064 598904
rect 217041 598846 220064 598848
rect 57329 598843 57395 598846
rect 138841 598843 138907 598846
rect 217041 598843 217107 598846
rect 429193 598362 429259 598365
rect 428812 598360 429259 598362
rect 428812 598304 429198 598360
rect 429254 598304 429259 598360
rect 428812 598302 429259 598304
rect 429193 598299 429259 598302
rect 203241 598226 203307 598229
rect 281993 598226 282059 598229
rect 200836 598224 203307 598226
rect 120766 597682 120826 598196
rect 200836 598168 203246 598224
rect 203302 598168 203307 598224
rect 200836 598166 203307 598168
rect 280876 598224 282059 598226
rect 280876 598168 281998 598224
rect 282054 598168 282059 598224
rect 280876 598166 282059 598168
rect 203241 598163 203307 598166
rect 281993 598163 282059 598166
rect 120993 597682 121059 597685
rect 120766 597680 121059 597682
rect 120766 597624 120998 597680
rect 121054 597624 121059 597680
rect 120766 597622 121059 597624
rect 120993 597619 121059 597622
rect 317965 597682 318031 597685
rect 509926 597682 509986 597992
rect 511257 597682 511323 597685
rect 317965 597680 320068 597682
rect 317965 597624 317970 597680
rect 318026 597624 320068 597680
rect 317965 597622 320068 597624
rect 509926 597680 511323 597682
rect 509926 597624 511262 597680
rect 511318 597624 511323 597680
rect 509926 597622 511323 597624
rect 317965 597619 318031 597622
rect 511257 597619 511323 597622
rect -960 596988 480 597228
rect 57421 596186 57487 596189
rect 137461 596186 137527 596189
rect 217777 596186 217843 596189
rect 57421 596184 60076 596186
rect 57421 596128 57426 596184
rect 57482 596128 60076 596184
rect 57421 596126 60076 596128
rect 137461 596184 140032 596186
rect 137461 596128 137466 596184
rect 137522 596128 140032 596184
rect 137461 596126 140032 596128
rect 217777 596184 220064 596186
rect 217777 596128 217782 596184
rect 217838 596128 220064 596184
rect 217777 596126 220064 596128
rect 57421 596123 57487 596126
rect 137461 596123 137527 596126
rect 217777 596123 217843 596126
rect 122097 595506 122163 595509
rect 202045 595506 202111 595509
rect 281809 595506 281875 595509
rect 120796 595504 122163 595506
rect 120796 595448 122102 595504
rect 122158 595448 122163 595504
rect 120796 595446 122163 595448
rect 200836 595504 202111 595506
rect 200836 595448 202050 595504
rect 202106 595448 202111 595504
rect 200836 595446 202111 595448
rect 280876 595504 281875 595506
rect 280876 595448 281814 595504
rect 281870 595448 281875 595504
rect 280876 595446 281875 595448
rect 122097 595443 122163 595446
rect 202045 595443 202111 595446
rect 281809 595443 281875 595446
rect 583520 595084 584960 595324
rect 429377 593602 429443 593605
rect 428812 593600 429443 593602
rect 428812 593544 429382 593600
rect 429438 593544 429443 593600
rect 428812 593542 429443 593544
rect 429377 593539 429443 593542
rect 317965 592922 318031 592925
rect 317965 592920 320068 592922
rect 317965 592864 317970 592920
rect 318026 592864 320068 592920
rect 317965 592862 320068 592864
rect 317965 592859 318031 592862
rect 59261 592786 59327 592789
rect 136633 592786 136699 592789
rect 216673 592786 216739 592789
rect 59261 592784 60076 592786
rect 59261 592728 59266 592784
rect 59322 592728 60076 592784
rect 59261 592726 60076 592728
rect 136633 592784 140032 592786
rect 136633 592728 136638 592784
rect 136694 592728 140032 592784
rect 136633 592726 140032 592728
rect 216673 592784 220064 592786
rect 216673 592728 216678 592784
rect 216734 592728 220064 592784
rect 216673 592726 220064 592728
rect 59261 592723 59327 592726
rect 136633 592723 136699 592726
rect 216673 592723 216739 592726
rect 457621 592650 457687 592653
rect 460062 592650 460122 593232
rect 457621 592648 460122 592650
rect 457621 592592 457626 592648
rect 457682 592592 460122 592648
rect 457621 592590 460122 592592
rect 457621 592587 457687 592590
rect 123477 592106 123543 592109
rect 201033 592106 201099 592109
rect 282913 592106 282979 592109
rect 120796 592104 123543 592106
rect 120796 592048 123482 592104
rect 123538 592048 123543 592104
rect 120796 592046 123543 592048
rect 200836 592104 201099 592106
rect 200836 592048 201038 592104
rect 201094 592048 201099 592104
rect 200836 592046 201099 592048
rect 280876 592104 282979 592106
rect 280876 592048 282918 592104
rect 282974 592048 282979 592104
rect 280876 592046 282979 592048
rect 123477 592043 123543 592046
rect 201033 592043 201099 592046
rect 282913 592043 282979 592046
rect 58433 590066 58499 590069
rect 136633 590066 136699 590069
rect 216673 590066 216739 590069
rect 58433 590064 60076 590066
rect 58433 590008 58438 590064
rect 58494 590008 60076 590064
rect 58433 590006 60076 590008
rect 136633 590064 140032 590066
rect 136633 590008 136638 590064
rect 136694 590008 140032 590064
rect 136633 590006 140032 590008
rect 216673 590064 220064 590066
rect 216673 590008 216678 590064
rect 216734 590008 220064 590064
rect 216673 590006 220064 590008
rect 58433 590003 58499 590006
rect 136633 590003 136699 590006
rect 216673 590003 216739 590006
rect 121545 589386 121611 589389
rect 203333 589386 203399 589389
rect 281165 589386 281231 589389
rect 120796 589384 121611 589386
rect 120796 589328 121550 589384
rect 121606 589328 121611 589384
rect 120796 589326 121611 589328
rect 200836 589384 203399 589386
rect 200836 589328 203338 589384
rect 203394 589328 203399 589384
rect 200836 589326 203399 589328
rect 280876 589384 281231 589386
rect 280876 589328 281170 589384
rect 281226 589328 281231 589384
rect 280876 589326 281231 589328
rect 509926 589386 509986 589832
rect 512177 589386 512243 589389
rect 509926 589384 512243 589386
rect 509926 589328 512182 589384
rect 512238 589328 512243 589384
rect 509926 589326 512243 589328
rect 121545 589323 121611 589326
rect 203333 589323 203399 589326
rect 281165 589323 281231 589326
rect 512177 589323 512243 589326
rect 429469 588162 429535 588165
rect 428812 588160 429535 588162
rect 428812 588104 429474 588160
rect 429530 588104 429535 588160
rect 428812 588102 429535 588104
rect 429469 588099 429535 588102
rect 57145 586666 57211 586669
rect 139301 586666 139367 586669
rect 216673 586666 216739 586669
rect 57145 586664 60076 586666
rect 57145 586608 57150 586664
rect 57206 586608 60076 586664
rect 57145 586606 60076 586608
rect 139301 586664 140032 586666
rect 139301 586608 139306 586664
rect 139362 586608 140032 586664
rect 139301 586606 140032 586608
rect 216673 586664 220064 586666
rect 216673 586608 216678 586664
rect 216734 586608 220064 586664
rect 216673 586606 220064 586608
rect 57145 586603 57211 586606
rect 139301 586603 139367 586606
rect 216673 586603 216739 586606
rect 317413 586530 317479 586533
rect 317413 586528 317522 586530
rect 317413 586472 317418 586528
rect 317474 586472 317522 586528
rect 317413 586467 317522 586472
rect 317462 586394 317522 586467
rect 320038 586394 320098 587452
rect 317462 586334 320098 586394
rect 122281 585986 122347 585989
rect 202229 585986 202295 585989
rect 283557 585986 283623 585989
rect 120796 585984 122347 585986
rect 120796 585928 122286 585984
rect 122342 585928 122347 585984
rect 120796 585926 122347 585928
rect 200836 585984 202295 585986
rect 200836 585928 202234 585984
rect 202290 585928 202295 585984
rect 200836 585926 202295 585928
rect 280876 585984 283623 585986
rect 280876 585928 283562 585984
rect 283618 585928 283623 585984
rect 280876 585926 283623 585928
rect 122281 585923 122347 585926
rect 202229 585923 202295 585926
rect 283557 585923 283623 585926
rect -960 584490 480 584580
rect 3509 584490 3575 584493
rect -960 584488 3575 584490
rect -960 584432 3514 584488
rect 3570 584432 3575 584488
rect -960 584430 3575 584432
rect -960 584340 480 584430
rect 3509 584427 3575 584430
rect 58709 583946 58775 583949
rect 137921 583946 137987 583949
rect 219157 583946 219223 583949
rect 58709 583944 60076 583946
rect 58709 583888 58714 583944
rect 58770 583888 60076 583944
rect 58709 583886 60076 583888
rect 137921 583944 140032 583946
rect 137921 583888 137926 583944
rect 137982 583888 140032 583944
rect 137921 583886 140032 583888
rect 219157 583944 220064 583946
rect 219157 583888 219162 583944
rect 219218 583888 220064 583944
rect 219157 583886 220064 583888
rect 58709 583883 58775 583886
rect 137921 583883 137987 583886
rect 219157 583883 219223 583886
rect 430849 583402 430915 583405
rect 428812 583400 430915 583402
rect 428812 583344 430854 583400
rect 430910 583344 430915 583400
rect 428812 583342 430915 583344
rect 430849 583339 430915 583342
rect 123569 583266 123635 583269
rect 201125 583266 201191 583269
rect 281625 583266 281691 583269
rect 120796 583264 123635 583266
rect 120796 583208 123574 583264
rect 123630 583208 123635 583264
rect 120796 583206 123635 583208
rect 200836 583264 201191 583266
rect 200836 583208 201130 583264
rect 201186 583208 201191 583264
rect 200836 583206 201191 583208
rect 280876 583264 281691 583266
rect 280876 583208 281630 583264
rect 281686 583208 281691 583264
rect 280876 583206 281691 583208
rect 123569 583203 123635 583206
rect 201125 583203 201191 583206
rect 281625 583203 281691 583206
rect 316677 582722 316743 582725
rect 316677 582720 320068 582722
rect 316677 582664 316682 582720
rect 316738 582664 320068 582720
rect 316677 582662 320068 582664
rect 316677 582659 316743 582662
rect 583520 582164 584960 582404
rect 57053 580546 57119 580549
rect 138565 580546 138631 580549
rect 218145 580546 218211 580549
rect 57053 580544 60076 580546
rect 57053 580488 57058 580544
rect 57114 580488 60076 580544
rect 57053 580486 60076 580488
rect 138565 580544 140032 580546
rect 138565 580488 138570 580544
rect 138626 580488 140032 580544
rect 138565 580486 140032 580488
rect 218145 580544 220064 580546
rect 218145 580488 218150 580544
rect 218206 580488 220064 580544
rect 218145 580486 220064 580488
rect 57053 580483 57119 580486
rect 138565 580483 138631 580486
rect 218145 580483 218211 580486
rect 121085 579866 121151 579869
rect 203425 579866 203491 579869
rect 281257 579866 281323 579869
rect 120796 579864 121151 579866
rect 120796 579808 121090 579864
rect 121146 579808 121151 579864
rect 120796 579806 121151 579808
rect 200836 579864 203491 579866
rect 200836 579808 203430 579864
rect 203486 579808 203491 579864
rect 200836 579806 203491 579808
rect 280876 579864 281323 579866
rect 280876 579808 281262 579864
rect 281318 579808 281323 579864
rect 280876 579806 281323 579808
rect 121085 579803 121151 579806
rect 203425 579803 203491 579806
rect 281257 579803 281323 579806
rect 430941 578642 431007 578645
rect 428812 578640 431007 578642
rect 428812 578584 430946 578640
rect 431002 578584 431007 578640
rect 428812 578582 431007 578584
rect 430941 578579 431007 578582
rect 317505 577962 317571 577965
rect 317505 577960 320068 577962
rect 317505 577904 317510 577960
rect 317566 577904 320068 577960
rect 317505 577902 320068 577904
rect 317505 577899 317571 577902
rect 138473 577826 138539 577829
rect 216673 577826 216739 577829
rect 138473 577824 140032 577826
rect 59537 577790 59603 577793
rect 59537 577788 60076 577790
rect 59537 577732 59542 577788
rect 59598 577732 60076 577788
rect 138473 577768 138478 577824
rect 138534 577768 140032 577824
rect 138473 577766 140032 577768
rect 216673 577824 220064 577826
rect 216673 577768 216678 577824
rect 216734 577768 220064 577824
rect 216673 577766 220064 577768
rect 138473 577763 138539 577766
rect 216673 577763 216739 577766
rect 59537 577730 60076 577732
rect 59537 577727 59603 577730
rect 121177 577146 121243 577149
rect 201217 577146 201283 577149
rect 281533 577146 281599 577149
rect 120796 577144 121243 577146
rect 120796 577088 121182 577144
rect 121238 577088 121243 577144
rect 120796 577086 121243 577088
rect 200836 577144 201283 577146
rect 200836 577088 201222 577144
rect 201278 577088 201283 577144
rect 200836 577086 201283 577088
rect 280876 577144 281599 577146
rect 280876 577088 281538 577144
rect 281594 577088 281599 577144
rect 280876 577086 281599 577088
rect 121177 577083 121243 577086
rect 201217 577083 201283 577086
rect 281533 577083 281599 577086
rect 428414 573341 428474 573852
rect 428365 573336 428474 573341
rect 428365 573280 428370 573336
rect 428426 573280 428474 573336
rect 428365 573278 428474 573280
rect 428365 573275 428431 573278
rect 317965 573202 318031 573205
rect 317965 573200 320068 573202
rect 317965 573144 317970 573200
rect 318026 573144 320068 573200
rect 317965 573142 320068 573144
rect 317965 573139 318031 573142
rect -960 571828 480 572068
rect 580901 569530 580967 569533
rect 583520 569530 584960 569620
rect 580901 569528 584960 569530
rect 580901 569472 580906 569528
rect 580962 569472 584960 569528
rect 580901 569470 584960 569472
rect 580901 569467 580967 569470
rect 583520 569380 584960 569470
rect 431033 569122 431099 569125
rect 428812 569120 431099 569122
rect 428812 569064 431038 569120
rect 431094 569064 431099 569120
rect 428812 569062 431099 569064
rect 431033 569059 431099 569062
rect 317965 568442 318031 568445
rect 317965 568440 320068 568442
rect 317965 568384 317970 568440
rect 318026 568384 320068 568440
rect 317965 568382 320068 568384
rect 317965 568379 318031 568382
rect 428414 563821 428474 564332
rect 428414 563816 428523 563821
rect 428414 563760 428462 563816
rect 428518 563760 428523 563816
rect 428414 563758 428523 563760
rect 428457 563755 428523 563758
rect 317965 563682 318031 563685
rect 317965 563680 320068 563682
rect 317965 563624 317970 563680
rect 318026 563624 320068 563680
rect 317965 563622 320068 563624
rect 317965 563619 318031 563622
rect 431125 559602 431191 559605
rect 428812 559600 431191 559602
rect 428812 559544 431130 559600
rect 431186 559544 431191 559600
rect 428812 559542 431191 559544
rect 431125 559539 431191 559542
rect -960 559330 480 559420
rect 2773 559330 2839 559333
rect -960 559328 2839 559330
rect -960 559272 2778 559328
rect 2834 559272 2839 559328
rect -960 559270 2839 559272
rect -960 559180 480 559270
rect 2773 559267 2839 559270
rect 317965 558922 318031 558925
rect 317965 558920 320068 558922
rect 317965 558864 317970 558920
rect 318026 558864 320068 558920
rect 317965 558862 320068 558864
rect 317965 558859 318031 558862
rect 217593 557562 217659 557565
rect 217961 557562 218027 557565
rect 217593 557560 218027 557562
rect 217593 557504 217598 557560
rect 217654 557504 217966 557560
rect 218022 557504 218027 557560
rect 217593 557502 218027 557504
rect 217593 557499 217659 557502
rect 217961 557499 218027 557502
rect 248689 556746 248755 556749
rect 300669 556746 300735 556749
rect 248689 556744 300735 556746
rect 248689 556688 248694 556744
rect 248750 556688 300674 556744
rect 300730 556688 300735 556744
rect 248689 556686 300735 556688
rect 248689 556683 248755 556686
rect 300669 556683 300735 556686
rect 580165 556746 580231 556749
rect 583520 556746 584960 556836
rect 580165 556744 584960 556746
rect 580165 556688 580170 556744
rect 580226 556688 584960 556744
rect 580165 556686 584960 556688
rect 580165 556683 580231 556686
rect 258717 556610 258783 556613
rect 303153 556610 303219 556613
rect 258717 556608 303219 556610
rect 258717 556552 258722 556608
rect 258778 556552 303158 556608
rect 303214 556552 303219 556608
rect 583520 556596 584960 556686
rect 258717 556550 303219 556552
rect 258717 556547 258783 556550
rect 303153 556547 303219 556550
rect 255129 556474 255195 556477
rect 300485 556474 300551 556477
rect 255129 556472 300551 556474
rect 255129 556416 255134 556472
rect 255190 556416 300490 556472
rect 300546 556416 300551 556472
rect 255129 556414 300551 556416
rect 255129 556411 255195 556414
rect 300485 556411 300551 556414
rect 290917 556338 290983 556341
rect 318333 556338 318399 556341
rect 290917 556336 318399 556338
rect 290917 556280 290922 556336
rect 290978 556280 318338 556336
rect 318394 556280 318399 556336
rect 290917 556278 318399 556280
rect 290917 556275 290983 556278
rect 318333 556275 318399 556278
rect 241513 556202 241579 556205
rect 319897 556202 319963 556205
rect 241513 556200 319963 556202
rect 241513 556144 241518 556200
rect 241574 556144 319902 556200
rect 319958 556144 319963 556200
rect 241513 556142 319963 556144
rect 241513 556139 241579 556142
rect 319897 556139 319963 556142
rect 3417 554842 3483 554845
rect 318517 554842 318583 554845
rect 431217 554842 431283 554845
rect 3417 554840 318583 554842
rect 3417 554784 3422 554840
rect 3478 554784 318522 554840
rect 318578 554784 318583 554840
rect 3417 554782 318583 554784
rect 428812 554840 431283 554842
rect 428812 554784 431222 554840
rect 431278 554784 431283 554840
rect 428812 554782 431283 554784
rect 3417 554779 3483 554782
rect 318517 554779 318583 554782
rect 431217 554779 431283 554782
rect 317965 554162 318031 554165
rect 317965 554160 320068 554162
rect 317965 554104 317970 554160
rect 318026 554104 320068 554160
rect 317965 554102 320068 554104
rect 317965 554099 318031 554102
rect 431309 550082 431375 550085
rect 428812 550080 431375 550082
rect 428812 550024 431314 550080
rect 431370 550024 431375 550080
rect 428812 550022 431375 550024
rect 431309 550019 431375 550022
rect 317413 549402 317479 549405
rect 317413 549400 320068 549402
rect 317413 549344 317418 549400
rect 317474 549344 320068 549400
rect 317413 549342 320068 549344
rect 317413 549339 317479 549342
rect 303245 547498 303311 547501
rect 299828 547496 303311 547498
rect 299828 547440 303250 547496
rect 303306 547440 303311 547496
rect 299828 547438 303311 547440
rect 303245 547435 303311 547438
rect -960 546668 480 546908
rect 429285 545322 429351 545325
rect 428812 545320 429351 545322
rect 428812 545264 429290 545320
rect 429346 545264 429351 545320
rect 428812 545262 429351 545264
rect 429285 545259 429351 545262
rect 317965 544642 318031 544645
rect 317965 544640 320068 544642
rect 317965 544584 317970 544640
rect 318026 544584 320068 544640
rect 317965 544582 320068 544584
rect 317965 544579 318031 544582
rect 583520 543812 584960 544052
rect 430573 540562 430639 540565
rect 428812 540560 430639 540562
rect 428812 540504 430578 540560
rect 430634 540504 430639 540560
rect 428812 540502 430639 540504
rect 430573 540499 430639 540502
rect 318701 539882 318767 539885
rect 318701 539880 320068 539882
rect 318701 539824 318706 539880
rect 318762 539824 320068 539880
rect 318701 539822 320068 539824
rect 318701 539819 318767 539822
rect 428549 535938 428615 535941
rect 428549 535936 428658 535938
rect 428549 535880 428554 535936
rect 428610 535880 428658 535936
rect 428549 535875 428658 535880
rect 428598 535772 428658 535875
rect 303153 535530 303219 535533
rect 430614 535530 430620 535532
rect 303153 535528 430620 535530
rect 303153 535472 303158 535528
rect 303214 535472 430620 535528
rect 303153 535470 430620 535472
rect 303153 535467 303219 535470
rect 430614 535468 430620 535470
rect 430684 535468 430690 535532
rect 319897 535394 319963 535397
rect 430798 535394 430804 535396
rect 319897 535392 430804 535394
rect 319897 535336 319902 535392
rect 319958 535336 430804 535392
rect 319897 535334 430804 535336
rect 319897 535331 319963 535334
rect 430798 535332 430804 535334
rect 430868 535332 430874 535396
rect -960 534156 480 534396
rect 324865 534034 324931 534037
rect 436737 534034 436803 534037
rect 324865 534032 436803 534034
rect 324865 533976 324870 534032
rect 324926 533976 436742 534032
rect 436798 533976 436803 534032
rect 324865 533974 436803 533976
rect 324865 533971 324931 533974
rect 436737 533971 436803 533974
rect 319713 532674 319779 532677
rect 337653 532674 337719 532677
rect 319713 532672 337719 532674
rect 319713 532616 319718 532672
rect 319774 532616 337658 532672
rect 337714 532616 337719 532672
rect 319713 532614 337719 532616
rect 319713 532611 319779 532614
rect 337653 532611 337719 532614
rect 302325 532538 302391 532541
rect 299828 532536 302391 532538
rect 299828 532480 302330 532536
rect 302386 532480 302391 532536
rect 299828 532478 302391 532480
rect 302325 532475 302391 532478
rect 583520 531028 584960 531268
rect 57697 525058 57763 525061
rect 57697 525056 60076 525058
rect 57697 525000 57702 525056
rect 57758 525000 60076 525056
rect 57697 524998 60076 525000
rect 57697 524995 57763 524998
rect -960 521658 480 521748
rect 3417 521658 3483 521661
rect -960 521656 3483 521658
rect -960 521600 3422 521656
rect 3478 521600 3483 521656
rect -960 521598 3483 521600
rect -960 521508 480 521598
rect 3417 521595 3483 521598
rect 580901 518394 580967 518397
rect 583520 518394 584960 518484
rect 580901 518392 584960 518394
rect 580901 518336 580906 518392
rect 580962 518336 584960 518392
rect 580901 518334 584960 518336
rect 580901 518331 580967 518334
rect 583520 518244 584960 518334
rect 302969 517578 303035 517581
rect 299828 517576 303035 517578
rect 299828 517520 302974 517576
rect 303030 517520 303035 517576
rect 299828 517518 303035 517520
rect 302969 517515 303035 517518
rect -960 509146 480 509236
rect 2773 509146 2839 509149
rect -960 509144 2839 509146
rect -960 509088 2778 509144
rect 2834 509088 2839 509144
rect -960 509086 2839 509088
rect -960 508996 480 509086
rect 2773 509083 2839 509086
rect 583520 505460 584960 505700
rect 302877 502618 302943 502621
rect 299828 502616 302943 502618
rect 299828 502560 302882 502616
rect 302938 502560 302943 502616
rect 299828 502558 302943 502560
rect 302877 502555 302943 502558
rect -960 496348 480 496588
rect 580165 492826 580231 492829
rect 583520 492826 584960 492916
rect 580165 492824 584960 492826
rect 580165 492768 580170 492824
rect 580226 492768 584960 492824
rect 580165 492766 584960 492768
rect 580165 492763 580231 492766
rect 583520 492676 584960 492766
rect 59302 492492 59308 492556
rect 59372 492554 59378 492556
rect 72877 492554 72943 492557
rect 59372 492552 72943 492554
rect 59372 492496 72882 492552
rect 72938 492496 72943 492552
rect 59372 492494 72943 492496
rect 59372 492492 59378 492494
rect 72877 492491 72943 492494
rect 185761 492554 185827 492557
rect 196566 492554 196572 492556
rect 185761 492552 196572 492554
rect 185761 492496 185766 492552
rect 185822 492496 196572 492552
rect 185761 492494 196572 492496
rect 185761 492491 185827 492494
rect 196566 492492 196572 492494
rect 196636 492492 196642 492556
rect 212809 492554 212875 492557
rect 213310 492554 213316 492556
rect 212809 492552 213316 492554
rect 212809 492496 212814 492552
rect 212870 492496 213316 492552
rect 212809 492494 213316 492496
rect 212809 492491 212875 492494
rect 213310 492492 213316 492494
rect 213380 492492 213386 492556
rect 217358 492492 217364 492556
rect 217428 492554 217434 492556
rect 217777 492554 217843 492557
rect 217428 492552 217843 492554
rect 217428 492496 217782 492552
rect 217838 492496 217843 492552
rect 217428 492494 217843 492496
rect 217428 492492 217434 492494
rect 217777 492491 217843 492494
rect 219934 492492 219940 492556
rect 220004 492554 220010 492556
rect 224401 492554 224467 492557
rect 220004 492552 224467 492554
rect 220004 492496 224406 492552
rect 224462 492496 224467 492552
rect 220004 492494 224467 492496
rect 220004 492492 220010 492494
rect 224401 492491 224467 492494
rect 235901 492554 235967 492557
rect 357934 492554 357940 492556
rect 235901 492552 357940 492554
rect 235901 492496 235906 492552
rect 235962 492496 357940 492552
rect 235901 492494 357940 492496
rect 235901 492491 235967 492494
rect 357934 492492 357940 492494
rect 358004 492492 358010 492556
rect 71957 492418 72023 492421
rect 77753 492418 77819 492421
rect 71957 492416 77819 492418
rect 71957 492360 71962 492416
rect 72018 492360 77758 492416
rect 77814 492360 77819 492416
rect 71957 492358 77819 492360
rect 71957 492355 72023 492358
rect 77753 492355 77819 492358
rect 150249 492418 150315 492421
rect 197854 492418 197860 492420
rect 150249 492416 197860 492418
rect 150249 492360 150254 492416
rect 150310 492360 197860 492416
rect 150249 492358 197860 492360
rect 150249 492355 150315 492358
rect 197854 492356 197860 492358
rect 197924 492356 197930 492420
rect 217225 492418 217291 492421
rect 217542 492418 217548 492420
rect 217225 492416 217548 492418
rect 217225 492360 217230 492416
rect 217286 492360 217548 492416
rect 217225 492358 217548 492360
rect 217225 492355 217291 492358
rect 217542 492356 217548 492358
rect 217612 492356 217618 492420
rect 235809 492418 235875 492421
rect 360694 492418 360700 492420
rect 235809 492416 360700 492418
rect 235809 492360 235814 492416
rect 235870 492360 360700 492416
rect 235809 492358 360700 492360
rect 235809 492355 235875 492358
rect 360694 492356 360700 492358
rect 360764 492356 360770 492420
rect 46790 492220 46796 492284
rect 46860 492282 46866 492284
rect 66161 492282 66227 492285
rect 46860 492280 66227 492282
rect 46860 492224 66166 492280
rect 66222 492224 66227 492280
rect 46860 492222 66227 492224
rect 46860 492220 46866 492222
rect 66161 492219 66227 492222
rect 68921 492282 68987 492285
rect 78581 492282 78647 492285
rect 68921 492280 78647 492282
rect 68921 492224 68926 492280
rect 68982 492224 78586 492280
rect 78642 492224 78647 492280
rect 68921 492222 78647 492224
rect 68921 492219 68987 492222
rect 78581 492219 78647 492222
rect 147765 492282 147831 492285
rect 191189 492282 191255 492285
rect 147765 492280 191255 492282
rect 147765 492224 147770 492280
rect 147826 492224 191194 492280
rect 191250 492224 191255 492280
rect 147765 492222 191255 492224
rect 147765 492219 147831 492222
rect 191189 492219 191255 492222
rect 200849 492282 200915 492285
rect 201350 492282 201356 492284
rect 200849 492280 201356 492282
rect 200849 492224 200854 492280
rect 200910 492224 201356 492280
rect 200849 492222 201356 492224
rect 200849 492219 200915 492222
rect 201350 492220 201356 492222
rect 201420 492220 201426 492284
rect 201769 492282 201835 492285
rect 202638 492282 202644 492284
rect 201769 492280 202644 492282
rect 201769 492224 201774 492280
rect 201830 492224 202644 492280
rect 201769 492222 202644 492224
rect 201769 492219 201835 492222
rect 202638 492220 202644 492222
rect 202708 492220 202714 492284
rect 235257 492282 235323 492285
rect 364926 492282 364932 492284
rect 235257 492280 364932 492282
rect 235257 492224 235262 492280
rect 235318 492224 364932 492280
rect 235257 492222 364932 492224
rect 235257 492219 235323 492222
rect 364926 492220 364932 492222
rect 364996 492220 365002 492284
rect 53598 492084 53604 492148
rect 53668 492146 53674 492148
rect 76005 492146 76071 492149
rect 53668 492144 76071 492146
rect 53668 492088 76010 492144
rect 76066 492088 76071 492144
rect 53668 492086 76071 492088
rect 53668 492084 53674 492086
rect 76005 492083 76071 492086
rect 149145 492146 149211 492149
rect 200665 492146 200731 492149
rect 201166 492146 201172 492148
rect 149145 492144 200498 492146
rect 149145 492088 149150 492144
rect 149206 492088 200498 492144
rect 149145 492086 200498 492088
rect 149145 492083 149211 492086
rect 50838 491948 50844 492012
rect 50908 492010 50914 492012
rect 77293 492010 77359 492013
rect 50908 492008 77359 492010
rect 50908 491952 77298 492008
rect 77354 491952 77359 492008
rect 50908 491950 77359 491952
rect 50908 491948 50914 491950
rect 77293 491947 77359 491950
rect 146569 492010 146635 492013
rect 200205 492010 200271 492013
rect 146569 492008 200271 492010
rect 146569 491952 146574 492008
rect 146630 491952 200210 492008
rect 200266 491952 200271 492008
rect 146569 491950 200271 491952
rect 200438 492010 200498 492086
rect 200665 492144 201172 492146
rect 200665 492088 200670 492144
rect 200726 492088 201172 492144
rect 200665 492086 201172 492088
rect 200665 492083 200731 492086
rect 201166 492084 201172 492086
rect 201236 492084 201242 492148
rect 205725 492146 205791 492149
rect 206870 492146 206876 492148
rect 205725 492144 206876 492146
rect 205725 492088 205730 492144
rect 205786 492088 206876 492144
rect 205725 492086 206876 492088
rect 205725 492083 205791 492086
rect 206870 492084 206876 492086
rect 206940 492084 206946 492148
rect 233233 492146 233299 492149
rect 367686 492146 367692 492148
rect 233233 492144 367692 492146
rect 233233 492088 233238 492144
rect 233294 492088 367692 492144
rect 233233 492086 367692 492088
rect 233233 492083 233299 492086
rect 367686 492084 367692 492086
rect 367756 492084 367762 492148
rect 204846 492010 204852 492012
rect 200438 491950 204852 492010
rect 146569 491947 146635 491950
rect 200205 491947 200271 491950
rect 204846 491948 204852 491950
rect 204916 491948 204922 492012
rect 232313 492010 232379 492013
rect 371734 492010 371740 492012
rect 232313 492008 371740 492010
rect 232313 491952 232318 492008
rect 232374 491952 371740 492008
rect 232313 491950 371740 491952
rect 232313 491947 232379 491950
rect 371734 491948 371740 491950
rect 371804 491948 371810 492012
rect 46606 491812 46612 491876
rect 46676 491874 46682 491876
rect 80789 491874 80855 491877
rect 46676 491872 80855 491874
rect 46676 491816 80794 491872
rect 80850 491816 80855 491872
rect 46676 491814 80855 491816
rect 46676 491812 46682 491814
rect 80789 491811 80855 491814
rect 145097 491874 145163 491877
rect 205030 491874 205036 491876
rect 145097 491872 205036 491874
rect 145097 491816 145102 491872
rect 145158 491816 205036 491872
rect 145097 491814 205036 491816
rect 145097 491811 145163 491814
rect 205030 491812 205036 491814
rect 205100 491812 205106 491876
rect 219198 491812 219204 491876
rect 219268 491874 219274 491876
rect 224861 491874 224927 491877
rect 219268 491872 224927 491874
rect 219268 491816 224866 491872
rect 224922 491816 224927 491872
rect 219268 491814 224927 491816
rect 219268 491812 219274 491814
rect 224861 491811 224927 491814
rect 234153 491874 234219 491877
rect 374494 491874 374500 491876
rect 234153 491872 374500 491874
rect 234153 491816 234158 491872
rect 234214 491816 374500 491872
rect 234153 491814 374500 491816
rect 234153 491811 234219 491814
rect 374494 491812 374500 491814
rect 374564 491812 374570 491876
rect 59118 491676 59124 491740
rect 59188 491738 59194 491740
rect 68645 491738 68711 491741
rect 59188 491736 68711 491738
rect 59188 491680 68650 491736
rect 68706 491680 68711 491736
rect 59188 491678 68711 491680
rect 59188 491676 59194 491678
rect 68645 491675 68711 491678
rect 187049 491738 187115 491741
rect 196750 491738 196756 491740
rect 187049 491736 196756 491738
rect 187049 491680 187054 491736
rect 187110 491680 196756 491736
rect 187049 491678 196756 491680
rect 187049 491675 187115 491678
rect 196750 491676 196756 491678
rect 196820 491676 196826 491740
rect 197629 491738 197695 491741
rect 198038 491738 198044 491740
rect 197629 491736 198044 491738
rect 197629 491680 197634 491736
rect 197690 491680 198044 491736
rect 197629 491678 198044 491680
rect 197629 491675 197695 491678
rect 198038 491676 198044 491678
rect 198108 491676 198114 491740
rect 200205 491738 200271 491741
rect 205214 491738 205220 491740
rect 200205 491736 205220 491738
rect 200205 491680 200210 491736
rect 200266 491680 205220 491736
rect 200205 491678 205220 491680
rect 200205 491675 200271 491678
rect 205214 491676 205220 491678
rect 205284 491676 205290 491740
rect 55070 491540 55076 491604
rect 55140 491602 55146 491604
rect 74257 491602 74323 491605
rect 55140 491600 74323 491602
rect 55140 491544 74262 491600
rect 74318 491544 74323 491600
rect 55140 491542 74323 491544
rect 55140 491540 55146 491542
rect 74257 491539 74323 491542
rect 197353 491602 197419 491605
rect 198406 491602 198412 491604
rect 197353 491600 198412 491602
rect 197353 491544 197358 491600
rect 197414 491544 198412 491600
rect 197353 491542 198412 491544
rect 197353 491539 197419 491542
rect 198406 491540 198412 491542
rect 198476 491540 198482 491604
rect 211153 491602 211219 491605
rect 211654 491602 211660 491604
rect 211153 491600 211660 491602
rect 211153 491544 211158 491600
rect 211214 491544 211660 491600
rect 211153 491542 211660 491544
rect 211153 491539 211219 491542
rect 211654 491540 211660 491542
rect 211724 491540 211730 491604
rect 191189 491466 191255 491469
rect 200614 491466 200620 491468
rect 191189 491464 200620 491466
rect 191189 491408 191194 491464
rect 191250 491408 200620 491464
rect 191189 491406 200620 491408
rect 191189 491403 191255 491406
rect 200614 491404 200620 491406
rect 200684 491404 200690 491468
rect 50286 491268 50292 491332
rect 50356 491330 50362 491332
rect 50521 491330 50587 491333
rect 52361 491332 52427 491333
rect 52310 491330 52316 491332
rect 50356 491328 50587 491330
rect 50356 491272 50526 491328
rect 50582 491272 50587 491328
rect 50356 491270 50587 491272
rect 52270 491270 52316 491330
rect 52380 491328 52427 491332
rect 52422 491272 52427 491328
rect 50356 491268 50362 491270
rect 50521 491267 50587 491270
rect 52310 491268 52316 491270
rect 52380 491268 52427 491272
rect 52361 491267 52427 491268
rect 197721 491330 197787 491333
rect 198590 491330 198596 491332
rect 197721 491328 198596 491330
rect 197721 491272 197726 491328
rect 197782 491272 198596 491328
rect 197721 491270 198596 491272
rect 197721 491267 197787 491270
rect 198590 491268 198596 491270
rect 198660 491268 198666 491332
rect 153745 490514 153811 490517
rect 213862 490514 213868 490516
rect 153745 490512 213868 490514
rect 153745 490456 153750 490512
rect 153806 490456 213868 490512
rect 153745 490454 213868 490456
rect 153745 490451 153811 490454
rect 213862 490452 213868 490454
rect 213932 490452 213938 490516
rect 57094 489636 57100 489700
rect 57164 489698 57170 489700
rect 120349 489698 120415 489701
rect 57164 489696 120415 489698
rect 57164 489640 120354 489696
rect 120410 489640 120415 489696
rect 57164 489638 120415 489640
rect 57164 489636 57170 489638
rect 120349 489635 120415 489638
rect 50521 489562 50587 489565
rect 115657 489562 115723 489565
rect 50521 489560 115723 489562
rect 50521 489504 50526 489560
rect 50582 489504 115662 489560
rect 115718 489504 115723 489560
rect 50521 489502 115723 489504
rect 50521 489499 50587 489502
rect 115657 489499 115723 489502
rect 50613 489426 50679 489429
rect 120257 489426 120323 489429
rect 50613 489424 120323 489426
rect 50613 489368 50618 489424
rect 50674 489368 120262 489424
rect 120318 489368 120323 489424
rect 50613 489366 120323 489368
rect 50613 489363 50679 489366
rect 120257 489363 120323 489366
rect 49049 489290 49115 489293
rect 120165 489290 120231 489293
rect 49049 489288 120231 489290
rect 49049 489232 49054 489288
rect 49110 489232 120170 489288
rect 120226 489232 120231 489288
rect 49049 489230 120231 489232
rect 49049 489227 49115 489230
rect 120165 489227 120231 489230
rect 46841 489154 46907 489157
rect 125777 489154 125843 489157
rect 46841 489152 125843 489154
rect 46841 489096 46846 489152
rect 46902 489096 125782 489152
rect 125838 489096 125843 489152
rect 46841 489094 125843 489096
rect 46841 489091 46907 489094
rect 125777 489091 125843 489094
rect 171409 489154 171475 489157
rect 206502 489154 206508 489156
rect 171409 489152 206508 489154
rect 171409 489096 171414 489152
rect 171470 489096 206508 489152
rect 171409 489094 206508 489096
rect 171409 489091 171475 489094
rect 206502 489092 206508 489094
rect 206572 489092 206578 489156
rect 129641 487794 129707 487797
rect 199142 487794 199148 487796
rect 129641 487792 199148 487794
rect 129641 487736 129646 487792
rect 129702 487736 199148 487792
rect 129641 487734 199148 487736
rect 129641 487731 129707 487734
rect 199142 487732 199148 487734
rect 199212 487732 199218 487796
rect 236545 487794 236611 487797
rect 378174 487794 378180 487796
rect 236545 487792 378180 487794
rect 236545 487736 236550 487792
rect 236606 487736 378180 487792
rect 236545 487734 378180 487736
rect 236545 487731 236611 487734
rect 378174 487732 378180 487734
rect 378244 487732 378250 487796
rect 47710 486916 47716 486980
rect 47780 486978 47786 486980
rect 121453 486978 121519 486981
rect 47780 486976 121519 486978
rect 47780 486920 121458 486976
rect 121514 486920 121519 486976
rect 47780 486918 121519 486920
rect 47780 486916 47786 486918
rect 121453 486915 121519 486918
rect 43713 486842 43779 486845
rect 121637 486842 121703 486845
rect 43713 486840 121703 486842
rect 43713 486784 43718 486840
rect 43774 486784 121642 486840
rect 121698 486784 121703 486840
rect 43713 486782 121703 486784
rect 43713 486779 43779 486782
rect 121637 486779 121703 486782
rect 43805 486706 43871 486709
rect 123017 486706 123083 486709
rect 43805 486704 123083 486706
rect 43805 486648 43810 486704
rect 43866 486648 123022 486704
rect 123078 486648 123083 486704
rect 43805 486646 123083 486648
rect 43805 486643 43871 486646
rect 123017 486643 123083 486646
rect 46749 486570 46815 486573
rect 127065 486570 127131 486573
rect 46749 486568 127131 486570
rect 46749 486512 46754 486568
rect 46810 486512 127070 486568
rect 127126 486512 127131 486568
rect 46749 486510 127131 486512
rect 46749 486507 46815 486510
rect 127065 486507 127131 486510
rect 147765 486570 147831 486573
rect 210366 486570 210372 486572
rect 147765 486568 210372 486570
rect 147765 486512 147770 486568
rect 147826 486512 210372 486568
rect 147765 486510 210372 486512
rect 147765 486507 147831 486510
rect 210366 486508 210372 486510
rect 210436 486508 210442 486572
rect 42333 486434 42399 486437
rect 127157 486434 127223 486437
rect 42333 486432 127223 486434
rect 42333 486376 42338 486432
rect 42394 486376 127162 486432
rect 127218 486376 127223 486432
rect 42333 486374 127223 486376
rect 42333 486371 42399 486374
rect 127157 486371 127223 486374
rect 143717 486434 143783 486437
rect 208894 486434 208900 486436
rect 143717 486432 208900 486434
rect 143717 486376 143722 486432
rect 143778 486376 208900 486432
rect 143717 486374 208900 486376
rect 143717 486371 143783 486374
rect 208894 486372 208900 486374
rect 208964 486372 208970 486436
rect -960 483836 480 484076
rect 47894 483924 47900 483988
rect 47964 483986 47970 483988
rect 122833 483986 122899 483989
rect 47964 483984 122899 483986
rect 47964 483928 122838 483984
rect 122894 483928 122899 483984
rect 47964 483926 122899 483928
rect 47964 483924 47970 483926
rect 122833 483923 122899 483926
rect 44950 483788 44956 483852
rect 45020 483850 45026 483852
rect 125685 483850 125751 483853
rect 45020 483848 125751 483850
rect 45020 483792 125690 483848
rect 125746 483792 125751 483848
rect 45020 483790 125751 483792
rect 45020 483788 45026 483790
rect 125685 483787 125751 483790
rect 44766 483652 44772 483716
rect 44836 483714 44842 483716
rect 126973 483714 127039 483717
rect 44836 483712 127039 483714
rect 44836 483656 126978 483712
rect 127034 483656 127039 483712
rect 44836 483654 127039 483656
rect 44836 483652 44842 483654
rect 126973 483651 127039 483654
rect 145005 483714 145071 483717
rect 206134 483714 206140 483716
rect 145005 483712 206140 483714
rect 145005 483656 145010 483712
rect 145066 483656 206140 483712
rect 145005 483654 206140 483656
rect 145005 483651 145071 483654
rect 206134 483652 206140 483654
rect 206204 483652 206210 483716
rect 229185 483714 229251 483717
rect 374678 483714 374684 483716
rect 229185 483712 374684 483714
rect 229185 483656 229190 483712
rect 229246 483656 374684 483712
rect 229185 483654 374684 483656
rect 229185 483651 229251 483654
rect 374678 483652 374684 483654
rect 374748 483652 374754 483716
rect 583520 479892 584960 480132
rect 150525 479498 150591 479501
rect 200798 479498 200804 479500
rect 150525 479496 200804 479498
rect 150525 479440 150530 479496
rect 150586 479440 200804 479496
rect 150525 479438 200804 479440
rect 150525 479435 150591 479438
rect 200798 479436 200804 479438
rect 200868 479436 200874 479500
rect 231945 479498 232011 479501
rect 378726 479498 378732 479500
rect 231945 479496 378732 479498
rect 231945 479440 231950 479496
rect 232006 479440 378732 479496
rect 231945 479438 378732 479440
rect 231945 479435 232011 479438
rect 378726 479436 378732 479438
rect 378796 479436 378802 479500
rect 179597 478274 179663 478277
rect 217174 478274 217180 478276
rect 179597 478272 217180 478274
rect 179597 478216 179602 478272
rect 179658 478216 217180 478272
rect 179597 478214 217180 478216
rect 179597 478211 179663 478214
rect 217174 478212 217180 478214
rect 217244 478212 217250 478276
rect 143533 478138 143599 478141
rect 206318 478138 206324 478140
rect 143533 478136 206324 478138
rect 143533 478080 143538 478136
rect 143594 478080 206324 478136
rect 143533 478078 206324 478080
rect 143533 478075 143599 478078
rect 206318 478076 206324 478078
rect 206388 478076 206394 478140
rect 231853 478138 231919 478141
rect 370446 478138 370452 478140
rect 231853 478136 370452 478138
rect 231853 478080 231858 478136
rect 231914 478080 370452 478136
rect 231853 478078 370452 478080
rect 231853 478075 231919 478078
rect 370446 478076 370452 478078
rect 370516 478076 370522 478140
rect 151813 476778 151879 476781
rect 208342 476778 208348 476780
rect 151813 476776 208348 476778
rect 151813 476720 151818 476776
rect 151874 476720 208348 476776
rect 151813 476718 208348 476720
rect 151813 476715 151879 476718
rect 208342 476716 208348 476718
rect 208412 476716 208418 476780
rect 292573 476778 292639 476781
rect 359774 476778 359780 476780
rect 292573 476776 359780 476778
rect 292573 476720 292578 476776
rect 292634 476720 359780 476776
rect 292573 476718 359780 476720
rect 292573 476715 292639 476718
rect 359774 476716 359780 476718
rect 359844 476716 359850 476780
rect 153193 475554 153259 475557
rect 219014 475554 219020 475556
rect 153193 475552 219020 475554
rect 153193 475496 153198 475552
rect 153254 475496 219020 475552
rect 153193 475494 219020 475496
rect 153193 475491 153259 475494
rect 219014 475492 219020 475494
rect 219084 475492 219090 475556
rect 146293 475418 146359 475421
rect 214414 475418 214420 475420
rect 146293 475416 214420 475418
rect 146293 475360 146298 475416
rect 146354 475360 214420 475416
rect 146293 475358 214420 475360
rect 146293 475355 146359 475358
rect 214414 475356 214420 475358
rect 214484 475356 214490 475420
rect 223573 475418 223639 475421
rect 375966 475418 375972 475420
rect 223573 475416 375972 475418
rect 223573 475360 223578 475416
rect 223634 475360 375972 475416
rect 223573 475358 375972 475360
rect 223573 475355 223639 475358
rect 375966 475356 375972 475358
rect 376036 475356 376042 475420
rect 157425 474058 157491 474061
rect 208526 474058 208532 474060
rect 157425 474056 208532 474058
rect 157425 474000 157430 474056
rect 157486 474000 208532 474056
rect 157425 473998 208532 474000
rect 157425 473995 157491 473998
rect 208526 473996 208532 473998
rect 208596 473996 208602 474060
rect 278957 474058 279023 474061
rect 377254 474058 377260 474060
rect 278957 474056 377260 474058
rect 278957 474000 278962 474056
rect 279018 474000 377260 474056
rect 278957 473998 377260 474000
rect 278957 473995 279023 473998
rect 377254 473996 377260 473998
rect 377324 473996 377330 474060
rect 144913 472562 144979 472565
rect 207974 472562 207980 472564
rect 144913 472560 207980 472562
rect 144913 472504 144918 472560
rect 144974 472504 207980 472560
rect 144913 472502 207980 472504
rect 144913 472499 144979 472502
rect 207974 472500 207980 472502
rect 208044 472500 208050 472564
rect 233325 472562 233391 472565
rect 376150 472562 376156 472564
rect 233325 472560 376156 472562
rect 233325 472504 233330 472560
rect 233386 472504 376156 472560
rect 233325 472502 376156 472504
rect 233325 472499 233391 472502
rect 376150 472500 376156 472502
rect 376220 472500 376226 472564
rect -960 471338 480 471428
rect 3509 471338 3575 471341
rect -960 471336 3575 471338
rect -960 471280 3514 471336
rect 3570 471280 3575 471336
rect -960 471278 3575 471280
rect -960 471188 480 471278
rect 3509 471275 3575 471278
rect 278865 471202 278931 471205
rect 359958 471202 359964 471204
rect 278865 471200 359964 471202
rect 278865 471144 278870 471200
rect 278926 471144 359964 471200
rect 278865 471142 359964 471144
rect 278865 471139 278931 471142
rect 359958 471140 359964 471142
rect 360028 471140 360034 471204
rect 164325 469978 164391 469981
rect 214598 469978 214604 469980
rect 164325 469976 214604 469978
rect 164325 469920 164330 469976
rect 164386 469920 214604 469976
rect 164325 469918 214604 469920
rect 164325 469915 164391 469918
rect 214598 469916 214604 469918
rect 214668 469916 214674 469980
rect 156045 469842 156111 469845
rect 215334 469842 215340 469844
rect 156045 469840 215340 469842
rect 156045 469784 156050 469840
rect 156106 469784 215340 469840
rect 156045 469782 215340 469784
rect 156045 469779 156111 469782
rect 215334 469780 215340 469782
rect 215404 469780 215410 469844
rect 155953 468482 156019 468485
rect 212574 468482 212580 468484
rect 155953 468480 212580 468482
rect 155953 468424 155958 468480
rect 156014 468424 212580 468480
rect 155953 468422 212580 468424
rect 155953 468419 156019 468422
rect 212574 468420 212580 468422
rect 212644 468420 212650 468484
rect 226425 467258 226491 467261
rect 363454 467258 363460 467260
rect 226425 467256 363460 467258
rect 226425 467200 226430 467256
rect 226486 467200 363460 467256
rect 226425 467198 363460 467200
rect 226425 467195 226491 467198
rect 363454 467196 363460 467198
rect 363524 467196 363530 467260
rect 172697 467122 172763 467125
rect 202270 467122 202276 467124
rect 172697 467120 202276 467122
rect 172697 467064 172702 467120
rect 172758 467064 202276 467120
rect 172697 467062 202276 467064
rect 172697 467059 172763 467062
rect 202270 467060 202276 467062
rect 202340 467060 202346 467124
rect 233233 467122 233299 467125
rect 378910 467122 378916 467124
rect 233233 467120 378916 467122
rect 233233 467064 233238 467120
rect 233294 467064 378916 467120
rect 233233 467062 378916 467064
rect 233233 467059 233299 467062
rect 378910 467060 378916 467062
rect 378980 467060 378986 467124
rect 580901 467122 580967 467125
rect 583520 467122 584960 467212
rect 580901 467120 584960 467122
rect 580901 467064 580906 467120
rect 580962 467064 584960 467120
rect 580901 467062 584960 467064
rect 580901 467059 580967 467062
rect 583520 466972 584960 467062
rect 53557 466306 53623 466309
rect 84377 466306 84443 466309
rect 53557 466304 84443 466306
rect 53557 466248 53562 466304
rect 53618 466248 84382 466304
rect 84438 466248 84443 466304
rect 53557 466246 84443 466248
rect 53557 466243 53623 466246
rect 84377 466243 84443 466246
rect 53649 466170 53715 466173
rect 85757 466170 85823 466173
rect 53649 466168 85823 466170
rect 53649 466112 53654 466168
rect 53710 466112 85762 466168
rect 85818 466112 85823 466168
rect 53649 466110 85823 466112
rect 53649 466107 53715 466110
rect 85757 466107 85823 466110
rect 52177 466034 52243 466037
rect 84285 466034 84351 466037
rect 52177 466032 84351 466034
rect 52177 465976 52182 466032
rect 52238 465976 84290 466032
rect 84346 465976 84351 466032
rect 52177 465974 84351 465976
rect 52177 465971 52243 465974
rect 84285 465971 84351 465974
rect 169845 466034 169911 466037
rect 207657 466034 207723 466037
rect 169845 466032 207723 466034
rect 169845 465976 169850 466032
rect 169906 465976 207662 466032
rect 207718 465976 207723 466032
rect 169845 465974 207723 465976
rect 169845 465971 169911 465974
rect 207657 465971 207723 465974
rect 59997 465898 60063 465901
rect 92657 465898 92723 465901
rect 59997 465896 92723 465898
rect 59997 465840 60002 465896
rect 60058 465840 92662 465896
rect 92718 465840 92723 465896
rect 59997 465838 92723 465840
rect 59997 465835 60063 465838
rect 92657 465835 92723 465838
rect 160277 465898 160343 465901
rect 204897 465898 204963 465901
rect 160277 465896 204963 465898
rect 160277 465840 160282 465896
rect 160338 465840 204902 465896
rect 204958 465840 204963 465896
rect 160277 465838 204963 465840
rect 160277 465835 160343 465838
rect 204897 465835 204963 465838
rect 48078 465700 48084 465764
rect 48148 465762 48154 465764
rect 81525 465762 81591 465765
rect 48148 465760 81591 465762
rect 48148 465704 81530 465760
rect 81586 465704 81591 465760
rect 48148 465702 81591 465704
rect 48148 465700 48154 465702
rect 81525 465699 81591 465702
rect 147673 465762 147739 465765
rect 218697 465762 218763 465765
rect 147673 465760 218763 465762
rect 147673 465704 147678 465760
rect 147734 465704 218702 465760
rect 218758 465704 218763 465760
rect 147673 465702 218763 465704
rect 147673 465699 147739 465702
rect 218697 465699 218763 465702
rect 265065 465762 265131 465765
rect 359406 465762 359412 465764
rect 265065 465760 359412 465762
rect 265065 465704 265070 465760
rect 265126 465704 359412 465760
rect 265065 465702 359412 465704
rect 265065 465699 265131 465702
rect 359406 465700 359412 465702
rect 359476 465700 359482 465764
rect 58934 463388 58940 463452
rect 59004 463450 59010 463452
rect 69197 463450 69263 463453
rect 59004 463448 69263 463450
rect 59004 463392 69202 463448
rect 69258 463392 69263 463448
rect 59004 463390 69263 463392
rect 59004 463388 59010 463390
rect 69197 463387 69263 463390
rect 183645 463450 183711 463453
rect 199326 463450 199332 463452
rect 183645 463448 199332 463450
rect 183645 463392 183650 463448
rect 183706 463392 199332 463448
rect 183645 463390 199332 463392
rect 183645 463387 183711 463390
rect 199326 463388 199332 463390
rect 199396 463388 199402 463452
rect 46422 463252 46428 463316
rect 46492 463314 46498 463316
rect 70485 463314 70551 463317
rect 46492 463312 70551 463314
rect 46492 463256 70490 463312
rect 70546 463256 70551 463312
rect 46492 463254 70551 463256
rect 46492 463252 46498 463254
rect 70485 463251 70551 463254
rect 169753 463314 169819 463317
rect 209221 463314 209287 463317
rect 169753 463312 209287 463314
rect 169753 463256 169758 463312
rect 169814 463256 209226 463312
rect 209282 463256 209287 463312
rect 169753 463254 209287 463256
rect 169753 463251 169819 463254
rect 209221 463251 209287 463254
rect 53414 463116 53420 463180
rect 53484 463178 53490 463180
rect 80145 463178 80211 463181
rect 53484 463176 80211 463178
rect 53484 463120 80150 463176
rect 80206 463120 80211 463176
rect 53484 463118 80211 463120
rect 53484 463116 53490 463118
rect 80145 463115 80211 463118
rect 158713 463178 158779 463181
rect 202086 463178 202092 463180
rect 158713 463176 202092 463178
rect 158713 463120 158718 463176
rect 158774 463120 202092 463176
rect 158713 463118 202092 463120
rect 158713 463115 158779 463118
rect 202086 463116 202092 463118
rect 202156 463116 202162 463180
rect 49417 463042 49483 463045
rect 93853 463042 93919 463045
rect 49417 463040 93919 463042
rect 49417 462984 49422 463040
rect 49478 462984 93858 463040
rect 93914 462984 93919 463040
rect 49417 462982 93919 462984
rect 49417 462979 49483 462982
rect 93853 462979 93919 462982
rect 169937 463042 170003 463045
rect 216070 463042 216076 463044
rect 169937 463040 216076 463042
rect 169937 462984 169942 463040
rect 169998 462984 216076 463040
rect 169937 462982 216076 462984
rect 169937 462979 170003 462982
rect 216070 462980 216076 462982
rect 216140 462980 216146 463044
rect 296713 463042 296779 463045
rect 376702 463042 376708 463044
rect 296713 463040 376708 463042
rect 296713 462984 296718 463040
rect 296774 462984 376708 463040
rect 296713 462982 376708 462984
rect 296713 462979 296779 462982
rect 376702 462980 376708 462982
rect 376772 462980 376778 463044
rect 49325 462906 49391 462909
rect 93945 462906 94011 462909
rect 49325 462904 94011 462906
rect 49325 462848 49330 462904
rect 49386 462848 93950 462904
rect 94006 462848 94011 462904
rect 49325 462846 94011 462848
rect 49325 462843 49391 462846
rect 93945 462843 94011 462846
rect 107653 462906 107719 462909
rect 198774 462906 198780 462908
rect 107653 462904 198780 462906
rect 107653 462848 107658 462904
rect 107714 462848 198780 462904
rect 107653 462846 198780 462848
rect 107653 462843 107719 462846
rect 198774 462844 198780 462846
rect 198844 462844 198850 462908
rect 258165 462906 258231 462909
rect 359590 462906 359596 462908
rect 258165 462904 359596 462906
rect 258165 462848 258170 462904
rect 258226 462848 359596 462904
rect 258165 462846 359596 462848
rect 258165 462843 258231 462846
rect 359590 462844 359596 462846
rect 359660 462844 359666 462908
rect 179638 462164 179644 462228
rect 179708 462226 179714 462228
rect 180057 462226 180123 462229
rect 179708 462224 180123 462226
rect 179708 462168 180062 462224
rect 180118 462168 180123 462224
rect 179708 462166 180123 462168
rect 179708 462164 179714 462166
rect 180057 462163 180123 462166
rect 510838 462164 510844 462228
rect 510908 462226 510914 462228
rect 511257 462226 511323 462229
rect 510908 462224 511323 462226
rect 510908 462168 511262 462224
rect 511318 462168 511323 462224
rect 510908 462166 511323 462168
rect 510908 462164 510914 462166
rect 511257 462163 511323 462166
rect 171317 461682 171383 461685
rect 202454 461682 202460 461684
rect 171317 461680 202460 461682
rect 171317 461624 171322 461680
rect 171378 461624 202460 461680
rect 171317 461622 202460 461624
rect 171317 461619 171383 461622
rect 202454 461620 202460 461622
rect 202524 461620 202530 461684
rect 60222 461484 60228 461548
rect 60292 461546 60298 461548
rect 73153 461546 73219 461549
rect 60292 461544 73219 461546
rect 60292 461488 73158 461544
rect 73214 461488 73219 461544
rect 60292 461486 73219 461488
rect 60292 461484 60298 461486
rect 73153 461483 73219 461486
rect 161565 461546 161631 461549
rect 203190 461546 203196 461548
rect 161565 461544 203196 461546
rect 161565 461488 161570 461544
rect 161626 461488 203196 461544
rect 161565 461486 203196 461488
rect 161565 461483 161631 461486
rect 203190 461484 203196 461486
rect 203260 461484 203266 461548
rect 178309 461412 178375 461413
rect 178309 461408 178356 461412
rect 178420 461410 178426 461412
rect 178309 461352 178314 461408
rect 178309 461348 178356 461352
rect 178420 461350 178466 461410
rect 178420 461348 178426 461350
rect 198958 461348 198964 461412
rect 199028 461410 199034 461412
rect 199561 461410 199627 461413
rect 199028 461408 199627 461410
rect 199028 461352 199566 461408
rect 199622 461352 199627 461408
rect 199028 461350 199627 461352
rect 199028 461348 199034 461350
rect 178309 461347 178375 461348
rect 199561 461347 199627 461350
rect 339677 461276 339743 461277
rect 339677 461272 339724 461276
rect 339788 461274 339794 461276
rect 339677 461216 339682 461272
rect 339677 461212 339724 461216
rect 339788 461214 339834 461274
rect 339788 461212 339794 461214
rect 339677 461211 339743 461212
rect 190913 461004 190979 461005
rect 338297 461004 338363 461005
rect 350993 461004 351059 461005
rect 190862 461002 190868 461004
rect 190822 460942 190868 461002
rect 190932 461000 190979 461004
rect 338246 461002 338252 461004
rect 190974 460944 190979 461000
rect 190862 460940 190868 460942
rect 190932 460940 190979 460944
rect 338206 460942 338252 461002
rect 338316 461000 338363 461004
rect 350942 461002 350948 461004
rect 338358 460944 338363 461000
rect 338246 460940 338252 460942
rect 338316 460940 338363 460944
rect 350902 460942 350948 461002
rect 351012 461000 351059 461004
rect 351054 460944 351059 461000
rect 350942 460940 350948 460942
rect 351012 460940 351059 460944
rect 190913 460939 190979 460940
rect 338297 460939 338363 460940
rect 350993 460939 351059 460940
rect 498469 461004 498535 461005
rect 499849 461004 499915 461005
rect 498469 461000 498516 461004
rect 498580 461002 498586 461004
rect 499798 461002 499804 461004
rect 498469 460944 498474 461000
rect 498469 460940 498516 460944
rect 498580 460942 498626 461002
rect 499758 460942 499804 461002
rect 499868 461000 499915 461004
rect 499910 460944 499915 461000
rect 498580 460940 498586 460942
rect 499798 460940 499804 460942
rect 499868 460940 499915 460944
rect 498469 460939 498535 460940
rect 499849 460939 499915 460940
rect 58750 460804 58756 460868
rect 58820 460866 58826 460868
rect 69013 460866 69079 460869
rect 58820 460864 69079 460866
rect 58820 460808 69018 460864
rect 69074 460808 69079 460864
rect 58820 460806 69079 460808
rect 58820 460804 58826 460806
rect 69013 460803 69079 460806
rect 54886 460668 54892 460732
rect 54956 460730 54962 460732
rect 71773 460730 71839 460733
rect 54956 460728 71839 460730
rect 54956 460672 71778 460728
rect 71834 460672 71839 460728
rect 54956 460670 71839 460672
rect 54956 460668 54962 460670
rect 71773 460667 71839 460670
rect 50470 460532 50476 460596
rect 50540 460594 50546 460596
rect 69105 460594 69171 460597
rect 50540 460592 69171 460594
rect 50540 460536 69110 460592
rect 69166 460536 69171 460592
rect 50540 460534 69171 460536
rect 50540 460532 50546 460534
rect 69105 460531 69171 460534
rect 55622 460396 55628 460460
rect 55692 460458 55698 460460
rect 74625 460458 74691 460461
rect 55692 460456 74691 460458
rect 55692 460400 74630 460456
rect 74686 460400 74691 460456
rect 55692 460398 74691 460400
rect 55692 460396 55698 460398
rect 74625 460395 74691 460398
rect 166993 460458 167059 460461
rect 203006 460458 203012 460460
rect 166993 460456 203012 460458
rect 166993 460400 166998 460456
rect 167054 460400 203012 460456
rect 166993 460398 203012 460400
rect 166993 460395 167059 460398
rect 203006 460396 203012 460398
rect 203076 460396 203082 460460
rect 54702 460260 54708 460324
rect 54772 460322 54778 460324
rect 76005 460322 76071 460325
rect 54772 460320 76071 460322
rect 54772 460264 76010 460320
rect 76066 460264 76071 460320
rect 54772 460262 76071 460264
rect 54772 460260 54778 460262
rect 76005 460259 76071 460262
rect 154573 460322 154639 460325
rect 209814 460322 209820 460324
rect 154573 460320 209820 460322
rect 154573 460264 154578 460320
rect 154634 460264 209820 460320
rect 154573 460262 209820 460264
rect 154573 460259 154639 460262
rect 209814 460260 209820 460262
rect 209884 460260 209890 460324
rect 52126 460124 52132 460188
rect 52196 460186 52202 460188
rect 74717 460186 74783 460189
rect 52196 460184 74783 460186
rect 52196 460128 74722 460184
rect 74778 460128 74783 460184
rect 52196 460126 74783 460128
rect 52196 460124 52202 460126
rect 74717 460123 74783 460126
rect 157333 460186 157399 460189
rect 218646 460186 218652 460188
rect 157333 460184 218652 460186
rect 157333 460128 157338 460184
rect 157394 460128 218652 460184
rect 157333 460126 218652 460128
rect 157333 460123 157399 460126
rect 218646 460124 218652 460126
rect 218716 460124 218722 460188
rect 298093 460186 298159 460189
rect 376886 460186 376892 460188
rect 298093 460184 376892 460186
rect 298093 460128 298098 460184
rect 298154 460128 376892 460184
rect 298093 460126 376892 460128
rect 298093 460123 298159 460126
rect 376886 460124 376892 460126
rect 376956 460124 376962 460188
rect 58566 459988 58572 460052
rect 58636 460050 58642 460052
rect 67725 460050 67791 460053
rect 58636 460048 67791 460050
rect 58636 459992 67730 460048
rect 67786 459992 67791 460048
rect 58636 459990 67791 459992
rect 58636 459988 58642 459990
rect 67725 459987 67791 459990
rect 48630 459580 48636 459644
rect 48700 459642 48706 459644
rect 49233 459642 49299 459645
rect 48700 459640 49299 459642
rect 48700 459584 49238 459640
rect 49294 459584 49299 459640
rect 48700 459582 49299 459584
rect 48700 459580 48706 459582
rect 49233 459579 49299 459582
rect 50654 459580 50660 459644
rect 50724 459642 50730 459644
rect 50981 459642 51047 459645
rect 50724 459640 51047 459642
rect 50724 459584 50986 459640
rect 51042 459584 51047 459640
rect 50724 459582 51047 459584
rect 50724 459580 50730 459582
rect 50981 459579 51047 459582
rect 51758 459580 51764 459644
rect 51828 459642 51834 459644
rect 52269 459642 52335 459645
rect 51828 459640 52335 459642
rect 51828 459584 52274 459640
rect 52330 459584 52335 459640
rect 51828 459582 52335 459584
rect 51828 459580 51834 459582
rect 52269 459579 52335 459582
rect 53230 459580 53236 459644
rect 53300 459642 53306 459644
rect 53465 459642 53531 459645
rect 55489 459644 55555 459645
rect 55438 459642 55444 459644
rect 53300 459640 53531 459642
rect 53300 459584 53470 459640
rect 53526 459584 53531 459640
rect 53300 459582 53531 459584
rect 55398 459582 55444 459642
rect 55508 459640 55555 459644
rect 55550 459584 55555 459640
rect 53300 459580 53306 459582
rect 53465 459579 53531 459582
rect 55438 459580 55444 459582
rect 55508 459580 55555 459584
rect 216990 459580 216996 459644
rect 217060 459642 217066 459644
rect 220997 459642 221063 459645
rect 217060 459640 221063 459642
rect 217060 459584 221002 459640
rect 221058 459584 221063 459640
rect 217060 459582 221063 459584
rect 217060 459580 217066 459582
rect 55489 459579 55555 459580
rect 220997 459579 221063 459582
rect 186313 459506 186379 459509
rect 213453 459506 213519 459509
rect 186313 459504 213519 459506
rect 186313 459448 186318 459504
rect 186374 459448 213458 459504
rect 213514 459448 213519 459504
rect 186313 459446 213519 459448
rect 186313 459443 186379 459446
rect 213453 459443 213519 459446
rect 172513 459370 172579 459373
rect 205398 459370 205404 459372
rect 172513 459368 205404 459370
rect 172513 459312 172518 459368
rect 172574 459312 205404 459368
rect 172513 459310 205404 459312
rect 172513 459307 172579 459310
rect 205398 459308 205404 459310
rect 205468 459308 205474 459372
rect 171133 459234 171199 459237
rect 208158 459234 208164 459236
rect 171133 459232 208164 459234
rect 171133 459176 171138 459232
rect 171194 459176 208164 459232
rect 171133 459174 208164 459176
rect 171133 459171 171199 459174
rect 208158 459172 208164 459174
rect 208228 459172 208234 459236
rect 57462 459036 57468 459100
rect 57532 459098 57538 459100
rect 80053 459098 80119 459101
rect 57532 459096 80119 459098
rect 57532 459040 80058 459096
rect 80114 459040 80119 459096
rect 57532 459038 80119 459040
rect 57532 459036 57538 459038
rect 80053 459035 80119 459038
rect 161473 459098 161539 459101
rect 206461 459098 206527 459101
rect 161473 459096 206527 459098
rect 161473 459040 161478 459096
rect 161534 459040 206466 459096
rect 206522 459040 206527 459096
rect 161473 459038 206527 459040
rect 161473 459035 161539 459038
rect 206461 459035 206527 459038
rect -960 458826 480 458916
rect 57830 458900 57836 458964
rect 57900 458962 57906 458964
rect 89897 458962 89963 458965
rect 57900 458960 89963 458962
rect 57900 458904 89902 458960
rect 89958 458904 89963 458960
rect 57900 458902 89963 458904
rect 57900 458900 57906 458902
rect 89897 458899 89963 458902
rect 162853 458962 162919 458965
rect 213126 458962 213132 458964
rect 162853 458960 213132 458962
rect 162853 458904 162858 458960
rect 162914 458904 213132 458960
rect 162853 458902 213132 458904
rect 162853 458899 162919 458902
rect 213126 458900 213132 458902
rect 213196 458900 213202 458964
rect 2773 458826 2839 458829
rect -960 458824 2839 458826
rect -960 458768 2778 458824
rect 2834 458768 2839 458824
rect -960 458766 2839 458768
rect -960 458676 480 458766
rect 2773 458763 2839 458766
rect 57646 458764 57652 458828
rect 57716 458826 57722 458828
rect 91277 458826 91343 458829
rect 57716 458824 91343 458826
rect 57716 458768 91282 458824
rect 91338 458768 91343 458824
rect 57716 458766 91343 458768
rect 57716 458764 57722 458766
rect 91277 458763 91343 458766
rect 150433 458826 150499 458829
rect 215886 458826 215892 458828
rect 150433 458824 215892 458826
rect 150433 458768 150438 458824
rect 150494 458768 215892 458824
rect 150433 458766 215892 458768
rect 150433 458763 150499 458766
rect 215886 458764 215892 458766
rect 215956 458764 215962 458828
rect 199009 454746 199075 454749
rect 358813 454746 358879 454749
rect 516593 454746 516659 454749
rect 196558 454744 199075 454746
rect 196558 454688 199014 454744
rect 199070 454688 199075 454744
rect 196558 454686 199075 454688
rect 196558 454190 196618 454686
rect 199009 454683 199075 454686
rect 356562 454744 358879 454746
rect 356562 454688 358818 454744
rect 358874 454688 358879 454744
rect 356562 454686 358879 454688
rect 356562 454190 356622 454686
rect 358813 454683 358879 454686
rect 516558 454744 516659 454746
rect 516558 454688 516598 454744
rect 516654 454688 516659 454744
rect 516558 454683 516659 454688
rect 516558 454202 516618 454683
rect 518893 454202 518959 454205
rect 516558 454200 518959 454202
rect 516558 454144 518898 454200
rect 518954 454144 518959 454200
rect 583520 454188 584960 454428
rect 516558 454142 518959 454144
rect 518893 454139 518959 454142
rect -960 446164 480 446404
rect 579889 441554 579955 441557
rect 583520 441554 584960 441644
rect 579889 441552 584960 441554
rect 579889 441496 579894 441552
rect 579950 441496 584960 441552
rect 579889 441494 584960 441496
rect 579889 441491 579955 441494
rect 583520 441404 584960 441494
rect -960 433516 480 433756
rect 583520 428620 584960 428860
rect -960 421154 480 421244
rect 3141 421154 3207 421157
rect -960 421152 3207 421154
rect -960 421096 3146 421152
rect 3202 421096 3207 421152
rect -960 421094 3207 421096
rect -960 421004 480 421094
rect 3141 421091 3207 421094
rect 580901 415986 580967 415989
rect 583520 415986 584960 416076
rect 580901 415984 584960 415986
rect 580901 415928 580906 415984
rect 580962 415928 584960 415984
rect 580901 415926 584960 415928
rect 580901 415923 580967 415926
rect 583520 415836 584960 415926
rect 57237 412450 57303 412453
rect 57237 412448 60062 412450
rect 57237 412392 57242 412448
rect 57298 412392 60062 412448
rect 57237 412390 60062 412392
rect 57237 412387 57303 412390
rect 60002 411894 60062 412390
rect 217869 411906 217935 411909
rect 219390 411906 220064 411924
rect 217869 411904 220064 411906
rect 217869 411848 217874 411904
rect 217930 411864 220064 411904
rect 377581 411906 377647 411909
rect 379470 411906 380052 411924
rect 377581 411904 380052 411906
rect 217930 411848 219450 411864
rect 217869 411846 219450 411848
rect 377581 411848 377586 411904
rect 377642 411864 380052 411904
rect 377642 411848 379530 411864
rect 377581 411846 379530 411848
rect 217869 411843 217935 411846
rect 377581 411843 377647 411846
rect 57237 411226 57303 411229
rect 57237 411224 60062 411226
rect 57237 411168 57242 411224
rect 57298 411168 60062 411224
rect 57237 411166 60062 411168
rect 57237 411163 57303 411166
rect 60002 410942 60062 411166
rect 216765 410954 216831 410957
rect 217685 410954 217751 410957
rect 219390 410954 220064 410972
rect 216765 410952 220064 410954
rect 216765 410896 216770 410952
rect 216826 410896 217690 410952
rect 217746 410912 220064 410952
rect 377765 410954 377831 410957
rect 379470 410954 380052 410972
rect 377765 410952 380052 410954
rect 217746 410896 219450 410912
rect 216765 410894 219450 410896
rect 377765 410896 377770 410952
rect 377826 410912 380052 410952
rect 377826 410896 379530 410912
rect 377765 410894 379530 410896
rect 216765 410891 216831 410894
rect 217685 410891 217751 410894
rect 377765 410891 377831 410894
rect 377305 410002 377371 410005
rect 377765 410002 377831 410005
rect 377305 410000 377831 410002
rect 377305 409944 377310 410000
rect 377366 409944 377770 410000
rect 377826 409944 377831 410000
rect 377305 409942 377831 409944
rect 377305 409939 377371 409942
rect 377765 409939 377831 409942
rect 216765 408778 216831 408781
rect 219390 408778 220064 408796
rect 216765 408776 220064 408778
rect 57237 408642 57303 408645
rect 60002 408642 60062 408766
rect 216765 408720 216770 408776
rect 216826 408736 220064 408776
rect 377857 408778 377923 408781
rect 379470 408778 380052 408796
rect 377857 408776 380052 408778
rect 216826 408720 219450 408736
rect 216765 408718 219450 408720
rect 377857 408720 377862 408776
rect 377918 408736 380052 408776
rect 377918 408720 379530 408736
rect 377857 408718 379530 408720
rect 216765 408715 216831 408718
rect 377857 408715 377923 408718
rect 57237 408640 60062 408642
rect -960 408506 480 408596
rect 57237 408584 57242 408640
rect 57298 408584 60062 408640
rect 57237 408582 60062 408584
rect 57237 408579 57303 408582
rect 2773 408506 2839 408509
rect -960 408504 2839 408506
rect -960 408448 2778 408504
rect 2834 408448 2839 408504
rect -960 408446 2839 408448
rect -960 408356 480 408446
rect 2773 408443 2839 408446
rect 217225 407826 217291 407829
rect 217961 407826 218027 407829
rect 219390 407826 220064 407844
rect 217225 407824 220064 407826
rect 57237 407282 57303 407285
rect 60002 407282 60062 407814
rect 217225 407768 217230 407824
rect 217286 407768 217966 407824
rect 218022 407784 220064 407824
rect 377029 407826 377095 407829
rect 377397 407826 377463 407829
rect 379470 407826 380052 407844
rect 377029 407824 380052 407826
rect 218022 407768 219450 407784
rect 217225 407766 219450 407768
rect 377029 407768 377034 407824
rect 377090 407768 377402 407824
rect 377458 407784 380052 407824
rect 377458 407768 379530 407784
rect 377029 407766 379530 407768
rect 217225 407763 217291 407766
rect 217961 407763 218027 407766
rect 377029 407763 377095 407766
rect 377397 407763 377463 407766
rect 57237 407280 60062 407282
rect 57237 407224 57242 407280
rect 57298 407224 60062 407280
rect 57237 407222 60062 407224
rect 57237 407219 57303 407222
rect 217593 406058 217659 406061
rect 219390 406058 220064 406076
rect 217593 406056 220064 406058
rect 57237 405786 57303 405789
rect 60002 405786 60062 406046
rect 217593 406000 217598 406056
rect 217654 406016 220064 406056
rect 377397 406058 377463 406061
rect 377949 406058 378015 406061
rect 379470 406058 380052 406076
rect 377397 406056 380052 406058
rect 217654 406000 219450 406016
rect 217593 405998 219450 406000
rect 377397 406000 377402 406056
rect 377458 406000 377954 406056
rect 378010 406016 380052 406056
rect 378010 406000 379530 406016
rect 377397 405998 379530 406000
rect 217593 405995 217659 405998
rect 377397 405995 377463 405998
rect 377949 405995 378015 405998
rect 57237 405784 60062 405786
rect 57237 405728 57242 405784
rect 57298 405728 60062 405784
rect 57237 405726 60062 405728
rect 57237 405723 57303 405726
rect 216857 404970 216923 404973
rect 219390 404970 220064 404988
rect 216857 404968 220064 404970
rect 57237 404426 57303 404429
rect 60002 404426 60062 404958
rect 216857 404912 216862 404968
rect 216918 404928 220064 404968
rect 377673 404970 377739 404973
rect 379470 404970 380052 404988
rect 377673 404968 380052 404970
rect 216918 404912 219450 404928
rect 216857 404910 219450 404912
rect 377673 404912 377678 404968
rect 377734 404928 380052 404968
rect 377734 404912 379530 404928
rect 377673 404910 379530 404912
rect 216857 404907 216923 404910
rect 377673 404907 377739 404910
rect 57237 404424 60062 404426
rect 57237 404368 57242 404424
rect 57298 404368 60062 404424
rect 57237 404366 60062 404368
rect 57237 404363 57303 404366
rect 217317 404290 217383 404293
rect 217961 404290 218027 404293
rect 217317 404288 218027 404290
rect 217317 404232 217322 404288
rect 217378 404232 217966 404288
rect 218022 404232 218027 404288
rect 217317 404230 218027 404232
rect 217317 404227 217383 404230
rect 217961 404227 218027 404230
rect 217961 403202 218027 403205
rect 219390 403202 220064 403220
rect 217961 403200 220064 403202
rect 57237 403066 57303 403069
rect 60002 403066 60062 403190
rect 217961 403144 217966 403200
rect 218022 403160 220064 403200
rect 377765 403202 377831 403205
rect 379470 403202 380052 403220
rect 377765 403200 380052 403202
rect 218022 403144 219450 403160
rect 217961 403142 219450 403144
rect 377765 403144 377770 403200
rect 377826 403160 380052 403200
rect 377826 403144 379530 403160
rect 377765 403142 379530 403144
rect 217961 403139 218027 403142
rect 377765 403139 377831 403142
rect 57237 403064 60062 403066
rect 57237 403008 57242 403064
rect 57298 403008 60062 403064
rect 583520 403052 584960 403292
rect 57237 403006 60062 403008
rect 57237 403003 57303 403006
rect -960 395844 480 396084
rect 199193 394634 199259 394637
rect 199745 394634 199811 394637
rect 196558 394632 199811 394634
rect 196558 394576 199198 394632
rect 199254 394576 199750 394632
rect 199806 394576 199811 394632
rect 196558 394574 199811 394576
rect 196558 394350 196618 394574
rect 199193 394571 199259 394574
rect 199745 394571 199811 394574
rect 356562 393818 356622 394350
rect 358905 393818 358971 393821
rect 356562 393816 358971 393818
rect 356562 393760 358910 393816
rect 358966 393760 358971 393816
rect 356562 393758 358971 393760
rect 516558 393818 516618 394350
rect 519169 393818 519235 393821
rect 516558 393816 519235 393818
rect 516558 393760 519174 393816
rect 519230 393760 519235 393816
rect 516558 393758 519235 393760
rect 358905 393755 358971 393758
rect 519169 393755 519235 393758
rect 199561 392730 199627 392733
rect 196558 392728 199627 392730
rect 196558 392672 199566 392728
rect 199622 392672 199627 392728
rect 196558 392670 199627 392672
rect 199561 392667 199627 392670
rect 356562 392186 356622 392718
rect 359917 392186 359983 392189
rect 356562 392184 359983 392186
rect 356562 392128 359922 392184
rect 359978 392128 359983 392184
rect 356562 392126 359983 392128
rect 516558 392186 516618 392718
rect 519353 392186 519419 392189
rect 516558 392184 519419 392186
rect 516558 392128 519358 392184
rect 519414 392128 519419 392184
rect 516558 392126 519419 392128
rect 359917 392123 359983 392126
rect 519353 392123 519419 392126
rect 199377 391370 199443 391373
rect 196558 391368 199443 391370
rect 196558 391312 199382 391368
rect 199438 391312 199443 391368
rect 196558 391310 199443 391312
rect 199377 391307 199443 391310
rect 356562 390826 356622 391358
rect 358997 390826 359063 390829
rect 356562 390824 359063 390826
rect 356562 390768 359002 390824
rect 359058 390768 359063 390824
rect 356562 390766 359063 390768
rect 516558 390826 516618 391358
rect 518985 390826 519051 390829
rect 516558 390824 519051 390826
rect 516558 390768 518990 390824
rect 519046 390768 519051 390824
rect 516558 390766 519051 390768
rect 358997 390763 359063 390766
rect 518985 390763 519051 390766
rect 578877 390418 578943 390421
rect 583520 390418 584960 390508
rect 578877 390416 584960 390418
rect 578877 390360 578882 390416
rect 578938 390360 584960 390416
rect 578877 390358 584960 390360
rect 578877 390355 578943 390358
rect 583520 390268 584960 390358
rect 199469 389874 199535 389877
rect 196558 389872 199535 389874
rect 196558 389816 199474 389872
rect 199530 389816 199535 389872
rect 196558 389814 199535 389816
rect 199469 389811 199535 389814
rect 356562 389330 356622 389862
rect 359825 389330 359891 389333
rect 356562 389328 359891 389330
rect 356562 389272 359830 389328
rect 359886 389272 359891 389328
rect 356562 389270 359891 389272
rect 516558 389330 516618 389862
rect 519077 389330 519143 389333
rect 516558 389328 519143 389330
rect 516558 389272 519082 389328
rect 519138 389272 519143 389328
rect 516558 389270 519143 389272
rect 359825 389267 359891 389270
rect 519077 389267 519143 389270
rect 199469 389194 199535 389197
rect 199653 389194 199719 389197
rect 199469 389192 199719 389194
rect 199469 389136 199474 389192
rect 199530 389136 199658 389192
rect 199714 389136 199719 389192
rect 199469 389134 199719 389136
rect 199469 389131 199535 389134
rect 199653 389131 199719 389134
rect 196558 388514 196618 388638
rect 199142 388514 199148 388516
rect 196558 388454 199148 388514
rect 199142 388452 199148 388454
rect 199212 388514 199218 388516
rect 199510 388514 199516 388516
rect 199212 388454 199516 388514
rect 199212 388452 199218 388454
rect 199510 388452 199516 388454
rect 199580 388452 199586 388516
rect 356562 388106 356622 388638
rect 359089 388106 359155 388109
rect 356562 388104 359155 388106
rect 356562 388048 359094 388104
rect 359150 388048 359155 388104
rect 356562 388046 359155 388048
rect 516558 388106 516618 388638
rect 519261 388106 519327 388109
rect 516558 388104 519327 388106
rect 516558 388048 519266 388104
rect 519322 388048 519327 388104
rect 516558 388046 519327 388048
rect 359089 388043 359155 388046
rect 519261 388043 519327 388046
rect 57237 384978 57303 384981
rect 216673 384978 216739 384981
rect 219390 384978 220064 384996
rect 57237 384976 60062 384978
rect 57237 384920 57242 384976
rect 57298 384920 60062 384976
rect 57237 384918 60062 384920
rect 216673 384976 220064 384978
rect 216673 384920 216678 384976
rect 216734 384936 220064 384976
rect 376937 384978 377003 384981
rect 379470 384978 380052 384996
rect 376937 384976 380052 384978
rect 216734 384920 219450 384936
rect 216673 384918 219450 384920
rect 376937 384920 376942 384976
rect 376998 384936 380052 384976
rect 376998 384920 379530 384936
rect 376937 384918 379530 384920
rect 57237 384915 57303 384918
rect 216673 384915 216739 384918
rect 376937 384915 377003 384918
rect -960 383196 480 383436
rect 57513 383346 57579 383349
rect 59494 383346 60032 383364
rect 57513 383344 60032 383346
rect 57513 383288 57518 383344
rect 57574 383304 60032 383344
rect 216673 383346 216739 383349
rect 219390 383346 220064 383364
rect 216673 383344 220064 383346
rect 57574 383288 59554 383304
rect 57513 383286 59554 383288
rect 216673 383288 216678 383344
rect 216734 383304 220064 383344
rect 376937 383346 377003 383349
rect 379470 383346 380052 383364
rect 376937 383344 380052 383346
rect 216734 383288 219450 383304
rect 216673 383286 219450 383288
rect 376937 383288 376942 383344
rect 376998 383304 380052 383344
rect 376998 383288 379530 383304
rect 376937 383286 379530 383288
rect 57513 383283 57579 383286
rect 216673 383283 216739 383286
rect 376937 383283 377003 383286
rect 56869 383074 56935 383077
rect 217041 383074 217107 383077
rect 219390 383074 220064 383092
rect 56869 383072 60062 383074
rect 56869 383016 56874 383072
rect 56930 383016 60062 383072
rect 56869 383014 60062 383016
rect 217041 383072 220064 383074
rect 217041 383016 217046 383072
rect 217102 383032 220064 383072
rect 376845 383074 376911 383077
rect 379470 383074 380052 383092
rect 376845 383072 380052 383074
rect 217102 383016 219450 383032
rect 217041 383014 219450 383016
rect 376845 383016 376850 383072
rect 376906 383032 380052 383072
rect 376906 383016 379530 383032
rect 376845 383014 379530 383016
rect 56869 383011 56935 383014
rect 217041 383011 217107 383014
rect 376845 383011 376911 383014
rect 48630 380972 48636 381036
rect 48700 381034 48706 381036
rect 49601 381034 49667 381037
rect 48700 381032 49667 381034
rect 48700 380976 49606 381032
rect 49662 380976 49667 381032
rect 48700 380974 49667 380976
rect 48700 380972 48706 380974
rect 49601 380971 49667 380974
rect 583520 377484 584960 377724
rect 50286 375260 50292 375324
rect 50356 375322 50362 375324
rect 50981 375322 51047 375325
rect 50356 375320 51047 375322
rect 50356 375264 50986 375320
rect 51042 375264 51047 375320
rect 50356 375262 51047 375264
rect 50356 375260 50362 375262
rect 50981 375259 51047 375262
rect 198038 375260 198044 375324
rect 198108 375322 198114 375324
rect 198641 375322 198707 375325
rect 198108 375320 198707 375322
rect 198108 375264 198646 375320
rect 198702 375264 198707 375320
rect 198108 375262 198707 375264
rect 198108 375260 198114 375262
rect 198641 375259 198707 375262
rect 217041 375322 217107 375325
rect 217961 375322 218027 375325
rect 217041 375320 218027 375322
rect 217041 375264 217046 375320
rect 217102 375264 217966 375320
rect 218022 375264 218027 375320
rect 217041 375262 218027 375264
rect 217041 375259 217107 375262
rect 217961 375259 218027 375262
rect 51073 375050 51139 375053
rect 105445 375052 105511 375053
rect 105445 375050 105492 375052
rect 51073 375048 103530 375050
rect 51073 374992 51078 375048
rect 51134 374992 103530 375048
rect 51073 374990 103530 374992
rect 105400 375048 105492 375050
rect 105400 374992 105450 375048
rect 105400 374990 105492 374992
rect 51073 374987 51139 374990
rect 103470 374914 103530 374990
rect 105445 374988 105492 374990
rect 105556 374988 105562 375052
rect 217041 375050 217107 375053
rect 263685 375052 263751 375053
rect 263685 375050 263732 375052
rect 113130 375048 217107 375050
rect 113130 374992 217046 375048
rect 217102 374992 217107 375048
rect 113130 374990 217107 374992
rect 263640 375048 263732 375050
rect 263640 374992 263690 375048
rect 263640 374990 263732 374992
rect 105445 374987 105511 374988
rect 113130 374914 113190 374990
rect 217041 374987 217107 374990
rect 263685 374988 263732 374990
rect 263796 374988 263802 375052
rect 311801 375050 311867 375053
rect 407757 375052 407823 375053
rect 418245 375052 418311 375053
rect 440325 375052 440391 375053
rect 443085 375052 443151 375053
rect 315246 375050 315252 375052
rect 311801 375048 315252 375050
rect 311801 374992 311806 375048
rect 311862 374992 315252 375048
rect 311801 374990 315252 374992
rect 263685 374987 263751 374988
rect 311801 374987 311867 374990
rect 315246 374988 315252 374990
rect 315316 374988 315322 375052
rect 407757 375050 407804 375052
rect 407712 375048 407804 375050
rect 407712 374992 407762 375048
rect 407712 374990 407804 374992
rect 407757 374988 407804 374990
rect 407868 374988 407874 375052
rect 418245 375050 418292 375052
rect 418200 375048 418292 375050
rect 418200 374992 418250 375048
rect 418200 374990 418292 374992
rect 418245 374988 418292 374990
rect 418356 374988 418362 375052
rect 440325 375050 440372 375052
rect 440280 375048 440372 375050
rect 440280 374992 440330 375048
rect 440280 374990 440372 374992
rect 440325 374988 440372 374990
rect 440436 374988 440442 375052
rect 443085 375050 443132 375052
rect 443040 375048 443132 375050
rect 443040 374992 443090 375048
rect 443040 374990 443132 374992
rect 443085 374988 443132 374990
rect 443196 374988 443202 375052
rect 407757 374987 407823 374988
rect 418245 374987 418311 374988
rect 440325 374987 440391 374988
rect 443085 374987 443151 374988
rect 140957 374916 141023 374917
rect 103470 374854 113190 374914
rect 140920 374852 140926 374916
rect 140990 374914 141023 374916
rect 140990 374912 141082 374914
rect 141018 374856 141082 374912
rect 140990 374854 141082 374856
rect 140990 374852 141023 374854
rect 140957 374851 141023 374852
rect 314561 374778 314627 374781
rect 317822 374778 317828 374780
rect 314561 374776 317828 374778
rect 314561 374720 314566 374776
rect 314622 374720 317828 374776
rect 314561 374718 317828 374720
rect 314561 374715 314627 374718
rect 317822 374716 317828 374718
rect 317892 374716 317898 374780
rect 163405 374644 163471 374645
rect 165981 374644 166047 374645
rect 163360 374580 163366 374644
rect 163430 374642 163471 374644
rect 163430 374640 163522 374642
rect 163466 374584 163522 374640
rect 163430 374582 163522 374584
rect 163430 374580 163471 374582
rect 165944 374580 165950 374644
rect 166014 374642 166047 374644
rect 179321 374642 179387 374645
rect 200573 374642 200639 374645
rect 410701 374644 410767 374645
rect 410701 374642 410742 374644
rect 166014 374640 166106 374642
rect 166042 374584 166106 374640
rect 166014 374582 166106 374584
rect 179321 374640 200639 374642
rect 179321 374584 179326 374640
rect 179382 374584 200578 374640
rect 200634 374584 200639 374640
rect 179321 374582 200639 374584
rect 410650 374640 410742 374642
rect 410650 374584 410706 374640
rect 410650 374582 410742 374584
rect 166014 374580 166047 374582
rect 163405 374579 163471 374580
rect 165981 374579 166047 374580
rect 179321 374579 179387 374582
rect 200573 374579 200639 374582
rect 410701 374580 410742 374582
rect 410806 374580 410812 374644
rect 410701 374579 410767 374580
rect 143533 374508 143599 374509
rect 153469 374508 153535 374509
rect 158529 374508 158595 374509
rect 160921 374508 160987 374509
rect 244273 374508 244339 374509
rect 143504 374444 143510 374508
rect 143574 374506 143599 374508
rect 143574 374504 143666 374506
rect 143594 374448 143666 374504
rect 143574 374446 143666 374448
rect 143574 374444 143599 374446
rect 153432 374444 153438 374508
rect 153502 374506 153535 374508
rect 153502 374504 153594 374506
rect 153530 374448 153594 374504
rect 153502 374446 153594 374448
rect 153502 374444 153535 374446
rect 158478 374444 158484 374508
rect 158548 374506 158595 374508
rect 158548 374504 158640 374506
rect 158590 374448 158640 374504
rect 158548 374446 158640 374448
rect 158548 374444 158595 374446
rect 160912 374444 160918 374508
rect 160982 374506 160988 374508
rect 160982 374446 161074 374506
rect 160982 374444 160988 374446
rect 244222 374444 244228 374508
rect 244292 374506 244339 374508
rect 248689 374508 248755 374509
rect 250069 374508 250135 374509
rect 271137 374508 271203 374509
rect 275829 374508 275895 374509
rect 248689 374506 248702 374508
rect 244292 374504 244384 374506
rect 244334 374448 244384 374504
rect 244292 374446 244384 374448
rect 248610 374504 248702 374506
rect 248610 374448 248694 374504
rect 248610 374446 248702 374448
rect 244292 374444 244339 374446
rect 143533 374443 143599 374444
rect 153469 374443 153535 374444
rect 158529 374443 158595 374444
rect 160921 374443 160987 374444
rect 244273 374443 244339 374444
rect 248689 374444 248702 374446
rect 248766 374444 248772 374508
rect 250056 374444 250062 374508
rect 250126 374506 250135 374508
rect 271136 374506 271142 374508
rect 250126 374504 250218 374506
rect 250130 374448 250218 374504
rect 250126 374446 250218 374448
rect 271050 374446 271142 374506
rect 250126 374444 250135 374446
rect 271136 374444 271142 374446
rect 271206 374444 271212 374508
rect 275760 374506 275766 374508
rect 275738 374446 275766 374506
rect 275760 374444 275766 374446
rect 275830 374504 275895 374508
rect 320909 374508 320975 374509
rect 433333 374508 433399 374509
rect 433609 374508 433675 374509
rect 320909 374506 320918 374508
rect 275830 374448 275834 374504
rect 275890 374448 275895 374504
rect 275830 374444 275895 374448
rect 320826 374504 320918 374506
rect 320826 374448 320914 374504
rect 320826 374446 320918 374448
rect 248689 374443 248755 374444
rect 250069 374443 250135 374444
rect 271137 374443 271203 374444
rect 275829 374443 275895 374444
rect 320909 374444 320918 374446
rect 320982 374444 320988 374508
rect 433312 374444 433318 374508
rect 433382 374506 433399 374508
rect 433382 374504 433474 374506
rect 433394 374448 433474 374504
rect 433382 374446 433474 374448
rect 433382 374444 433399 374446
rect 433584 374444 433590 374508
rect 433654 374506 433675 374508
rect 445937 374508 446003 374509
rect 448237 374508 448303 374509
rect 445937 374506 445966 374508
rect 433654 374504 433746 374506
rect 433670 374448 433746 374504
rect 433654 374446 433746 374448
rect 445874 374504 445966 374506
rect 445874 374448 445942 374504
rect 445874 374446 445966 374448
rect 433654 374444 433675 374446
rect 320909 374443 320975 374444
rect 433333 374443 433399 374444
rect 433609 374443 433675 374444
rect 445937 374444 445966 374446
rect 446030 374444 446036 374508
rect 448237 374506 448278 374508
rect 448186 374504 448278 374506
rect 448186 374448 448242 374504
rect 448186 374446 448278 374448
rect 448237 374444 448278 374446
rect 448342 374444 448348 374508
rect 445937 374443 446003 374444
rect 448237 374443 448303 374444
rect 148961 374372 149027 374373
rect 148910 374308 148916 374372
rect 148980 374370 149027 374372
rect 148980 374368 149072 374370
rect 149022 374312 149072 374368
rect 148980 374310 149072 374312
rect 148980 374308 149027 374310
rect 148961 374307 149027 374308
rect 146201 374236 146267 374237
rect 415669 374236 415735 374237
rect 434805 374236 434871 374237
rect 146150 374172 146156 374236
rect 146220 374234 146267 374236
rect 146220 374232 146312 374234
rect 146262 374176 146312 374232
rect 146220 374174 146312 374176
rect 146220 374172 146267 374174
rect 217542 374172 217548 374236
rect 217612 374234 217618 374236
rect 415669 374234 415716 374236
rect 217612 374174 219450 374234
rect 415624 374232 415716 374234
rect 415624 374176 415674 374232
rect 415624 374174 415716 374176
rect 217612 374172 217618 374174
rect 146201 374171 146267 374172
rect 219390 374101 219450 374174
rect 415669 374172 415716 374174
rect 415780 374172 415786 374236
rect 434805 374234 434852 374236
rect 434760 374232 434852 374234
rect 434760 374176 434810 374232
rect 434760 374174 434852 374176
rect 434805 374172 434852 374174
rect 434916 374172 434922 374236
rect 415669 374171 415735 374172
rect 434805 374171 434871 374172
rect 219390 374098 219499 374101
rect 266302 374098 266308 374100
rect 219390 374096 266308 374098
rect 219390 374040 219438 374096
rect 219494 374040 266308 374096
rect 219390 374038 266308 374040
rect 219433 374035 219499 374038
rect 266302 374036 266308 374038
rect 266372 374036 266378 374100
rect 50797 373962 50863 373965
rect 216857 373962 216923 373965
rect 258073 373964 258139 373965
rect 50797 373960 216923 373962
rect 50797 373904 50802 373960
rect 50858 373904 216862 373960
rect 216918 373904 216923 373960
rect 50797 373902 216923 373904
rect 50797 373899 50863 373902
rect 216857 373899 216923 373902
rect 258022 373900 258028 373964
rect 258092 373962 258139 373964
rect 375189 373962 375255 373965
rect 376886 373962 376892 373964
rect 258092 373960 258184 373962
rect 258134 373904 258184 373960
rect 258092 373902 258184 373904
rect 375189 373960 376892 373962
rect 375189 373904 375194 373960
rect 375250 373904 376892 373960
rect 375189 373902 376892 373904
rect 258092 373900 258139 373902
rect 258073 373899 258139 373900
rect 375189 373899 375255 373902
rect 376886 373900 376892 373902
rect 376956 373962 376962 373964
rect 435214 373962 435220 373964
rect 376956 373902 435220 373962
rect 376956 373900 376962 373902
rect 435214 373900 435220 373902
rect 435284 373900 435290 373964
rect 98126 373764 98132 373828
rect 98196 373826 98202 373828
rect 98361 373826 98427 373829
rect 98196 373824 98427 373826
rect 98196 373768 98366 373824
rect 98422 373768 98427 373824
rect 98196 373766 98427 373768
rect 98196 373764 98202 373766
rect 98361 373763 98427 373766
rect 103278 373764 103284 373828
rect 103348 373826 103354 373828
rect 103513 373826 103579 373829
rect 110413 373828 110479 373829
rect 110413 373826 110460 373828
rect 103348 373824 103579 373826
rect 103348 373768 103518 373824
rect 103574 373768 103579 373824
rect 103348 373766 103579 373768
rect 110368 373824 110460 373826
rect 110368 373768 110418 373824
rect 110368 373766 110460 373768
rect 103348 373764 103354 373766
rect 103513 373763 103579 373766
rect 110413 373764 110460 373766
rect 110524 373764 110530 373828
rect 113130 373766 205650 373826
rect 110413 373763 110479 373764
rect 95049 373692 95115 373693
rect 94998 373690 95004 373692
rect 94958 373630 95004 373690
rect 95068 373688 95115 373692
rect 95110 373632 95115 373688
rect 94998 373628 95004 373630
rect 95068 373628 95115 373632
rect 95918 373628 95924 373692
rect 95988 373690 95994 373692
rect 96153 373690 96219 373693
rect 95988 373688 96219 373690
rect 95988 373632 96158 373688
rect 96214 373632 96219 373688
rect 95988 373630 96219 373632
rect 95988 373628 95994 373630
rect 95049 373627 95115 373628
rect 96153 373627 96219 373630
rect 97574 373628 97580 373692
rect 97644 373690 97650 373692
rect 113130 373690 113190 373766
rect 113541 373692 113607 373693
rect 116117 373692 116183 373693
rect 118325 373692 118391 373693
rect 121361 373692 121427 373693
rect 124121 373692 124187 373693
rect 113541 373690 113588 373692
rect 97644 373630 113190 373690
rect 113496 373688 113588 373690
rect 113496 373632 113546 373688
rect 113496 373630 113588 373632
rect 97644 373628 97650 373630
rect 113541 373628 113588 373630
rect 113652 373628 113658 373692
rect 116117 373690 116164 373692
rect 116072 373688 116164 373690
rect 116072 373632 116122 373688
rect 116072 373630 116164 373632
rect 116117 373628 116164 373630
rect 116228 373628 116234 373692
rect 118325 373690 118372 373692
rect 118280 373688 118372 373690
rect 118280 373632 118330 373688
rect 118280 373630 118372 373632
rect 118325 373628 118372 373630
rect 118436 373628 118442 373692
rect 121310 373690 121316 373692
rect 121270 373630 121316 373690
rect 121380 373688 121427 373692
rect 124070 373690 124076 373692
rect 121422 373632 121427 373688
rect 121310 373628 121316 373630
rect 121380 373628 121427 373632
rect 124030 373630 124076 373690
rect 124140 373688 124187 373692
rect 125685 373692 125751 373693
rect 128905 373692 128971 373693
rect 125685 373690 125732 373692
rect 124182 373632 124187 373688
rect 124070 373628 124076 373630
rect 124140 373628 124187 373632
rect 125640 373688 125732 373690
rect 125640 373632 125690 373688
rect 125640 373630 125732 373632
rect 113541 373627 113607 373628
rect 116117 373627 116183 373628
rect 118325 373627 118391 373628
rect 121361 373627 121427 373628
rect 124121 373627 124187 373628
rect 125685 373628 125732 373630
rect 125796 373628 125802 373692
rect 128854 373690 128860 373692
rect 128814 373630 128860 373690
rect 128924 373688 128971 373692
rect 128966 373632 128971 373688
rect 128854 373628 128860 373630
rect 128924 373628 128971 373632
rect 125685 373627 125751 373628
rect 128905 373627 128971 373628
rect 131021 373692 131087 373693
rect 133689 373692 133755 373693
rect 136449 373692 136515 373693
rect 139209 373692 139275 373693
rect 151721 373692 151787 373693
rect 131021 373688 131068 373692
rect 131132 373690 131138 373692
rect 133638 373690 133644 373692
rect 131021 373632 131026 373688
rect 131021 373628 131068 373632
rect 131132 373630 131178 373690
rect 133598 373630 133644 373690
rect 133708 373688 133755 373692
rect 136398 373690 136404 373692
rect 133750 373632 133755 373688
rect 131132 373628 131138 373630
rect 133638 373628 133644 373630
rect 133708 373628 133755 373632
rect 136358 373630 136404 373690
rect 136468 373688 136515 373692
rect 139158 373690 139164 373692
rect 136510 373632 136515 373688
rect 136398 373628 136404 373630
rect 136468 373628 136515 373632
rect 139118 373630 139164 373690
rect 139228 373688 139275 373692
rect 151670 373690 151676 373692
rect 139270 373632 139275 373688
rect 139158 373628 139164 373630
rect 139228 373628 139275 373632
rect 151630 373630 151676 373690
rect 151740 373688 151787 373692
rect 151782 373632 151787 373688
rect 151670 373628 151676 373630
rect 151740 373628 151787 373632
rect 205590 373690 205650 373766
rect 212758 373764 212764 373828
rect 212828 373826 212834 373828
rect 213821 373826 213887 373829
rect 404813 373828 404879 373829
rect 421005 373828 421071 373829
rect 423029 373828 423095 373829
rect 425421 373828 425487 373829
rect 439405 373828 439471 373829
rect 460933 373828 460999 373829
rect 212828 373824 213887 373826
rect 212828 373768 213826 373824
rect 213882 373768 213887 373824
rect 212828 373766 213887 373768
rect 212828 373764 212834 373766
rect 213821 373763 213887 373766
rect 217358 373764 217364 373828
rect 217428 373826 217434 373828
rect 268510 373826 268516 373828
rect 217428 373766 268516 373826
rect 217428 373764 217434 373766
rect 268510 373764 268516 373766
rect 268580 373764 268586 373828
rect 404813 373826 404860 373828
rect 404768 373824 404860 373826
rect 404768 373768 404818 373824
rect 404768 373766 404860 373768
rect 404813 373764 404860 373766
rect 404924 373764 404930 373828
rect 421005 373826 421052 373828
rect 420960 373824 421052 373826
rect 420960 373768 421010 373824
rect 420960 373766 421052 373768
rect 421005 373764 421052 373766
rect 421116 373764 421122 373828
rect 423029 373826 423076 373828
rect 422984 373824 423076 373826
rect 422984 373768 423034 373824
rect 422984 373766 423076 373768
rect 423029 373764 423076 373766
rect 423140 373764 423146 373828
rect 425421 373826 425468 373828
rect 425376 373824 425468 373826
rect 425376 373768 425426 373824
rect 425376 373766 425468 373768
rect 425421 373764 425468 373766
rect 425532 373764 425538 373828
rect 439405 373824 439452 373828
rect 439516 373826 439522 373828
rect 439405 373768 439410 373824
rect 439405 373764 439452 373768
rect 439516 373766 439562 373826
rect 460933 373824 460980 373828
rect 461044 373826 461050 373828
rect 460933 373768 460938 373824
rect 439516 373764 439522 373766
rect 460933 373764 460980 373768
rect 461044 373766 461090 373826
rect 461044 373764 461050 373766
rect 404813 373763 404879 373764
rect 421005 373763 421071 373764
rect 423029 373763 423095 373764
rect 425421 373763 425487 373764
rect 439405 373763 439471 373764
rect 460933 373763 460999 373764
rect 212809 373690 212875 373693
rect 212993 373690 213059 373693
rect 236453 373692 236519 373693
rect 242893 373692 242959 373693
rect 450261 373692 450327 373693
rect 236453 373690 236500 373692
rect 205590 373688 213059 373690
rect 205590 373632 212814 373688
rect 212870 373632 212998 373688
rect 213054 373632 213059 373688
rect 205590 373630 213059 373632
rect 236408 373688 236500 373690
rect 236408 373632 236458 373688
rect 236408 373630 236500 373632
rect 131021 373627 131087 373628
rect 133689 373627 133755 373628
rect 136449 373627 136515 373628
rect 139209 373627 139275 373628
rect 151721 373627 151787 373628
rect 212809 373627 212875 373630
rect 212993 373627 213059 373630
rect 236453 373628 236500 373630
rect 236564 373628 236570 373692
rect 242893 373690 242940 373692
rect 242848 373688 242940 373690
rect 242848 373632 242898 373688
rect 242848 373630 242940 373632
rect 242893 373628 242940 373630
rect 243004 373628 243010 373692
rect 450261 373690 450308 373692
rect 450216 373688 450308 373690
rect 450216 373632 450266 373688
rect 450216 373630 450308 373632
rect 450261 373628 450308 373630
rect 450372 373628 450378 373692
rect 236453 373627 236519 373628
rect 242893 373627 242959 373628
rect 450261 373627 450327 373628
rect 98269 373556 98335 373557
rect 107837 373556 107903 373557
rect 156505 373556 156571 373557
rect 98269 373554 98316 373556
rect 98224 373552 98316 373554
rect 98224 373496 98274 373552
rect 98224 373494 98316 373496
rect 98269 373492 98316 373494
rect 98380 373492 98386 373556
rect 107837 373554 107884 373556
rect 107792 373552 107884 373554
rect 107792 373496 107842 373552
rect 107792 373494 107884 373496
rect 107837 373492 107884 373494
rect 107948 373492 107954 373556
rect 156454 373554 156460 373556
rect 156414 373494 156460 373554
rect 156524 373552 156571 373556
rect 452837 373556 452903 373557
rect 458173 373556 458239 373557
rect 462773 373556 462839 373557
rect 452837 373554 452884 373556
rect 156566 373496 156571 373552
rect 156454 373492 156460 373494
rect 156524 373492 156571 373496
rect 452792 373552 452884 373554
rect 452792 373496 452842 373552
rect 452792 373494 452884 373496
rect 98269 373491 98335 373492
rect 107837 373491 107903 373492
rect 156505 373491 156571 373492
rect 452837 373492 452884 373494
rect 452948 373492 452954 373556
rect 458173 373554 458220 373556
rect 458128 373552 458220 373554
rect 458128 373496 458178 373552
rect 458128 373494 458220 373496
rect 458173 373492 458220 373494
rect 458284 373492 458290 373556
rect 462773 373554 462820 373556
rect 462728 373552 462820 373554
rect 462728 373496 462778 373552
rect 462728 373494 462820 373496
rect 462773 373492 462820 373494
rect 462884 373492 462890 373556
rect 452837 373491 452903 373492
rect 458173 373491 458239 373492
rect 462773 373491 462839 373492
rect 90173 373420 90239 373421
rect 96061 373420 96127 373421
rect 90173 373418 90220 373420
rect 90128 373416 90220 373418
rect 90128 373360 90178 373416
rect 90128 373358 90220 373360
rect 90173 373356 90220 373358
rect 90284 373356 90290 373420
rect 96061 373418 96108 373420
rect 96016 373416 96108 373418
rect 96016 373360 96066 373416
rect 96016 373358 96108 373360
rect 96061 373356 96108 373358
rect 96172 373356 96178 373420
rect 208117 373418 208183 373421
rect 269205 373420 269271 373421
rect 455413 373420 455479 373421
rect 217358 373418 217364 373420
rect 208117 373416 217364 373418
rect 208117 373360 208122 373416
rect 208178 373360 217364 373416
rect 208117 373358 217364 373360
rect 90173 373355 90239 373356
rect 96061 373355 96127 373356
rect 208117 373355 208183 373358
rect 217358 373356 217364 373358
rect 217428 373356 217434 373420
rect 269205 373418 269252 373420
rect 269160 373416 269252 373418
rect 269160 373360 269210 373416
rect 269160 373358 269252 373360
rect 269205 373356 269252 373358
rect 269316 373356 269322 373420
rect 455413 373418 455460 373420
rect 455368 373416 455460 373418
rect 455368 373360 455418 373416
rect 455368 373358 455460 373360
rect 455413 373356 455460 373358
rect 455524 373356 455530 373420
rect 269205 373355 269271 373356
rect 455413 373355 455479 373356
rect 88333 373284 88399 373285
rect 100845 373284 100911 373285
rect 88333 373282 88380 373284
rect 88288 373280 88380 373282
rect 88288 373224 88338 373280
rect 88288 373222 88380 373224
rect 88333 373220 88380 373222
rect 88444 373220 88450 373284
rect 100845 373282 100892 373284
rect 100800 373280 100892 373282
rect 100800 373224 100850 373280
rect 100800 373222 100892 373224
rect 100845 373220 100892 373222
rect 100956 373220 100962 373284
rect 203057 373282 203123 373285
rect 213085 373282 213151 373285
rect 253933 373284 253999 373285
rect 255405 373284 255471 373285
rect 256693 373284 256759 373285
rect 235942 373282 235948 373284
rect 203057 373280 235948 373282
rect 203057 373224 203062 373280
rect 203118 373224 213090 373280
rect 213146 373224 235948 373280
rect 203057 373222 235948 373224
rect 88333 373219 88399 373220
rect 100845 373219 100911 373220
rect 203057 373219 203123 373222
rect 213085 373219 213151 373222
rect 235942 373220 235948 373222
rect 236012 373220 236018 373284
rect 253933 373282 253980 373284
rect 253888 373280 253980 373282
rect 253888 373224 253938 373280
rect 253888 373222 253980 373224
rect 253933 373220 253980 373222
rect 254044 373220 254050 373284
rect 255405 373282 255452 373284
rect 255360 373280 255452 373282
rect 255360 373224 255410 373280
rect 255360 373222 255452 373224
rect 255405 373220 255452 373222
rect 255516 373220 255522 373284
rect 256693 373282 256740 373284
rect 256648 373280 256740 373282
rect 256648 373224 256698 373280
rect 256648 373222 256740 373224
rect 256693 373220 256740 373222
rect 256804 373220 256810 373284
rect 253933 373219 253999 373220
rect 255405 373219 255471 373220
rect 256693 373219 256759 373220
rect 92381 373148 92447 373149
rect 93669 373148 93735 373149
rect 247125 373148 247191 373149
rect 261293 373148 261359 373149
rect 264973 373148 265039 373149
rect 300853 373148 300919 373149
rect 438209 373148 438275 373149
rect 92381 373144 92428 373148
rect 92492 373146 92498 373148
rect 93669 373146 93716 373148
rect 92381 373088 92386 373144
rect 92381 373084 92428 373088
rect 92492 373086 92538 373146
rect 93624 373144 93716 373146
rect 93624 373088 93674 373144
rect 93624 373086 93716 373088
rect 92492 373084 92498 373086
rect 93669 373084 93716 373086
rect 93780 373084 93786 373148
rect 247125 373146 247172 373148
rect 247080 373144 247172 373146
rect 247080 373088 247130 373144
rect 247080 373086 247172 373088
rect 247125 373084 247172 373086
rect 247236 373084 247242 373148
rect 261293 373146 261340 373148
rect 261248 373144 261340 373146
rect 261248 373088 261298 373144
rect 261248 373086 261340 373088
rect 261293 373084 261340 373086
rect 261404 373084 261410 373148
rect 264973 373146 265020 373148
rect 264928 373144 265020 373146
rect 264928 373088 264978 373144
rect 264928 373086 265020 373088
rect 264973 373084 265020 373086
rect 265084 373084 265090 373148
rect 300853 373146 300900 373148
rect 300808 373144 300900 373146
rect 300808 373088 300858 373144
rect 300808 373086 300900 373088
rect 300853 373084 300900 373086
rect 300964 373084 300970 373148
rect 438158 373146 438164 373148
rect 438118 373086 438164 373146
rect 438228 373144 438275 373148
rect 438270 373088 438275 373144
rect 438158 373084 438164 373086
rect 438228 373084 438275 373088
rect 92381 373083 92447 373084
rect 93669 373083 93735 373084
rect 247125 373083 247191 373084
rect 261293 373083 261359 373084
rect 264973 373083 265039 373084
rect 300853 373083 300919 373084
rect 438209 373083 438275 373084
rect 216622 372812 216628 372876
rect 216692 372874 216698 372876
rect 218145 372874 218211 372877
rect 219341 372874 219407 372877
rect 216692 372872 219407 372874
rect 216692 372816 218150 372872
rect 218206 372816 219346 372872
rect 219402 372816 219407 372872
rect 216692 372814 219407 372816
rect 216692 372812 216698 372814
rect 218145 372811 218211 372814
rect 219341 372811 219407 372814
rect 52126 372676 52132 372740
rect 52196 372738 52202 372740
rect 52269 372738 52335 372741
rect 52196 372736 52335 372738
rect 52196 372680 52274 372736
rect 52330 372680 52335 372736
rect 52196 372678 52335 372680
rect 52196 372676 52202 372678
rect 52269 372675 52335 372678
rect 55438 372676 55444 372740
rect 55508 372738 55514 372740
rect 56225 372738 56291 372741
rect 55508 372736 56291 372738
rect 55508 372680 56230 372736
rect 56286 372680 56291 372736
rect 55508 372678 56291 372680
rect 55508 372676 55514 372678
rect 56225 372675 56291 372678
rect 216673 372738 216739 372741
rect 216806 372738 216812 372740
rect 216673 372736 216812 372738
rect 216673 372680 216678 372736
rect 216734 372680 216812 372736
rect 216673 372678 216812 372680
rect 216673 372675 216739 372678
rect 216806 372676 216812 372678
rect 216876 372676 216882 372740
rect 375281 372738 375347 372741
rect 378041 372740 378107 372741
rect 376702 372738 376708 372740
rect 375281 372736 376708 372738
rect 375281 372680 375286 372736
rect 375342 372680 376708 372736
rect 375281 372678 376708 372680
rect 375281 372675 375347 372678
rect 376702 372676 376708 372678
rect 376772 372676 376778 372740
rect 377990 372738 377996 372740
rect 377950 372678 377996 372738
rect 378060 372736 378107 372740
rect 378102 372680 378107 372736
rect 377990 372676 377996 372678
rect 378060 372676 378107 372680
rect 378041 372675 378107 372676
rect 84745 372604 84811 372605
rect 86769 372604 86835 372605
rect 88057 372604 88123 372605
rect 89345 372604 89411 372605
rect 84694 372602 84700 372604
rect 84654 372542 84700 372602
rect 84764 372600 84811 372604
rect 86718 372602 86724 372604
rect 84806 372544 84811 372600
rect 84694 372540 84700 372542
rect 84764 372540 84811 372544
rect 86678 372542 86724 372602
rect 86788 372600 86835 372604
rect 88006 372602 88012 372604
rect 86830 372544 86835 372600
rect 86718 372540 86724 372542
rect 86788 372540 86835 372544
rect 87966 372542 88012 372602
rect 88076 372600 88123 372604
rect 89294 372602 89300 372604
rect 88118 372544 88123 372600
rect 88006 372540 88012 372542
rect 88076 372540 88123 372544
rect 89254 372542 89300 372602
rect 89364 372600 89411 372604
rect 89406 372544 89411 372600
rect 89294 372540 89300 372542
rect 89364 372540 89411 372544
rect 90030 372540 90036 372604
rect 90100 372602 90106 372604
rect 90909 372602 90975 372605
rect 91553 372604 91619 372605
rect 93393 372604 93459 372605
rect 100017 372604 100083 372605
rect 104617 372604 104683 372605
rect 91502 372602 91508 372604
rect 90100 372600 90975 372602
rect 90100 372544 90914 372600
rect 90970 372544 90975 372600
rect 90100 372542 90975 372544
rect 91462 372542 91508 372602
rect 91572 372600 91619 372604
rect 93342 372602 93348 372604
rect 91614 372544 91619 372600
rect 90100 372540 90106 372542
rect 84745 372539 84811 372540
rect 86769 372539 86835 372540
rect 88057 372539 88123 372540
rect 89345 372539 89411 372540
rect 90909 372539 90975 372542
rect 91502 372540 91508 372542
rect 91572 372540 91619 372544
rect 93302 372542 93348 372602
rect 93412 372600 93459 372604
rect 99966 372602 99972 372604
rect 93454 372544 93459 372600
rect 93342 372540 93348 372542
rect 93412 372540 93459 372544
rect 99926 372542 99972 372602
rect 100036 372600 100083 372604
rect 104566 372602 104572 372604
rect 100078 372544 100083 372600
rect 99966 372540 99972 372542
rect 100036 372540 100083 372544
rect 104526 372542 104572 372602
rect 104636 372600 104683 372604
rect 104678 372544 104683 372600
rect 104566 372540 104572 372542
rect 104636 372540 104683 372544
rect 112846 372540 112852 372604
rect 112916 372602 112922 372604
rect 112989 372602 113055 372605
rect 112916 372600 113055 372602
rect 112916 372544 112994 372600
rect 113050 372544 113055 372600
rect 112916 372542 113055 372544
rect 112916 372540 112922 372542
rect 91553 372539 91619 372540
rect 93393 372539 93459 372540
rect 100017 372539 100083 372540
rect 104617 372539 104683 372540
rect 112989 372539 113055 372542
rect 114461 372604 114527 372605
rect 114461 372600 114508 372604
rect 114572 372602 114578 372604
rect 114461 372544 114466 372600
rect 114461 372540 114508 372544
rect 114572 372542 114618 372602
rect 114572 372540 114578 372542
rect 208342 372540 208348 372604
rect 208412 372602 208418 372604
rect 209681 372602 209747 372605
rect 208412 372600 209747 372602
rect 208412 372544 209686 372600
rect 209742 372544 209747 372600
rect 208412 372542 209747 372544
rect 208412 372540 208418 372542
rect 114461 372539 114527 372540
rect 209681 372539 209747 372542
rect 238109 372604 238175 372605
rect 239121 372604 239187 372605
rect 238109 372600 238156 372604
rect 238220 372602 238226 372604
rect 239070 372602 239076 372604
rect 238109 372544 238114 372600
rect 238109 372540 238156 372544
rect 238220 372542 238266 372602
rect 239030 372542 239076 372602
rect 239140 372600 239187 372604
rect 239182 372544 239187 372600
rect 238220 372540 238226 372542
rect 239070 372540 239076 372542
rect 239140 372540 239187 372544
rect 238109 372539 238175 372540
rect 239121 372539 239187 372540
rect 244273 372602 244339 372605
rect 244774 372602 244780 372604
rect 244273 372600 244780 372602
rect 244273 372544 244278 372600
rect 244334 372544 244780 372600
rect 244273 372542 244780 372544
rect 244273 372539 244339 372542
rect 244774 372540 244780 372542
rect 244844 372540 244850 372604
rect 251173 372602 251239 372605
rect 251950 372602 251956 372604
rect 251173 372600 251956 372602
rect 251173 372544 251178 372600
rect 251234 372544 251956 372600
rect 251173 372542 251956 372544
rect 251173 372539 251239 372542
rect 251950 372540 251956 372542
rect 252020 372540 252026 372604
rect 252553 372602 252619 372605
rect 259453 372604 259519 372605
rect 252870 372602 252876 372604
rect 252553 372600 252876 372602
rect 252553 372544 252558 372600
rect 252614 372544 252876 372600
rect 252553 372542 252876 372544
rect 252553 372539 252619 372542
rect 252870 372540 252876 372542
rect 252940 372540 252946 372604
rect 259453 372602 259500 372604
rect 259408 372600 259500 372602
rect 259408 372544 259458 372600
rect 259408 372542 259500 372544
rect 259453 372540 259500 372542
rect 259564 372540 259570 372604
rect 259637 372602 259703 372605
rect 262213 372604 262279 372605
rect 260046 372602 260052 372604
rect 259637 372600 260052 372602
rect 259637 372544 259642 372600
rect 259698 372544 260052 372600
rect 259637 372542 260052 372544
rect 259453 372539 259519 372540
rect 259637 372539 259703 372542
rect 260046 372540 260052 372542
rect 260116 372540 260122 372604
rect 262213 372602 262260 372604
rect 262168 372600 262260 372602
rect 262168 372544 262218 372600
rect 262168 372542 262260 372544
rect 262213 372540 262260 372542
rect 262324 372540 262330 372604
rect 266353 372602 266419 372605
rect 267038 372602 267044 372604
rect 266353 372600 267044 372602
rect 266353 372544 266358 372600
rect 266414 372544 267044 372600
rect 266353 372542 267044 372544
rect 262213 372539 262279 372540
rect 266353 372539 266419 372542
rect 267038 372540 267044 372542
rect 267108 372540 267114 372604
rect 271873 372602 271939 372605
rect 272558 372602 272564 372604
rect 271873 372600 272564 372602
rect 271873 372544 271878 372600
rect 271934 372544 272564 372600
rect 271873 372542 272564 372544
rect 271873 372539 271939 372542
rect 272558 372540 272564 372542
rect 272628 372540 272634 372604
rect 273253 372602 273319 372605
rect 273846 372602 273852 372604
rect 273253 372600 273852 372602
rect 273253 372544 273258 372600
rect 273314 372544 273852 372600
rect 273253 372542 273852 372544
rect 273253 372539 273319 372542
rect 273846 372540 273852 372542
rect 273916 372540 273922 372604
rect 326061 372602 326127 372605
rect 326654 372602 326660 372604
rect 326061 372600 326660 372602
rect 326061 372544 326066 372600
rect 326122 372544 326660 372600
rect 326061 372542 326660 372544
rect 326061 372539 326127 372542
rect 326654 372540 326660 372542
rect 326724 372540 326730 372604
rect 425053 372602 425119 372605
rect 426433 372604 426499 372605
rect 425278 372602 425284 372604
rect 425053 372600 425284 372602
rect 425053 372544 425058 372600
rect 425114 372544 425284 372600
rect 425053 372542 425284 372544
rect 425053 372539 425119 372542
rect 425278 372540 425284 372542
rect 425348 372540 425354 372604
rect 426382 372540 426388 372604
rect 426452 372602 426499 372604
rect 427813 372602 427879 372605
rect 428590 372602 428596 372604
rect 426452 372600 426544 372602
rect 426494 372544 426544 372600
rect 426452 372542 426544 372544
rect 427813 372600 428596 372602
rect 427813 372544 427818 372600
rect 427874 372544 428596 372600
rect 427813 372542 428596 372544
rect 426452 372540 426499 372542
rect 426433 372539 426499 372540
rect 427813 372539 427879 372542
rect 428590 372540 428596 372542
rect 428660 372540 428666 372604
rect 79501 372466 79567 372469
rect 84561 372468 84627 372469
rect 79910 372466 79916 372468
rect 79501 372464 79916 372466
rect 79501 372408 79506 372464
rect 79562 372408 79916 372464
rect 79501 372406 79916 372408
rect 79501 372403 79567 372406
rect 79910 372404 79916 372406
rect 79980 372404 79986 372468
rect 84510 372466 84516 372468
rect 84470 372406 84516 372466
rect 84580 372464 84627 372468
rect 84622 372408 84627 372464
rect 84510 372404 84516 372406
rect 84580 372404 84627 372408
rect 84561 372403 84627 372404
rect 182725 372466 182791 372469
rect 183134 372466 183140 372468
rect 182725 372464 183140 372466
rect 182725 372408 182730 372464
rect 182786 372408 183140 372464
rect 182725 372406 183140 372408
rect 182725 372403 182791 372406
rect 183134 372404 183140 372406
rect 183204 372404 183210 372468
rect 213913 372466 213979 372469
rect 214281 372466 214347 372469
rect 278998 372466 279004 372468
rect 213913 372464 279004 372466
rect 213913 372408 213918 372464
rect 213974 372408 214286 372464
rect 214342 372408 279004 372464
rect 213913 372406 279004 372408
rect 213913 372403 213979 372406
rect 214281 372403 214347 372406
rect 278998 372404 279004 372406
rect 279068 372466 279074 372468
rect 280061 372466 280127 372469
rect 279068 372464 280127 372466
rect 279068 372408 280066 372464
rect 280122 372408 280127 372464
rect 279068 372406 280127 372408
rect 279068 372404 279074 372406
rect 280061 372403 280127 372406
rect 376702 372404 376708 372468
rect 376772 372466 376778 372468
rect 433558 372466 433564 372468
rect 376772 372406 433564 372466
rect 376772 372404 376778 372406
rect 433558 372404 433564 372406
rect 433628 372404 433634 372468
rect 78305 372332 78371 372333
rect 78254 372330 78260 372332
rect 78214 372270 78260 372330
rect 78324 372328 78371 372332
rect 78366 372272 78371 372328
rect 78254 372268 78260 372270
rect 78324 372268 78371 372272
rect 109534 372268 109540 372332
rect 109604 372330 109610 372332
rect 110137 372330 110203 372333
rect 109604 372328 110203 372330
rect 109604 372272 110142 372328
rect 110198 372272 110203 372328
rect 109604 372270 110203 372272
rect 109604 372268 109610 372270
rect 78305 372267 78371 372268
rect 110137 372267 110203 372270
rect 118182 372268 118188 372332
rect 118252 372330 118258 372332
rect 216305 372330 216371 372333
rect 277526 372330 277532 372332
rect 118252 372328 277532 372330
rect 118252 372272 216310 372328
rect 216366 372272 277532 372328
rect 118252 372270 277532 372272
rect 118252 372268 118258 372270
rect 216305 372267 216371 372270
rect 277526 372268 277532 372270
rect 277596 372268 277602 372332
rect 470593 372330 470659 372333
rect 470726 372330 470732 372332
rect 470593 372328 470732 372330
rect 470593 372272 470598 372328
rect 470654 372272 470732 372328
rect 470593 372270 470732 372272
rect 470593 372267 470659 372270
rect 470726 372268 470732 372270
rect 470796 372268 470802 372332
rect 113214 372132 113220 372196
rect 113284 372194 113290 372196
rect 211613 372194 211679 372197
rect 219525 372194 219591 372197
rect 273294 372194 273300 372196
rect 113284 372192 273300 372194
rect 113284 372136 211618 372192
rect 211674 372136 219530 372192
rect 219586 372136 273300 372192
rect 113284 372134 273300 372136
rect 113284 372132 113290 372134
rect 211613 372131 211679 372134
rect 219525 372131 219591 372134
rect 273294 372132 273300 372134
rect 273364 372132 273370 372196
rect 292573 372194 292639 372197
rect 343173 372196 343239 372197
rect 343449 372196 343515 372197
rect 292798 372194 292804 372196
rect 292573 372192 292804 372194
rect 292573 372136 292578 372192
rect 292634 372136 292804 372192
rect 292573 372134 292804 372136
rect 292573 372131 292639 372134
rect 292798 372132 292804 372134
rect 292868 372132 292874 372196
rect 343173 372192 343220 372196
rect 343284 372194 343290 372196
rect 343173 372136 343178 372192
rect 343173 372132 343220 372136
rect 343284 372134 343330 372194
rect 343284 372132 343290 372134
rect 343398 372132 343404 372196
rect 343468 372194 343515 372196
rect 400254 372194 400260 372196
rect 343468 372192 343560 372194
rect 343510 372136 343560 372192
rect 343468 372134 343560 372136
rect 393270 372134 400260 372194
rect 343468 372132 343515 372134
rect 343173 372131 343239 372132
rect 343449 372131 343515 372132
rect 81433 372058 81499 372061
rect 81934 372058 81940 372060
rect 81433 372056 81940 372058
rect 81433 372000 81438 372056
rect 81494 372000 81940 372056
rect 81433 371998 81940 372000
rect 81433 371995 81499 371998
rect 81934 371996 81940 371998
rect 82004 372058 82010 372060
rect 209497 372058 209563 372061
rect 222101 372058 222167 372061
rect 240542 372058 240548 372060
rect 82004 372056 219450 372058
rect 82004 372000 209502 372056
rect 209558 372000 219450 372056
rect 82004 371998 219450 372000
rect 82004 371996 82010 371998
rect 209497 371995 209563 371998
rect 183277 371924 183343 371925
rect 183277 371920 183324 371924
rect 183388 371922 183394 371924
rect 219390 371922 219450 371998
rect 222101 372056 240548 372058
rect 222101 372000 222106 372056
rect 222162 372000 240548 372056
rect 222101 371998 240548 372000
rect 222101 371995 222167 371998
rect 240542 371996 240548 371998
rect 240612 372058 240618 372060
rect 368381 372058 368447 372061
rect 393270 372058 393330 372134
rect 400254 372132 400260 372134
rect 400324 372132 400330 372196
rect 405733 372194 405799 372197
rect 503161 372196 503227 372197
rect 406142 372194 406148 372196
rect 405733 372192 406148 372194
rect 405733 372136 405738 372192
rect 405794 372136 406148 372192
rect 405733 372134 406148 372136
rect 405733 372131 405799 372134
rect 406142 372132 406148 372134
rect 406212 372132 406218 372196
rect 503110 372194 503116 372196
rect 503070 372134 503116 372194
rect 503180 372192 503227 372196
rect 503222 372136 503227 372192
rect 503110 372132 503116 372134
rect 503180 372132 503227 372136
rect 503161 372131 503227 372132
rect 240612 372056 393330 372058
rect 240612 372000 368386 372056
rect 368442 372000 393330 372056
rect 240612 371998 393330 372000
rect 396073 372058 396139 372061
rect 396206 372058 396212 372060
rect 396073 372056 396212 372058
rect 396073 372000 396078 372056
rect 396134 372000 396212 372056
rect 396073 371998 396212 372000
rect 240612 371996 240618 371998
rect 368381 371995 368447 371998
rect 396073 371995 396139 371998
rect 396206 371996 396212 371998
rect 396276 371996 396282 372060
rect 398833 372058 398899 372061
rect 398966 372058 398972 372060
rect 398833 372056 398972 372058
rect 398833 372000 398838 372056
rect 398894 372000 398972 372056
rect 398833 371998 398972 372000
rect 398833 371995 398899 371998
rect 398966 371996 398972 371998
rect 399036 371996 399042 372060
rect 241646 371922 241652 371924
rect 183277 371864 183282 371920
rect 183277 371860 183324 371864
rect 183388 371862 183434 371922
rect 219390 371862 241652 371922
rect 183388 371860 183394 371862
rect 241646 371860 241652 371862
rect 241716 371860 241722 371924
rect 245653 371922 245719 371925
rect 245878 371922 245884 371924
rect 245653 371920 245884 371922
rect 245653 371864 245658 371920
rect 245714 371864 245884 371920
rect 245653 371862 245884 371864
rect 183277 371859 183343 371860
rect 245653 371859 245719 371862
rect 245878 371860 245884 371862
rect 245948 371860 245954 371924
rect 246021 371922 246087 371925
rect 372429 371922 372495 371925
rect 397453 371924 397519 371925
rect 397453 371922 397500 371924
rect 246021 371920 393330 371922
rect 246021 371864 246026 371920
rect 246082 371864 372434 371920
rect 372490 371864 393330 371920
rect 246021 371862 393330 371864
rect 397408 371920 397500 371922
rect 397408 371864 397458 371920
rect 397408 371862 397500 371864
rect 246021 371859 246087 371862
rect 372429 371859 372495 371862
rect 76598 371724 76604 371788
rect 76668 371786 76674 371788
rect 76833 371786 76899 371789
rect 77201 371788 77267 371789
rect 77150 371786 77156 371788
rect 76668 371784 76899 371786
rect 76668 371728 76838 371784
rect 76894 371728 76899 371784
rect 76668 371726 76899 371728
rect 77110 371726 77156 371786
rect 77220 371784 77267 371788
rect 77262 371728 77267 371784
rect 76668 371724 76674 371726
rect 76833 371723 76899 371726
rect 77150 371724 77156 371726
rect 77220 371724 77267 371728
rect 119838 371724 119844 371788
rect 119908 371786 119914 371788
rect 213913 371786 213979 371789
rect 276013 371786 276079 371789
rect 276422 371786 276428 371788
rect 119908 371784 213979 371786
rect 119908 371728 213918 371784
rect 213974 371728 213979 371784
rect 119908 371726 213979 371728
rect 119908 371724 119914 371726
rect 77201 371723 77267 371724
rect 213913 371723 213979 371726
rect 219390 371784 276428 371786
rect 219390 371728 276018 371784
rect 276074 371728 276428 371784
rect 219390 371726 276428 371728
rect 102041 371652 102107 371653
rect 107009 371652 107075 371653
rect 108849 371652 108915 371653
rect 111609 371652 111675 371653
rect 101990 371650 101996 371652
rect 101950 371590 101996 371650
rect 102060 371648 102107 371652
rect 106958 371650 106964 371652
rect 102102 371592 102107 371648
rect 101990 371588 101996 371590
rect 102060 371588 102107 371592
rect 106918 371590 106964 371650
rect 107028 371648 107075 371652
rect 108798 371650 108804 371652
rect 107070 371592 107075 371648
rect 106958 371588 106964 371590
rect 107028 371588 107075 371592
rect 108758 371590 108804 371650
rect 108868 371648 108915 371652
rect 111558 371650 111564 371652
rect 108910 371592 108915 371648
rect 108798 371588 108804 371590
rect 108868 371588 108915 371592
rect 111518 371590 111564 371650
rect 111628 371648 111675 371652
rect 111670 371592 111675 371648
rect 111558 371588 111564 371590
rect 111628 371588 111675 371592
rect 117078 371588 117084 371652
rect 117148 371650 117154 371652
rect 216990 371650 216996 371652
rect 117148 371590 216996 371650
rect 117148 371588 117154 371590
rect 216990 371588 216996 371590
rect 217060 371650 217066 371652
rect 219390 371650 219450 371726
rect 276013 371723 276079 371726
rect 276422 371724 276428 371726
rect 276492 371724 276498 371788
rect 302233 371786 302299 371789
rect 302918 371786 302924 371788
rect 302233 371784 302924 371786
rect 302233 371728 302238 371784
rect 302294 371728 302924 371784
rect 302233 371726 302924 371728
rect 302233 371723 302299 371726
rect 302918 371724 302924 371726
rect 302988 371724 302994 371788
rect 393270 371786 393330 371862
rect 397453 371860 397500 371862
rect 397564 371860 397570 371924
rect 412817 371922 412883 371925
rect 413686 371922 413692 371924
rect 412817 371920 413692 371922
rect 412817 371864 412822 371920
rect 412878 371864 413692 371920
rect 412817 371862 413692 371864
rect 397453 371859 397519 371860
rect 412817 371859 412883 371862
rect 413686 371860 413692 371862
rect 413756 371860 413762 371924
rect 483013 371922 483079 371925
rect 483238 371922 483244 371924
rect 483013 371920 483244 371922
rect 483013 371864 483018 371920
rect 483074 371864 483244 371920
rect 483013 371862 483244 371864
rect 483013 371859 483079 371862
rect 483238 371860 483244 371862
rect 483308 371860 483314 371924
rect 402278 371786 402284 371788
rect 393270 371726 402284 371786
rect 402278 371724 402284 371726
rect 402348 371724 402354 371788
rect 409873 371786 409939 371789
rect 410006 371786 410012 371788
rect 409873 371784 410012 371786
rect 409873 371728 409878 371784
rect 409934 371728 410012 371784
rect 409873 371726 410012 371728
rect 409873 371723 409939 371726
rect 410006 371724 410012 371726
rect 410076 371724 410082 371788
rect 411253 371786 411319 371789
rect 430573 371788 430639 371789
rect 411846 371786 411852 371788
rect 411253 371784 411852 371786
rect 411253 371728 411258 371784
rect 411314 371728 411852 371784
rect 411253 371726 411852 371728
rect 411253 371723 411319 371726
rect 411846 371724 411852 371726
rect 411916 371724 411922 371788
rect 430573 371786 430620 371788
rect 430528 371784 430620 371786
rect 430528 371728 430578 371784
rect 430528 371726 430620 371728
rect 430573 371724 430620 371726
rect 430684 371724 430690 371788
rect 430573 371723 430639 371724
rect 217060 371590 219450 371650
rect 217060 371588 217066 371590
rect 241646 371588 241652 371652
rect 241716 371650 241722 371652
rect 246021 371650 246087 371653
rect 251173 371652 251239 371653
rect 251173 371650 251220 371652
rect 241716 371648 246087 371650
rect 241716 371592 246026 371648
rect 246082 371592 246087 371648
rect 241716 371590 246087 371592
rect 251128 371648 251220 371650
rect 251128 371592 251178 371648
rect 251128 371590 251220 371592
rect 241716 371588 241722 371590
rect 102041 371587 102107 371588
rect 107009 371587 107075 371588
rect 108849 371587 108915 371588
rect 111609 371587 111675 371588
rect 246021 371587 246087 371590
rect 251173 371588 251220 371590
rect 251284 371588 251290 371652
rect 258165 371650 258231 371653
rect 258390 371650 258396 371652
rect 258165 371648 258396 371650
rect 258165 371592 258170 371648
rect 258226 371592 258396 371648
rect 258165 371590 258396 371592
rect 251173 371587 251239 371588
rect 258165 371587 258231 371590
rect 258390 371588 258396 371590
rect 258460 371588 258466 371652
rect 407113 371650 407179 371653
rect 407246 371650 407252 371652
rect 407113 371648 407252 371650
rect 407113 371592 407118 371648
rect 407174 371592 407252 371648
rect 407113 371590 407252 371592
rect 407113 371587 407179 371590
rect 407246 371588 407252 371590
rect 407316 371588 407322 371652
rect 412633 371650 412699 371653
rect 412766 371650 412772 371652
rect 412633 371648 412772 371650
rect 412633 371592 412638 371648
rect 412694 371592 412772 371648
rect 412633 371590 412772 371592
rect 412633 371587 412699 371590
rect 412766 371588 412772 371590
rect 412836 371588 412842 371652
rect 465073 371650 465139 371653
rect 465390 371650 465396 371652
rect 465073 371648 465396 371650
rect 465073 371592 465078 371648
rect 465134 371592 465396 371648
rect 465073 371590 465396 371592
rect 465073 371587 465139 371590
rect 465390 371588 465396 371590
rect 465460 371588 465466 371652
rect 83825 371516 83891 371517
rect 83774 371514 83780 371516
rect 83734 371454 83780 371514
rect 83844 371512 83891 371516
rect 220905 371514 220971 371517
rect 222101 371514 222167 371517
rect 83886 371456 83891 371512
rect 83774 371452 83780 371454
rect 83844 371452 83891 371456
rect 83825 371451 83891 371452
rect 84150 371512 222167 371514
rect 84150 371456 220910 371512
rect 220966 371456 222106 371512
rect 222162 371456 222167 371512
rect 84150 371454 222167 371456
rect 80053 371378 80119 371381
rect 81014 371378 81020 371380
rect 80053 371376 81020 371378
rect 80053 371320 80058 371376
rect 80114 371320 81020 371376
rect 80053 371318 81020 371320
rect 80053 371315 80119 371318
rect 81014 371316 81020 371318
rect 81084 371378 81090 371380
rect 84150 371378 84210 371454
rect 220905 371451 220971 371454
rect 222101 371451 222167 371454
rect 247033 371514 247099 371517
rect 247902 371514 247908 371516
rect 247033 371512 247908 371514
rect 247033 371456 247038 371512
rect 247094 371456 247908 371512
rect 247033 371454 247908 371456
rect 247033 371451 247099 371454
rect 247902 371452 247908 371454
rect 247972 371452 247978 371516
rect 249793 371514 249859 371517
rect 250294 371514 250300 371516
rect 249793 371512 250300 371514
rect 249793 371456 249798 371512
rect 249854 371456 250300 371512
rect 249793 371454 250300 371456
rect 249793 371451 249859 371454
rect 250294 371452 250300 371454
rect 250364 371452 250370 371516
rect 252645 371514 252711 371517
rect 253606 371514 253612 371516
rect 252645 371512 253612 371514
rect 252645 371456 252650 371512
rect 252706 371456 253612 371512
rect 252645 371454 253612 371456
rect 252645 371451 252711 371454
rect 253606 371452 253612 371454
rect 253676 371452 253682 371516
rect 255313 371514 255379 371517
rect 256182 371514 256188 371516
rect 255313 371512 256188 371514
rect 255313 371456 255318 371512
rect 255374 371456 256188 371512
rect 255313 371454 256188 371456
rect 255313 371451 255379 371454
rect 256182 371452 256188 371454
rect 256252 371452 256258 371516
rect 260833 371514 260899 371517
rect 263593 371516 263659 371517
rect 260966 371514 260972 371516
rect 260833 371512 260972 371514
rect 260833 371456 260838 371512
rect 260894 371456 260972 371512
rect 260833 371454 260972 371456
rect 260833 371451 260899 371454
rect 260966 371452 260972 371454
rect 261036 371452 261042 371516
rect 263542 371452 263548 371516
rect 263612 371514 263659 371516
rect 264973 371514 265039 371517
rect 267733 371516 267799 371517
rect 265750 371514 265756 371516
rect 263612 371512 263704 371514
rect 263654 371456 263704 371512
rect 263612 371454 263704 371456
rect 264973 371512 265756 371514
rect 264973 371456 264978 371512
rect 265034 371456 265756 371512
rect 264973 371454 265756 371456
rect 263612 371452 263659 371454
rect 263593 371451 263659 371452
rect 264973 371451 265039 371454
rect 265750 371452 265756 371454
rect 265820 371452 265826 371516
rect 267733 371512 267780 371516
rect 267844 371514 267850 371516
rect 277301 371514 277367 371517
rect 411253 371516 411319 371517
rect 277526 371514 277532 371516
rect 267733 371456 267738 371512
rect 267733 371452 267780 371456
rect 267844 371454 267890 371514
rect 277301 371512 277532 371514
rect 277301 371456 277306 371512
rect 277362 371456 277532 371512
rect 277301 371454 277532 371456
rect 267844 371452 267850 371454
rect 267733 371451 267799 371452
rect 277301 371451 277367 371454
rect 277526 371452 277532 371454
rect 277596 371452 277602 371516
rect 411253 371514 411300 371516
rect 411208 371512 411300 371514
rect 411208 371456 411258 371512
rect 411208 371454 411300 371456
rect 411253 371452 411300 371454
rect 411364 371452 411370 371516
rect 418245 371514 418311 371517
rect 422293 371516 422359 371517
rect 418838 371514 418844 371516
rect 418245 371512 418844 371514
rect 418245 371456 418250 371512
rect 418306 371456 418844 371512
rect 418245 371454 418844 371456
rect 411253 371451 411319 371452
rect 418245 371451 418311 371454
rect 418838 371452 418844 371454
rect 418908 371452 418914 371516
rect 422293 371512 422340 371516
rect 422404 371514 422410 371516
rect 426433 371514 426499 371517
rect 427670 371514 427676 371516
rect 422293 371456 422298 371512
rect 422293 371452 422340 371456
rect 422404 371454 422450 371514
rect 426433 371512 427676 371514
rect 426433 371456 426438 371512
rect 426494 371456 427676 371512
rect 426433 371454 427676 371456
rect 422404 371452 422410 371454
rect 422293 371451 422359 371452
rect 426433 371451 426499 371454
rect 427670 371452 427676 371454
rect 427740 371452 427746 371516
rect 81084 371318 84210 371378
rect 81084 371316 81090 371318
rect 100702 371316 100708 371380
rect 100772 371378 100778 371380
rect 101673 371378 101739 371381
rect 102777 371380 102843 371381
rect 102726 371378 102732 371380
rect 100772 371376 101739 371378
rect 100772 371320 101678 371376
rect 101734 371320 101739 371376
rect 100772 371318 101739 371320
rect 102686 371318 102732 371378
rect 102796 371376 102843 371380
rect 102838 371320 102843 371376
rect 100772 371316 100778 371318
rect 101673 371315 101739 371318
rect 102726 371316 102732 371318
rect 102796 371316 102843 371320
rect 105302 371316 105308 371380
rect 105372 371378 105378 371380
rect 105629 371378 105695 371381
rect 105372 371376 105695 371378
rect 105372 371320 105634 371376
rect 105690 371320 105695 371376
rect 105372 371318 105695 371320
rect 105372 371316 105378 371318
rect 102777 371315 102843 371316
rect 105629 371315 105695 371318
rect 107510 371316 107516 371380
rect 107580 371316 107586 371380
rect 115790 371316 115796 371380
rect 115860 371378 115866 371380
rect 222009 371378 222075 371381
rect 270309 371378 270375 371381
rect 115860 371376 270375 371378
rect 115860 371320 222014 371376
rect 222070 371320 270314 371376
rect 270370 371320 270375 371376
rect 115860 371318 270375 371320
rect 115860 371316 115866 371318
rect 107518 371242 107578 371316
rect 222009 371315 222075 371318
rect 270309 371315 270375 371318
rect 270493 371378 270559 371381
rect 270902 371378 270908 371380
rect 270493 371376 270908 371378
rect 270493 371320 270498 371376
rect 270554 371320 270908 371376
rect 270493 371318 270908 371320
rect 270493 371315 270559 371318
rect 270902 371316 270908 371318
rect 270972 371316 270978 371380
rect 273253 371378 273319 371381
rect 273662 371378 273668 371380
rect 273253 371376 273668 371378
rect 273253 371320 273258 371376
rect 273314 371320 273668 371376
rect 273253 371318 273668 371320
rect 273253 371315 273319 371318
rect 273662 371316 273668 371318
rect 273732 371316 273738 371380
rect 276013 371378 276079 371381
rect 276238 371378 276244 371380
rect 276013 371376 276244 371378
rect 276013 371320 276018 371376
rect 276074 371320 276244 371376
rect 276013 371318 276244 371320
rect 276013 371315 276079 371318
rect 276238 371316 276244 371318
rect 276308 371316 276314 371380
rect 277393 371378 277459 371381
rect 278262 371378 278268 371380
rect 277393 371376 278268 371378
rect 277393 371320 277398 371376
rect 277454 371320 278268 371376
rect 277393 371318 278268 371320
rect 277393 371315 277459 371318
rect 278262 371316 278268 371318
rect 278332 371316 278338 371380
rect 280153 371378 280219 371381
rect 280286 371378 280292 371380
rect 280153 371376 280292 371378
rect 280153 371320 280158 371376
rect 280214 371320 280292 371376
rect 280153 371318 280292 371320
rect 280153 371315 280219 371318
rect 280286 371316 280292 371318
rect 280356 371316 280362 371380
rect 282913 371378 282979 371381
rect 283782 371378 283788 371380
rect 282913 371376 283788 371378
rect 282913 371320 282918 371376
rect 282974 371320 283788 371376
rect 282913 371318 283788 371320
rect 282913 371315 282979 371318
rect 283782 371316 283788 371318
rect 283852 371316 283858 371380
rect 285673 371378 285739 371381
rect 285806 371378 285812 371380
rect 285673 371376 285812 371378
rect 285673 371320 285678 371376
rect 285734 371320 285812 371376
rect 285673 371318 285812 371320
rect 285673 371315 285739 371318
rect 285806 371316 285812 371318
rect 285876 371316 285882 371380
rect 287237 371378 287303 371381
rect 287646 371378 287652 371380
rect 287237 371376 287652 371378
rect 287237 371320 287242 371376
rect 287298 371320 287652 371376
rect 287237 371318 287652 371320
rect 287237 371315 287303 371318
rect 287646 371316 287652 371318
rect 287716 371316 287722 371380
rect 289813 371378 289879 371381
rect 295333 371380 295399 371381
rect 298093 371380 298159 371381
rect 290590 371378 290596 371380
rect 289813 371376 290596 371378
rect 289813 371320 289818 371376
rect 289874 371320 290596 371376
rect 289813 371318 290596 371320
rect 289813 371315 289879 371318
rect 290590 371316 290596 371318
rect 290660 371316 290666 371380
rect 295333 371378 295380 371380
rect 295288 371376 295380 371378
rect 295288 371320 295338 371376
rect 295288 371318 295380 371320
rect 295333 371316 295380 371318
rect 295444 371316 295450 371380
rect 298093 371378 298140 371380
rect 298048 371376 298140 371378
rect 298048 371320 298098 371376
rect 298048 371318 298140 371320
rect 298093 371316 298140 371318
rect 298204 371316 298210 371380
rect 304993 371378 305059 371381
rect 305310 371378 305316 371380
rect 304993 371376 305316 371378
rect 304993 371320 304998 371376
rect 305054 371320 305316 371376
rect 304993 371318 305316 371320
rect 295333 371315 295399 371316
rect 298093 371315 298159 371316
rect 304993 371315 305059 371318
rect 305310 371316 305316 371318
rect 305380 371316 305386 371380
rect 307753 371378 307819 371381
rect 308622 371378 308628 371380
rect 307753 371376 308628 371378
rect 307753 371320 307758 371376
rect 307814 371320 308628 371376
rect 307753 371318 308628 371320
rect 307753 371315 307819 371318
rect 308622 371316 308628 371318
rect 308692 371316 308698 371380
rect 310513 371378 310579 371381
rect 310646 371378 310652 371380
rect 310513 371376 310652 371378
rect 310513 371320 310518 371376
rect 310574 371320 310652 371376
rect 310513 371318 310652 371320
rect 310513 371315 310579 371318
rect 310646 371316 310652 371318
rect 310716 371316 310722 371380
rect 313273 371378 313339 371381
rect 322933 371380 322999 371381
rect 313406 371378 313412 371380
rect 313273 371376 313412 371378
rect 313273 371320 313278 371376
rect 313334 371320 313412 371376
rect 313273 371318 313412 371320
rect 313273 371315 313339 371318
rect 313406 371316 313412 371318
rect 313476 371316 313482 371380
rect 322933 371378 322980 371380
rect 322888 371376 322980 371378
rect 322888 371320 322938 371376
rect 322888 371318 322980 371320
rect 322933 371316 322980 371318
rect 323044 371316 323050 371380
rect 396073 371378 396139 371381
rect 402973 371380 403039 371381
rect 396574 371378 396580 371380
rect 396073 371376 396580 371378
rect 396073 371320 396078 371376
rect 396134 371320 396580 371376
rect 396073 371318 396580 371320
rect 322933 371315 322999 371316
rect 396073 371315 396139 371318
rect 396574 371316 396580 371318
rect 396644 371316 396650 371380
rect 402973 371376 403020 371380
rect 403084 371378 403090 371380
rect 403249 371378 403315 371381
rect 408493 371380 408559 371381
rect 414013 371380 414079 371381
rect 403566 371378 403572 371380
rect 402973 371320 402978 371376
rect 402973 371316 403020 371320
rect 403084 371318 403130 371378
rect 403249 371376 403572 371378
rect 403249 371320 403254 371376
rect 403310 371320 403572 371376
rect 403249 371318 403572 371320
rect 403084 371316 403090 371318
rect 402973 371315 403039 371316
rect 403249 371315 403315 371318
rect 403566 371316 403572 371318
rect 403636 371316 403642 371380
rect 408493 371378 408540 371380
rect 408448 371376 408540 371378
rect 408448 371320 408498 371376
rect 408448 371318 408540 371320
rect 408493 371316 408540 371318
rect 408604 371316 408610 371380
rect 414013 371378 414060 371380
rect 413968 371376 414060 371378
rect 413968 371320 414018 371376
rect 413968 371318 414060 371320
rect 414013 371316 414060 371318
rect 414124 371316 414130 371380
rect 415393 371378 415459 371381
rect 416773 371380 416839 371381
rect 418153 371380 418219 371381
rect 415526 371378 415532 371380
rect 415393 371376 415532 371378
rect 415393 371320 415398 371376
rect 415454 371320 415532 371376
rect 415393 371318 415532 371320
rect 408493 371315 408559 371316
rect 414013 371315 414079 371316
rect 415393 371315 415459 371318
rect 415526 371316 415532 371318
rect 415596 371316 415602 371380
rect 416773 371378 416820 371380
rect 416728 371376 416820 371378
rect 416728 371320 416778 371376
rect 416728 371318 416820 371320
rect 416773 371316 416820 371318
rect 416884 371316 416890 371380
rect 418102 371316 418108 371380
rect 418172 371378 418219 371380
rect 419533 371378 419599 371381
rect 420310 371378 420316 371380
rect 418172 371376 418264 371378
rect 418214 371320 418264 371376
rect 418172 371318 418264 371320
rect 419533 371376 420316 371378
rect 419533 371320 419538 371376
rect 419594 371320 420316 371376
rect 419533 371318 420316 371320
rect 418172 371316 418219 371318
rect 416773 371315 416839 371316
rect 418153 371315 418219 371316
rect 419533 371315 419599 371318
rect 420310 371316 420316 371318
rect 420380 371316 420386 371380
rect 420913 371378 420979 371381
rect 421230 371378 421236 371380
rect 420913 371376 421236 371378
rect 420913 371320 420918 371376
rect 420974 371320 421236 371376
rect 420913 371318 421236 371320
rect 420913 371315 420979 371318
rect 421230 371316 421236 371318
rect 421300 371316 421306 371380
rect 423673 371378 423739 371381
rect 427813 371380 427879 371381
rect 423990 371378 423996 371380
rect 423673 371376 423996 371378
rect 423673 371320 423678 371376
rect 423734 371320 423996 371376
rect 423673 371318 423996 371320
rect 423673 371315 423739 371318
rect 423990 371316 423996 371318
rect 424060 371316 424066 371380
rect 427813 371378 427860 371380
rect 427768 371376 427860 371378
rect 427768 371320 427818 371376
rect 427768 371318 427860 371320
rect 427813 371316 427860 371318
rect 427924 371316 427930 371380
rect 429193 371378 429259 371381
rect 429326 371378 429332 371380
rect 429193 371376 429332 371378
rect 429193 371320 429198 371376
rect 429254 371320 429332 371376
rect 429193 371318 429332 371320
rect 427813 371315 427879 371316
rect 429193 371315 429259 371318
rect 429326 371316 429332 371318
rect 429396 371316 429402 371380
rect 430665 371378 430731 371381
rect 431166 371378 431172 371380
rect 430665 371376 431172 371378
rect 430665 371320 430670 371376
rect 430726 371320 431172 371376
rect 430665 371318 431172 371320
rect 430665 371315 430731 371318
rect 431166 371316 431172 371318
rect 431236 371316 431242 371380
rect 431953 371378 432019 371381
rect 432086 371378 432092 371380
rect 431953 371376 432092 371378
rect 431953 371320 431958 371376
rect 432014 371320 432092 371376
rect 431953 371318 432092 371320
rect 431953 371315 432019 371318
rect 432086 371316 432092 371318
rect 432156 371316 432162 371380
rect 436093 371378 436159 371381
rect 436318 371378 436324 371380
rect 436093 371376 436324 371378
rect 436093 371320 436098 371376
rect 436154 371320 436324 371376
rect 436093 371318 436324 371320
rect 436093 371315 436159 371318
rect 436318 371316 436324 371318
rect 436388 371316 436394 371380
rect 437473 371378 437539 371381
rect 438342 371378 438348 371380
rect 437473 371376 438348 371378
rect 437473 371320 437478 371376
rect 437534 371320 438348 371376
rect 437473 371318 438348 371320
rect 437473 371315 437539 371318
rect 438342 371316 438348 371318
rect 438412 371316 438418 371380
rect 467833 371378 467899 371381
rect 473353 371380 473419 371381
rect 467966 371378 467972 371380
rect 467833 371376 467972 371378
rect 467833 371320 467838 371376
rect 467894 371320 467972 371376
rect 467833 371318 467972 371320
rect 467833 371315 467899 371318
rect 467966 371316 467972 371318
rect 468036 371316 468042 371380
rect 473302 371316 473308 371380
rect 473372 371378 473419 371380
rect 480253 371380 480319 371381
rect 485773 371380 485839 371381
rect 473372 371376 473464 371378
rect 473414 371320 473464 371376
rect 473372 371318 473464 371320
rect 480253 371376 480300 371380
rect 480364 371378 480370 371380
rect 485773 371378 485820 371380
rect 480253 371320 480258 371376
rect 473372 371316 473419 371318
rect 473353 371315 473419 371316
rect 480253 371316 480300 371320
rect 480364 371318 480410 371378
rect 485728 371376 485820 371378
rect 485728 371320 485778 371376
rect 485728 371318 485820 371320
rect 480364 371316 480370 371318
rect 485773 371316 485820 371318
rect 485884 371316 485890 371380
rect 502333 371378 502399 371381
rect 503478 371378 503484 371380
rect 502333 371376 503484 371378
rect 502333 371320 502338 371376
rect 502394 371320 503484 371376
rect 502333 371318 503484 371320
rect 480253 371315 480319 371316
rect 485773 371315 485839 371316
rect 502333 371315 502399 371318
rect 503478 371316 503484 371318
rect 503548 371316 503554 371380
rect 107518 371182 200130 371242
rect 200070 371106 200130 371182
rect 208526 371180 208532 371244
rect 208596 371242 208602 371244
rect 209589 371242 209655 371245
rect 208596 371240 209655 371242
rect 208596 371184 209594 371240
rect 209650 371184 209655 371240
rect 208596 371182 209655 371184
rect 208596 371180 208602 371182
rect 209589 371179 209655 371182
rect 359958 371180 359964 371244
rect 360028 371242 360034 371244
rect 475326 371242 475332 371244
rect 360028 371182 475332 371242
rect 360028 371180 360034 371182
rect 475326 371180 475332 371182
rect 475396 371180 475402 371244
rect 216806 371106 216812 371108
rect 200070 371046 216812 371106
rect 216806 371044 216812 371046
rect 216876 371106 216882 371108
rect 218513 371106 218579 371109
rect 220721 371106 220787 371109
rect 216876 371104 220787 371106
rect 216876 371048 218518 371104
rect 218574 371048 220726 371104
rect 220782 371048 220787 371104
rect 216876 371046 220787 371048
rect 216876 371044 216882 371046
rect 218513 371043 218579 371046
rect 220721 371043 220787 371046
rect 377254 371044 377260 371108
rect 377324 371106 377330 371108
rect 478086 371106 478092 371108
rect 377324 371046 478092 371106
rect 377324 371044 377330 371046
rect 478086 371044 478092 371046
rect 478156 371044 478162 371108
rect -960 370834 480 370924
rect 3509 370834 3575 370837
rect -960 370832 3575 370834
rect -960 370776 3514 370832
rect 3570 370776 3575 370832
rect -960 370774 3575 370776
rect -960 370684 480 370774
rect 3509 370771 3575 370774
rect 110137 370562 110203 370565
rect 211705 370562 211771 370565
rect 216622 370562 216628 370564
rect 110137 370560 216628 370562
rect 110137 370504 110142 370560
rect 110198 370504 211710 370560
rect 211766 370504 216628 370560
rect 110137 370502 216628 370504
rect 110137 370499 110203 370502
rect 211705 370499 211771 370502
rect 216622 370500 216628 370502
rect 216692 370500 216698 370564
rect 377121 370426 377187 370429
rect 377806 370426 377812 370428
rect 377121 370424 377812 370426
rect 377121 370368 377126 370424
rect 377182 370368 377812 370424
rect 377121 370366 377812 370368
rect 377121 370363 377187 370366
rect 377806 370364 377812 370366
rect 377876 370364 377882 370428
rect 215334 369820 215340 369884
rect 215404 369882 215410 369884
rect 216581 369882 216647 369885
rect 215404 369880 216647 369882
rect 215404 369824 216586 369880
rect 216642 369824 216647 369880
rect 215404 369822 216647 369824
rect 215404 369820 215410 369822
rect 216581 369819 216647 369822
rect 379462 369820 379468 369884
rect 379532 369882 379538 369884
rect 379605 369882 379671 369885
rect 379532 369880 379671 369882
rect 379532 369824 379610 369880
rect 379666 369824 379671 369880
rect 379532 369822 379671 369824
rect 379532 369820 379538 369822
rect 379605 369819 379671 369822
rect 209814 369140 209820 369204
rect 209884 369202 209890 369204
rect 211061 369202 211127 369205
rect 209884 369200 211127 369202
rect 209884 369144 211066 369200
rect 211122 369144 211127 369200
rect 209884 369142 211127 369144
rect 209884 369140 209890 369142
rect 211061 369139 211127 369142
rect 211654 369140 211660 369204
rect 211724 369202 211730 369204
rect 212441 369202 212507 369205
rect 211724 369200 212507 369202
rect 211724 369144 212446 369200
rect 212502 369144 212507 369200
rect 211724 369142 212507 369144
rect 211724 369140 211730 369142
rect 212441 369139 212507 369142
rect 213310 369140 213316 369204
rect 213380 369202 213386 369204
rect 213729 369202 213795 369205
rect 213380 369200 213795 369202
rect 213380 369144 213734 369200
rect 213790 369144 213795 369200
rect 213380 369142 213795 369144
rect 213380 369140 213386 369142
rect 213729 369139 213795 369142
rect 213862 369140 213868 369204
rect 213932 369202 213938 369204
rect 215109 369202 215175 369205
rect 213932 369200 215175 369202
rect 213932 369144 215114 369200
rect 215170 369144 215175 369200
rect 213932 369142 215175 369144
rect 213932 369140 213938 369142
rect 215109 369139 215175 369142
rect 107009 369066 107075 369069
rect 218605 369066 218671 369069
rect 219617 369066 219683 369069
rect 107009 369064 219683 369066
rect 107009 369008 107014 369064
rect 107070 369008 218610 369064
rect 218666 369008 219622 369064
rect 219678 369008 219683 369064
rect 107009 369006 219683 369008
rect 107009 369003 107075 369006
rect 218605 369003 218671 369006
rect 219617 369003 219683 369006
rect 359774 369004 359780 369068
rect 359844 369066 359850 369068
rect 372981 369066 373047 369069
rect 420913 369066 420979 369069
rect 359844 369064 420979 369066
rect 359844 369008 372986 369064
rect 373042 369008 420918 369064
rect 420974 369008 420979 369064
rect 359844 369006 420979 369008
rect 359844 369004 359850 369006
rect 372981 369003 373047 369006
rect 420913 369003 420979 369006
rect 199377 366346 199443 366349
rect 199510 366346 199516 366348
rect 199377 366344 199516 366346
rect 199377 366288 199382 366344
rect 199438 366288 199516 366344
rect 199377 366286 199516 366288
rect 199377 366283 199443 366286
rect 199510 366284 199516 366286
rect 199580 366346 199586 366348
rect 359089 366346 359155 366349
rect 199580 366344 359155 366346
rect 199580 366288 359094 366344
rect 359150 366288 359155 366344
rect 199580 366286 359155 366288
rect 199580 366284 199586 366286
rect 359089 366283 359155 366286
rect 580901 364850 580967 364853
rect 583520 364850 584960 364940
rect 580901 364848 584960 364850
rect 580901 364792 580906 364848
rect 580962 364792 584960 364848
rect 580901 364790 584960 364792
rect 580901 364787 580967 364790
rect 583520 364700 584960 364790
rect -960 358322 480 358412
rect 2773 358322 2839 358325
rect -960 358320 2839 358322
rect -960 358264 2778 358320
rect 2834 358264 2839 358320
rect -960 358262 2839 358264
rect -960 358172 480 358262
rect 2773 358259 2839 358262
rect 178534 351868 178540 351932
rect 178604 351930 178610 351932
rect 179321 351930 179387 351933
rect 178604 351928 179387 351930
rect 178604 351872 179326 351928
rect 179382 351872 179387 351928
rect 178604 351870 179387 351872
rect 178604 351868 178610 351870
rect 179321 351867 179387 351870
rect 583520 351780 584960 352020
rect 179689 350572 179755 350573
rect 179638 350570 179644 350572
rect 179598 350510 179644 350570
rect 179708 350568 179755 350572
rect 179750 350512 179755 350568
rect 179638 350508 179644 350510
rect 179708 350508 179755 350512
rect 190862 350508 190868 350572
rect 190932 350570 190938 350572
rect 191281 350570 191347 350573
rect 190932 350568 191347 350570
rect 190932 350512 191286 350568
rect 191342 350512 191347 350568
rect 190932 350510 191347 350512
rect 190932 350508 190938 350510
rect 179689 350507 179755 350508
rect 191281 350507 191347 350510
rect 196617 350570 196683 350573
rect 338481 350572 338547 350573
rect 198958 350570 198964 350572
rect 196617 350568 198964 350570
rect 196617 350512 196622 350568
rect 196678 350512 198964 350568
rect 196617 350510 198964 350512
rect 196617 350507 196683 350510
rect 198958 350508 198964 350510
rect 199028 350508 199034 350572
rect 338430 350570 338436 350572
rect 338390 350510 338436 350570
rect 338500 350568 338547 350572
rect 338542 350512 338547 350568
rect 338430 350508 338436 350510
rect 338500 350508 338547 350512
rect 339718 350508 339724 350572
rect 339788 350570 339794 350572
rect 340505 350570 340571 350573
rect 339788 350568 340571 350570
rect 339788 350512 340510 350568
rect 340566 350512 340571 350568
rect 339788 350510 340571 350512
rect 339788 350508 339794 350510
rect 338481 350507 338547 350508
rect 340505 350507 340571 350510
rect 350942 350508 350948 350572
rect 351012 350570 351018 350572
rect 351637 350570 351703 350573
rect 351012 350568 351703 350570
rect 351012 350512 351642 350568
rect 351698 350512 351703 350568
rect 351012 350510 351703 350512
rect 351012 350508 351018 350510
rect 351637 350507 351703 350510
rect 498510 350508 498516 350572
rect 498580 350570 498586 350572
rect 499021 350570 499087 350573
rect 498580 350568 499087 350570
rect 498580 350512 499026 350568
rect 499082 350512 499087 350568
rect 498580 350510 499087 350512
rect 498580 350508 498586 350510
rect 499021 350507 499087 350510
rect 499798 350508 499804 350572
rect 499868 350570 499874 350572
rect 500585 350570 500651 350573
rect 510889 350572 510955 350573
rect 510838 350570 510844 350572
rect 499868 350568 500651 350570
rect 499868 350512 500590 350568
rect 500646 350512 500651 350568
rect 499868 350510 500651 350512
rect 510798 350510 510844 350570
rect 510908 350568 510955 350572
rect 510950 350512 510955 350568
rect 499868 350508 499874 350510
rect 500585 350507 500651 350510
rect 510838 350508 510844 350510
rect 510908 350508 510955 350512
rect 510889 350507 510955 350508
rect 218329 350434 218395 350437
rect 218830 350434 218836 350436
rect 218329 350432 218836 350434
rect 218329 350376 218334 350432
rect 218390 350376 218836 350432
rect 218329 350374 218836 350376
rect 218329 350371 218395 350374
rect 218830 350372 218836 350374
rect 218900 350372 218906 350436
rect 377254 349692 377260 349756
rect 377324 349754 377330 349756
rect 380985 349754 381051 349757
rect 377324 349752 381051 349754
rect 377324 349696 380990 349752
rect 381046 349696 381051 349752
rect 377324 349694 381051 349696
rect 377324 349692 377330 349694
rect 380985 349691 381051 349694
rect -960 345524 480 345764
rect 196558 344178 196618 344190
rect 198825 344178 198891 344181
rect 196558 344176 198891 344178
rect 196558 344120 198830 344176
rect 198886 344120 198891 344176
rect 196558 344118 198891 344120
rect 356562 344178 356622 344190
rect 358905 344178 358971 344181
rect 356562 344176 358971 344178
rect 356562 344120 358910 344176
rect 358966 344120 358971 344176
rect 356562 344118 358971 344120
rect 198825 344115 198891 344118
rect 358905 344115 358971 344118
rect 516558 343770 516618 344190
rect 518985 343770 519051 343773
rect 516558 343768 519051 343770
rect 516558 343712 518990 343768
rect 519046 343712 519051 343768
rect 516558 343710 519051 343712
rect 518985 343707 519051 343710
rect 580165 339146 580231 339149
rect 583520 339146 584960 339236
rect 580165 339144 584960 339146
rect 580165 339088 580170 339144
rect 580226 339088 584960 339144
rect 580165 339086 584960 339088
rect 580165 339083 580231 339086
rect 583520 338996 584960 339086
rect -960 333012 480 333252
rect 583520 326212 584960 326452
rect -960 320514 480 320604
rect -960 320454 6930 320514
rect -960 320364 480 320454
rect 6870 320242 6930 320454
rect 54334 320242 54340 320244
rect 6870 320182 54340 320242
rect 54334 320180 54340 320182
rect 54404 320180 54410 320244
rect 52913 319970 52979 319973
rect 57094 319970 57100 319972
rect 52913 319968 57100 319970
rect 52913 319912 52918 319968
rect 52974 319912 57100 319968
rect 52913 319910 57100 319912
rect 52913 319907 52979 319910
rect 57094 319908 57100 319910
rect 57164 319908 57170 319972
rect 580901 313578 580967 313581
rect 583520 313578 584960 313668
rect 580901 313576 584960 313578
rect 580901 313520 580906 313576
rect 580962 313520 584960 313576
rect 580901 313518 584960 313520
rect 580901 313515 580967 313518
rect 583520 313428 584960 313518
rect -960 308002 480 308092
rect 2773 308002 2839 308005
rect -960 308000 2839 308002
rect -960 307944 2778 308000
rect 2834 307944 2839 308000
rect -960 307942 2839 307944
rect -960 307852 480 307942
rect 2773 307939 2839 307942
rect 56777 301746 56843 301749
rect 57605 301746 57671 301749
rect 60002 301746 60062 301894
rect 217133 301882 217199 301885
rect 217869 301882 217935 301885
rect 219390 301882 220064 301924
rect 217133 301880 220064 301882
rect 217133 301824 217138 301880
rect 217194 301824 217874 301880
rect 217930 301864 220064 301880
rect 377213 301882 377279 301885
rect 377581 301882 377647 301885
rect 379470 301882 380052 301924
rect 377213 301880 380052 301882
rect 217930 301824 219450 301864
rect 217133 301822 219450 301824
rect 377213 301824 377218 301880
rect 377274 301824 377586 301880
rect 377642 301864 380052 301880
rect 377642 301824 379530 301864
rect 377213 301822 379530 301824
rect 217133 301819 217199 301822
rect 217869 301819 217935 301822
rect 377213 301819 377279 301822
rect 377581 301819 377647 301822
rect 56777 301744 60062 301746
rect 56777 301688 56782 301744
rect 56838 301688 57610 301744
rect 57666 301688 60062 301744
rect 56777 301686 60062 301688
rect 56777 301683 56843 301686
rect 57605 301683 57671 301686
rect 56593 300930 56659 300933
rect 57697 300930 57763 300933
rect 60002 300930 60062 300942
rect 56593 300928 60062 300930
rect 56593 300872 56598 300928
rect 56654 300872 57702 300928
rect 57758 300872 60062 300928
rect 56593 300870 60062 300872
rect 217685 300930 217751 300933
rect 219390 300930 220064 300972
rect 217685 300928 220064 300930
rect 217685 300872 217690 300928
rect 217746 300912 220064 300928
rect 376845 300930 376911 300933
rect 377397 300930 377463 300933
rect 379470 300930 380052 300972
rect 376845 300928 380052 300930
rect 217746 300872 219450 300912
rect 217685 300870 219450 300872
rect 376845 300872 376850 300928
rect 376906 300872 377402 300928
rect 377458 300912 380052 300928
rect 377458 300872 379530 300912
rect 376845 300870 379530 300872
rect 56593 300867 56659 300870
rect 57697 300867 57763 300870
rect 217685 300867 217751 300870
rect 376845 300867 376911 300870
rect 377397 300867 377463 300870
rect 583520 300644 584960 300884
rect 57697 299434 57763 299437
rect 57881 299434 57947 299437
rect 57697 299432 60062 299434
rect 57697 299376 57702 299432
rect 57758 299376 57886 299432
rect 57942 299376 60062 299432
rect 57697 299374 60062 299376
rect 57697 299371 57763 299374
rect 57881 299371 57947 299374
rect 60002 298766 60062 299374
rect 217777 298754 217843 298757
rect 219390 298754 220064 298796
rect 217777 298752 220064 298754
rect 217777 298696 217782 298752
rect 217838 298736 220064 298752
rect 376937 298754 377003 298757
rect 377857 298754 377923 298757
rect 379470 298754 380052 298796
rect 376937 298752 380052 298754
rect 217838 298696 219450 298736
rect 217777 298694 219450 298696
rect 376937 298696 376942 298752
rect 376998 298696 377862 298752
rect 377918 298736 380052 298752
rect 377918 298696 379530 298736
rect 376937 298694 379530 298696
rect 217777 298691 217843 298694
rect 376937 298691 377003 298694
rect 377857 298691 377923 298694
rect 216673 298074 216739 298077
rect 217317 298074 217383 298077
rect 216673 298072 219450 298074
rect 216673 298016 216678 298072
rect 216734 298016 217322 298072
rect 217378 298016 219450 298072
rect 216673 298014 219450 298016
rect 216673 298011 216739 298014
rect 217317 298011 217383 298014
rect 219390 297844 219450 298014
rect 57421 297802 57487 297805
rect 60002 297802 60062 297814
rect 57421 297800 60062 297802
rect 57421 297744 57426 297800
rect 57482 297744 60062 297800
rect 219390 297784 220064 297844
rect 377305 297802 377371 297805
rect 379470 297802 380052 297844
rect 377305 297800 380052 297802
rect 57421 297742 60062 297744
rect 377305 297744 377310 297800
rect 377366 297784 380052 297800
rect 377366 297744 379530 297784
rect 377305 297742 379530 297744
rect 57421 297739 57487 297742
rect 377305 297739 377371 297742
rect 57513 296034 57579 296037
rect 60002 296034 60062 296046
rect 57513 296032 60062 296034
rect 57513 295976 57518 296032
rect 57574 295976 60062 296032
rect 57513 295974 60062 295976
rect 216949 296034 217015 296037
rect 219390 296034 220064 296076
rect 216949 296032 220064 296034
rect 216949 295976 216954 296032
rect 217010 296016 220064 296032
rect 377949 296034 378015 296037
rect 379470 296034 380052 296076
rect 377949 296032 380052 296034
rect 217010 295976 219450 296016
rect 216949 295974 219450 295976
rect 377949 295976 377954 296032
rect 378010 296016 380052 296032
rect 378010 295976 379530 296016
rect 377949 295974 379530 295976
rect 57513 295971 57579 295974
rect 216949 295971 217015 295974
rect 377949 295971 378015 295974
rect -960 295204 480 295444
rect 216949 295354 217015 295357
rect 217501 295354 217567 295357
rect 216949 295352 217567 295354
rect 216949 295296 216954 295352
rect 217010 295296 217506 295352
rect 217562 295296 217567 295352
rect 216949 295294 217567 295296
rect 216949 295291 217015 295294
rect 217501 295291 217567 295294
rect 376753 295354 376819 295357
rect 377949 295354 378015 295357
rect 376753 295352 378015 295354
rect 376753 295296 376758 295352
rect 376814 295296 377954 295352
rect 378010 295296 378015 295352
rect 376753 295294 378015 295296
rect 376753 295291 376819 295294
rect 377949 295291 378015 295294
rect 57329 294946 57395 294949
rect 60002 294946 60062 294958
rect 57329 294944 60062 294946
rect 57329 294888 57334 294944
rect 57390 294888 60062 294944
rect 57329 294886 60062 294888
rect 216857 294946 216923 294949
rect 219390 294946 220064 294988
rect 216857 294944 220064 294946
rect 216857 294888 216862 294944
rect 216918 294928 220064 294944
rect 377673 294946 377739 294949
rect 379470 294946 380052 294988
rect 377673 294944 380052 294946
rect 216918 294888 219450 294928
rect 216857 294886 219450 294888
rect 377673 294888 377678 294944
rect 377734 294928 380052 294944
rect 377734 294888 379530 294928
rect 377673 294886 379530 294888
rect 57329 294883 57395 294886
rect 216857 294883 216923 294886
rect 377673 294883 377739 294886
rect 56685 293994 56751 293997
rect 57329 293994 57395 293997
rect 56685 293992 57395 293994
rect 56685 293936 56690 293992
rect 56746 293936 57334 293992
rect 57390 293936 57395 293992
rect 56685 293934 57395 293936
rect 56685 293931 56751 293934
rect 57329 293931 57395 293934
rect 216857 293994 216923 293997
rect 217409 293994 217475 293997
rect 216857 293992 217475 293994
rect 216857 293936 216862 293992
rect 216918 293936 217414 293992
rect 217470 293936 217475 293992
rect 216857 293934 217475 293936
rect 216857 293931 216923 293934
rect 217409 293931 217475 293934
rect 377121 293994 377187 293997
rect 377673 293994 377739 293997
rect 377121 293992 377739 293994
rect 377121 293936 377126 293992
rect 377182 293936 377678 293992
rect 377734 293936 377739 293992
rect 377121 293934 377739 293936
rect 377121 293931 377187 293934
rect 377673 293931 377739 293934
rect 57329 292634 57395 292637
rect 60002 292634 60062 293190
rect 217041 293178 217107 293181
rect 217869 293178 217935 293181
rect 219390 293178 220064 293220
rect 217041 293176 220064 293178
rect 217041 293120 217046 293176
rect 217102 293120 217874 293176
rect 217930 293160 220064 293176
rect 377765 293178 377831 293181
rect 379470 293178 380052 293220
rect 377765 293176 380052 293178
rect 217930 293120 219450 293160
rect 217041 293118 219450 293120
rect 377765 293120 377770 293176
rect 377826 293160 380052 293176
rect 377826 293120 379530 293160
rect 377765 293118 379530 293120
rect 217041 293115 217107 293118
rect 217869 293115 217935 293118
rect 377765 293115 377831 293118
rect 57329 292632 60062 292634
rect 57329 292576 57334 292632
rect 57390 292576 60062 292632
rect 57329 292574 60062 292576
rect 57329 292571 57395 292574
rect 583520 287860 584960 288100
rect 518893 284746 518959 284749
rect 519353 284746 519419 284749
rect 516558 284744 519419 284746
rect 516558 284688 518898 284744
rect 518954 284688 519358 284744
rect 519414 284688 519419 284744
rect 516558 284686 519419 284688
rect 516558 284350 516618 284686
rect 518893 284683 518959 284686
rect 519353 284683 519419 284686
rect 196558 284338 196618 284350
rect 198733 284338 198799 284341
rect 199837 284338 199903 284341
rect 196558 284336 199903 284338
rect 196558 284280 198738 284336
rect 198794 284280 199842 284336
rect 199898 284280 199903 284336
rect 196558 284278 199903 284280
rect 356562 284338 356622 284350
rect 358813 284338 358879 284341
rect 359641 284338 359707 284341
rect 356562 284336 359707 284338
rect 356562 284280 358818 284336
rect 358874 284280 359646 284336
rect 359702 284280 359707 284336
rect 356562 284278 359707 284280
rect 198733 284275 198799 284278
rect 199837 284275 199903 284278
rect 358813 284275 358879 284278
rect 359641 284275 359707 284278
rect -960 282692 480 282932
rect 196558 282706 196618 282718
rect 199285 282706 199351 282709
rect 199745 282706 199811 282709
rect 196558 282704 199811 282706
rect 196558 282648 199290 282704
rect 199346 282648 199750 282704
rect 199806 282648 199811 282704
rect 196558 282646 199811 282648
rect 199285 282643 199351 282646
rect 199745 282643 199811 282646
rect 356562 282434 356622 282718
rect 516558 282706 516618 282718
rect 519445 282706 519511 282709
rect 516558 282704 519511 282706
rect 516558 282648 519450 282704
rect 519506 282648 519511 282704
rect 516558 282646 519511 282648
rect 519445 282643 519511 282646
rect 359181 282434 359247 282437
rect 356562 282432 359247 282434
rect 356562 282376 359186 282432
rect 359242 282376 359247 282432
rect 356562 282374 359247 282376
rect 359181 282371 359247 282374
rect 359549 281482 359615 281485
rect 519077 281482 519143 281485
rect 519537 281482 519603 281485
rect 356562 281480 359615 281482
rect 356562 281424 359554 281480
rect 359610 281424 359615 281480
rect 356562 281422 359615 281424
rect 356562 281358 356622 281422
rect 359549 281419 359615 281422
rect 517102 281480 519603 281482
rect 517102 281424 519082 281480
rect 519138 281424 519542 281480
rect 519598 281424 519603 281480
rect 517102 281422 519603 281424
rect 517102 281388 517162 281422
rect 519077 281419 519143 281422
rect 519537 281419 519603 281422
rect 196558 281346 196618 281358
rect 199101 281346 199167 281349
rect 199469 281346 199535 281349
rect 196558 281344 199535 281346
rect 196558 281288 199106 281344
rect 199162 281288 199474 281344
rect 199530 281288 199535 281344
rect 516588 281328 517162 281388
rect 196558 281286 199535 281288
rect 199101 281283 199167 281286
rect 199469 281283 199535 281286
rect 198917 280122 198983 280125
rect 199653 280122 199719 280125
rect 358997 280122 359063 280125
rect 359365 280122 359431 280125
rect 196558 280120 199719 280122
rect 196558 280064 198922 280120
rect 198978 280064 199658 280120
rect 199714 280064 199719 280120
rect 196558 280062 199719 280064
rect 196558 279862 196618 280062
rect 198917 280059 198983 280062
rect 199653 280059 199719 280062
rect 356562 280120 359431 280122
rect 356562 280064 359002 280120
rect 359058 280064 359370 280120
rect 359426 280064 359431 280120
rect 356562 280062 359431 280064
rect 356562 279862 356622 280062
rect 358997 280059 359063 280062
rect 359365 280059 359431 280062
rect 516558 279850 516618 279862
rect 519169 279850 519235 279853
rect 519629 279850 519695 279853
rect 516558 279848 519695 279850
rect 516558 279792 519174 279848
rect 519230 279792 519634 279848
rect 519690 279792 519695 279848
rect 516558 279790 519695 279792
rect 519169 279787 519235 279790
rect 519629 279787 519695 279790
rect 359089 278762 359155 278765
rect 359457 278762 359523 278765
rect 356562 278760 359523 278762
rect 356562 278704 359094 278760
rect 359150 278704 359462 278760
rect 359518 278704 359523 278760
rect 356562 278702 359523 278704
rect 356562 278638 356622 278702
rect 359089 278699 359155 278702
rect 359457 278699 359523 278702
rect 196558 278626 196618 278638
rect 199009 278626 199075 278629
rect 196558 278624 199075 278626
rect 196558 278568 199014 278624
rect 199070 278568 199075 278624
rect 196558 278566 199075 278568
rect 516558 278626 516618 278638
rect 519261 278626 519327 278629
rect 516558 278624 519327 278626
rect 516558 278568 519266 278624
rect 519322 278568 519327 278624
rect 516558 278566 519327 278568
rect 199009 278563 199075 278566
rect 519261 278563 519327 278566
rect 57605 275634 57671 275637
rect 57605 275632 60062 275634
rect 57605 275576 57610 275632
rect 57666 275576 60062 275632
rect 57605 275574 60062 275576
rect 57605 275571 57671 275574
rect 60002 274966 60062 275574
rect 583520 275076 584960 275316
rect 216673 274954 216739 274957
rect 219390 274954 220064 274996
rect 216673 274952 220064 274954
rect 216673 274896 216678 274952
rect 216734 274936 220064 274952
rect 376845 274954 376911 274957
rect 379470 274954 380052 274996
rect 376845 274952 380052 274954
rect 216734 274896 219450 274936
rect 216673 274894 219450 274896
rect 376845 274896 376850 274952
rect 376906 274936 380052 274952
rect 376906 274896 379530 274936
rect 376845 274894 379530 274896
rect 216673 274891 216739 274894
rect 376845 274891 376911 274894
rect 57237 273322 57303 273325
rect 57881 273322 57947 273325
rect 59494 273322 60032 273364
rect 57237 273320 60032 273322
rect 57237 273264 57242 273320
rect 57298 273264 57886 273320
rect 57942 273304 60032 273320
rect 216673 273322 216739 273325
rect 219390 273322 220064 273364
rect 216673 273320 220064 273322
rect 57942 273264 59554 273304
rect 57237 273262 59554 273264
rect 216673 273264 216678 273320
rect 216734 273304 220064 273320
rect 376753 273322 376819 273325
rect 379470 273322 380052 273364
rect 376753 273320 380052 273322
rect 216734 273264 219450 273304
rect 216673 273262 219450 273264
rect 376753 273264 376758 273320
rect 376814 273304 380052 273320
rect 376814 273264 379530 273304
rect 376753 273262 379530 273264
rect 57237 273259 57303 273262
rect 57881 273259 57947 273262
rect 216673 273259 216739 273262
rect 376753 273259 376819 273262
rect 58985 273050 59051 273053
rect 60002 273050 60062 273062
rect 58985 273048 60062 273050
rect 58985 272992 58990 273048
rect 59046 272992 60062 273048
rect 58985 272990 60062 272992
rect 216673 273050 216739 273053
rect 219390 273050 220064 273092
rect 216673 273048 220064 273050
rect 216673 272992 216678 273048
rect 216734 273032 220064 273048
rect 376753 273050 376819 273053
rect 379470 273050 380052 273092
rect 376753 273048 380052 273050
rect 216734 272992 219450 273032
rect 216673 272990 219450 272992
rect 376753 272992 376758 273048
rect 376814 273032 380052 273048
rect 376814 272992 379530 273032
rect 376753 272990 379530 272992
rect 58985 272987 59051 272990
rect 216673 272987 216739 272990
rect 376753 272987 376819 272990
rect -960 270330 480 270420
rect -960 270270 674 270330
rect -960 270194 480 270270
rect 614 270194 674 270270
rect -960 270180 674 270194
rect 246 270134 674 270180
rect 246 269650 306 270134
rect 246 269590 6930 269650
rect 6870 269242 6930 269590
rect 53046 269242 53052 269244
rect 6870 269182 53052 269242
rect 53046 269180 53052 269182
rect 53116 269180 53122 269244
rect 250437 265028 250503 265029
rect 274173 265028 274239 265029
rect 250437 265024 250484 265028
rect 250548 265026 250554 265028
rect 250437 264968 250442 265024
rect 250437 264964 250484 264968
rect 250548 264966 250594 265026
rect 274173 265024 274220 265028
rect 274284 265026 274290 265028
rect 274173 264968 274178 265024
rect 250548 264964 250554 264966
rect 274173 264964 274220 264968
rect 274284 264966 274330 265026
rect 274284 264964 274290 264966
rect 250437 264963 250503 264964
rect 274173 264963 274239 264964
rect 58617 264890 58683 264893
rect 110965 264892 111031 264893
rect 125961 264892 126027 264893
rect 128353 264892 128419 264893
rect 93456 264890 93462 264892
rect 58617 264888 93462 264890
rect 58617 264832 58622 264888
rect 58678 264832 93462 264888
rect 58617 264830 93462 264832
rect 58617 264827 58683 264830
rect 93456 264828 93462 264830
rect 93526 264828 93532 264892
rect 110965 264888 111006 264892
rect 111070 264890 111076 264892
rect 110965 264832 110970 264888
rect 110965 264828 111006 264832
rect 111070 264830 111122 264890
rect 111070 264828 111076 264830
rect 125960 264828 125966 264892
rect 126030 264890 126036 264892
rect 128302 264890 128308 264892
rect 126030 264830 126118 264890
rect 128262 264830 128308 264890
rect 128372 264888 128419 264892
rect 128414 264832 128419 264888
rect 126030 264828 126036 264830
rect 128302 264828 128308 264830
rect 128372 264828 128419 264832
rect 110965 264827 111031 264828
rect 125961 264827 126027 264828
rect 128353 264827 128419 264828
rect 130929 264892 130995 264893
rect 133413 264892 133479 264893
rect 135897 264892 135963 264893
rect 138473 264892 138539 264893
rect 473445 264892 473511 264893
rect 130929 264888 130998 264892
rect 130929 264832 130934 264888
rect 130990 264832 130998 264888
rect 130929 264828 130998 264832
rect 131062 264890 131068 264892
rect 131062 264830 131086 264890
rect 133413 264888 133446 264892
rect 133510 264890 133516 264892
rect 135888 264890 135894 264892
rect 133413 264832 133418 264888
rect 131062 264828 131068 264830
rect 133413 264828 133446 264832
rect 133510 264830 133570 264890
rect 135806 264830 135894 264890
rect 133510 264828 133516 264830
rect 135888 264828 135894 264830
rect 135958 264828 135964 264892
rect 138472 264828 138478 264892
rect 138542 264890 138548 264892
rect 138542 264830 138630 264890
rect 138542 264828 138548 264830
rect 196750 264828 196756 264892
rect 196820 264890 196826 264892
rect 318464 264890 318470 264892
rect 196820 264830 318470 264890
rect 196820 264828 196826 264830
rect 318464 264828 318470 264830
rect 318534 264828 318540 264892
rect 359406 264828 359412 264892
rect 359476 264890 359482 264892
rect 473432 264890 473438 264892
rect 359476 264830 473186 264890
rect 473354 264830 473438 264890
rect 473502 264888 473511 264892
rect 473506 264832 473511 264888
rect 359476 264828 359482 264830
rect 130929 264827 130995 264828
rect 133413 264827 133479 264828
rect 135897 264827 135963 264828
rect 138473 264827 138539 264828
rect 140865 264756 140931 264757
rect 143533 264756 143599 264757
rect 140865 264752 140926 264756
rect 140865 264696 140870 264752
rect 140865 264692 140926 264696
rect 140990 264754 140996 264756
rect 143504 264754 143510 264756
rect 140990 264694 141022 264754
rect 143442 264694 143510 264754
rect 143574 264752 143599 264756
rect 143594 264696 143599 264752
rect 140990 264692 140996 264694
rect 143504 264692 143510 264694
rect 143574 264692 143599 264696
rect 140865 264691 140931 264692
rect 143533 264691 143599 264692
rect 145925 264756 145991 264757
rect 148501 264756 148567 264757
rect 468477 264756 468543 264757
rect 470961 264756 471027 264757
rect 145925 264752 145958 264756
rect 146022 264754 146028 264756
rect 145925 264696 145930 264752
rect 145925 264692 145958 264696
rect 146022 264694 146082 264754
rect 148501 264752 148542 264756
rect 148606 264754 148612 264756
rect 148501 264696 148506 264752
rect 146022 264692 146028 264694
rect 148501 264692 148542 264696
rect 148606 264694 148658 264754
rect 148606 264692 148612 264694
rect 196566 264692 196572 264756
rect 196636 264754 196642 264756
rect 310984 264754 310990 264756
rect 196636 264694 310990 264754
rect 196636 264692 196642 264694
rect 310984 264692 310990 264694
rect 311054 264692 311060 264756
rect 359590 264692 359596 264756
rect 359660 264754 359666 264756
rect 445960 264754 445966 264756
rect 359660 264694 445966 264754
rect 359660 264692 359666 264694
rect 445960 264692 445966 264694
rect 446030 264692 446036 264756
rect 468477 264752 468542 264756
rect 468477 264696 468482 264752
rect 468538 264696 468542 264752
rect 468477 264692 468542 264696
rect 468606 264754 468612 264756
rect 468606 264694 468634 264754
rect 470961 264752 470990 264756
rect 471054 264754 471060 264756
rect 473126 264754 473186 264830
rect 473432 264828 473438 264830
rect 473502 264828 473511 264832
rect 473445 264827 473511 264828
rect 480897 264892 480963 264893
rect 480897 264888 480918 264892
rect 480982 264890 480988 264892
rect 480897 264832 480902 264888
rect 480897 264828 480918 264832
rect 480982 264830 481054 264890
rect 480982 264828 480988 264830
rect 480897 264827 480963 264828
rect 483381 264756 483447 264757
rect 485957 264756 486023 264757
rect 478464 264754 478470 264756
rect 470961 264696 470966 264752
rect 468606 264692 468612 264694
rect 470961 264692 470990 264696
rect 471054 264694 471118 264754
rect 473126 264694 478470 264754
rect 471054 264692 471060 264694
rect 478464 264692 478470 264694
rect 478534 264692 478540 264756
rect 483360 264754 483366 264756
rect 483290 264694 483366 264754
rect 483430 264752 483447 264756
rect 485944 264754 485950 264756
rect 483442 264696 483447 264752
rect 483360 264692 483366 264694
rect 483430 264692 483447 264696
rect 485866 264694 485950 264754
rect 486014 264752 486023 264756
rect 486018 264696 486023 264752
rect 485944 264692 485950 264694
rect 486014 264692 486023 264696
rect 145925 264691 145991 264692
rect 148501 264691 148567 264692
rect 468477 264691 468543 264692
rect 470961 264691 471027 264692
rect 483381 264691 483447 264692
rect 485957 264691 486023 264692
rect 198181 264618 198247 264621
rect 291837 264618 291903 264621
rect 198181 264616 291903 264618
rect 198181 264560 198186 264616
rect 198242 264560 291842 264616
rect 291898 264560 291903 264616
rect 198181 264558 291903 264560
rect 198181 264555 198247 264558
rect 291837 264555 291903 264558
rect 293401 264620 293467 264621
rect 418429 264620 418495 264621
rect 421097 264620 421163 264621
rect 293401 264616 293446 264620
rect 293510 264618 293516 264620
rect 293401 264560 293406 264616
rect 293401 264556 293446 264560
rect 293510 264558 293558 264618
rect 418429 264616 418494 264620
rect 418429 264560 418434 264616
rect 418490 264560 418494 264616
rect 293510 264556 293516 264558
rect 418429 264556 418494 264560
rect 418558 264618 418564 264620
rect 421072 264618 421078 264620
rect 418558 264558 418586 264618
rect 421006 264558 421078 264618
rect 421142 264616 421163 264620
rect 421158 264560 421163 264616
rect 418558 264556 418564 264558
rect 421072 264556 421078 264558
rect 421142 264556 421163 264560
rect 293401 264555 293467 264556
rect 418429 264555 418495 264556
rect 421097 264555 421163 264556
rect 423489 264620 423555 264621
rect 425973 264620 426039 264621
rect 429745 264620 429811 264621
rect 475837 264620 475903 264621
rect 423489 264616 423526 264620
rect 423590 264618 423596 264620
rect 425968 264618 425974 264620
rect 423489 264560 423494 264616
rect 423489 264556 423526 264560
rect 423590 264558 423646 264618
rect 425882 264558 425974 264618
rect 423590 264556 423596 264558
rect 425968 264556 425974 264558
rect 426038 264556 426044 264620
rect 429745 264616 429782 264620
rect 429846 264618 429852 264620
rect 429745 264560 429750 264616
rect 429745 264556 429782 264560
rect 429846 264558 429902 264618
rect 475837 264616 475886 264620
rect 475950 264618 475956 264620
rect 475837 264560 475842 264616
rect 429846 264556 429852 264558
rect 475837 264556 475886 264560
rect 475950 264558 475994 264618
rect 475950 264556 475956 264558
rect 423489 264555 423555 264556
rect 425973 264555 426039 264556
rect 429745 264555 429811 264556
rect 475837 264555 475903 264556
rect 202321 264482 202387 264485
rect 300894 264482 300900 264484
rect 202321 264480 300900 264482
rect 202321 264424 202326 264480
rect 202382 264424 300900 264480
rect 202321 264422 300900 264424
rect 202321 264419 202387 264422
rect 300894 264420 300900 264422
rect 300964 264420 300970 264484
rect 211429 264346 211495 264349
rect 280797 264348 280863 264349
rect 283373 264348 283439 264349
rect 285949 264348 286015 264349
rect 288157 264348 288223 264349
rect 290917 264348 290983 264349
rect 211429 264344 277410 264346
rect 211429 264288 211434 264344
rect 211490 264288 277410 264344
rect 211429 264286 277410 264288
rect 211429 264283 211495 264286
rect 56869 264210 56935 264213
rect 60733 264210 60799 264213
rect 117998 264210 118004 264212
rect 56869 264208 118004 264210
rect 56869 264152 56874 264208
rect 56930 264152 60738 264208
rect 60794 264152 118004 264208
rect 56869 264150 118004 264152
rect 56869 264147 56935 264150
rect 60733 264147 60799 264150
rect 117998 264148 118004 264150
rect 118068 264148 118074 264212
rect 277350 264210 277410 264286
rect 280797 264344 280844 264348
rect 280908 264346 280914 264348
rect 280797 264288 280802 264344
rect 280797 264284 280844 264288
rect 280908 264286 280954 264346
rect 283373 264344 283420 264348
rect 283484 264346 283490 264348
rect 283373 264288 283378 264344
rect 280908 264284 280914 264286
rect 283373 264284 283420 264288
rect 283484 264286 283530 264346
rect 285949 264344 285996 264348
rect 286060 264346 286066 264348
rect 285949 264288 285954 264344
rect 283484 264284 283490 264286
rect 285949 264284 285996 264288
rect 286060 264286 286106 264346
rect 288157 264344 288204 264348
rect 288268 264346 288274 264348
rect 288157 264288 288162 264344
rect 286060 264284 286066 264286
rect 288157 264284 288204 264288
rect 288268 264286 288314 264346
rect 290917 264344 290964 264348
rect 291028 264346 291034 264348
rect 291837 264346 291903 264349
rect 298502 264346 298508 264348
rect 290917 264288 290922 264344
rect 288268 264284 288274 264286
rect 290917 264284 290964 264288
rect 291028 264286 291074 264346
rect 291837 264344 298508 264346
rect 291837 264288 291842 264344
rect 291898 264288 298508 264344
rect 291837 264286 298508 264288
rect 291028 264284 291034 264286
rect 280797 264283 280863 264284
rect 283373 264283 283439 264284
rect 285949 264283 286015 264284
rect 288157 264283 288223 264284
rect 290917 264283 290983 264284
rect 291837 264283 291903 264286
rect 298502 264284 298508 264286
rect 298572 264284 298578 264348
rect 295926 264210 295932 264212
rect 277350 264150 295932 264210
rect 295926 264148 295932 264150
rect 295996 264148 296002 264212
rect 51441 263666 51507 263669
rect 51758 263666 51764 263668
rect 51441 263664 51764 263666
rect 51441 263608 51446 263664
rect 51502 263608 51764 263664
rect 51441 263606 51764 263608
rect 51441 263603 51507 263606
rect 51758 263604 51764 263606
rect 51828 263604 51834 263668
rect 218421 263666 218487 263669
rect 415853 263668 415919 263669
rect 219014 263666 219020 263668
rect 218421 263664 219020 263666
rect 218421 263608 218426 263664
rect 218482 263608 219020 263664
rect 218421 263606 219020 263608
rect 218421 263603 218487 263606
rect 219014 263604 219020 263606
rect 219084 263604 219090 263668
rect 415853 263664 415900 263668
rect 415964 263666 415970 263668
rect 415853 263608 415858 263664
rect 415853 263604 415900 263608
rect 415964 263606 416010 263666
rect 415964 263604 415970 263606
rect 415853 263603 415919 263604
rect 80053 263530 80119 263533
rect 88333 263532 88399 263533
rect 89989 263532 90055 263533
rect 90725 263532 90791 263533
rect 91277 263532 91343 263533
rect 92381 263532 92447 263533
rect 80462 263530 80468 263532
rect 80053 263528 80468 263530
rect 80053 263472 80058 263528
rect 80114 263472 80468 263528
rect 80053 263470 80468 263472
rect 80053 263467 80119 263470
rect 80462 263468 80468 263470
rect 80532 263468 80538 263532
rect 88333 263528 88380 263532
rect 88444 263530 88450 263532
rect 88333 263472 88338 263528
rect 88333 263468 88380 263472
rect 88444 263470 88490 263530
rect 89989 263528 90036 263532
rect 90100 263530 90106 263532
rect 89989 263472 89994 263528
rect 88444 263468 88450 263470
rect 89989 263468 90036 263472
rect 90100 263470 90146 263530
rect 90725 263528 90772 263532
rect 90836 263530 90842 263532
rect 90725 263472 90730 263528
rect 90100 263468 90106 263470
rect 90725 263468 90772 263472
rect 90836 263470 90882 263530
rect 91277 263528 91324 263532
rect 91388 263530 91394 263532
rect 91277 263472 91282 263528
rect 90836 263468 90842 263470
rect 91277 263468 91324 263472
rect 91388 263470 91434 263530
rect 92381 263528 92428 263532
rect 92492 263530 92498 263532
rect 93577 263530 93643 263533
rect 96061 263532 96127 263533
rect 93710 263530 93716 263532
rect 92381 263472 92386 263528
rect 91388 263468 91394 263470
rect 92381 263468 92428 263472
rect 92492 263470 92538 263530
rect 93577 263528 93716 263530
rect 93577 263472 93582 263528
rect 93638 263472 93716 263528
rect 93577 263470 93716 263472
rect 92492 263468 92498 263470
rect 88333 263467 88399 263468
rect 89989 263467 90055 263468
rect 90725 263467 90791 263468
rect 91277 263467 91343 263468
rect 92381 263467 92447 263468
rect 93577 263467 93643 263470
rect 93710 263468 93716 263470
rect 93780 263468 93786 263532
rect 96061 263528 96108 263532
rect 96172 263530 96178 263532
rect 98085 263530 98151 263533
rect 101029 263532 101095 263533
rect 98494 263530 98500 263532
rect 96061 263472 96066 263528
rect 96061 263468 96108 263472
rect 96172 263470 96218 263530
rect 98085 263528 98500 263530
rect 98085 263472 98090 263528
rect 98146 263472 98500 263528
rect 98085 263470 98500 263472
rect 96172 263468 96178 263470
rect 96061 263467 96127 263468
rect 98085 263467 98151 263470
rect 98494 263468 98500 263470
rect 98564 263468 98570 263532
rect 101029 263528 101076 263532
rect 101140 263530 101146 263532
rect 101029 263472 101034 263528
rect 101029 263468 101076 263472
rect 101140 263470 101186 263530
rect 101140 263468 101146 263470
rect 103278 263468 103284 263532
rect 103348 263530 103354 263532
rect 103513 263530 103579 263533
rect 103348 263528 103579 263530
rect 103348 263472 103518 263528
rect 103574 263472 103579 263528
rect 103348 263470 103579 263472
rect 103348 263468 103354 263470
rect 101029 263467 101095 263468
rect 103513 263467 103579 263470
rect 105629 263530 105695 263533
rect 108205 263532 108271 263533
rect 105854 263530 105860 263532
rect 105629 263528 105860 263530
rect 105629 263472 105634 263528
rect 105690 263472 105860 263528
rect 105629 263470 105860 263472
rect 105629 263467 105695 263470
rect 105854 263468 105860 263470
rect 105924 263468 105930 263532
rect 108205 263528 108252 263532
rect 108316 263530 108322 263532
rect 109309 263530 109375 263533
rect 109718 263530 109724 263532
rect 108205 263472 108210 263528
rect 108205 263468 108252 263472
rect 108316 263470 108362 263530
rect 109309 263528 109724 263530
rect 109309 263472 109314 263528
rect 109370 263472 109724 263528
rect 109309 263470 109724 263472
rect 108316 263468 108322 263470
rect 108205 263467 108271 263468
rect 109309 263467 109375 263470
rect 109718 263468 109724 263470
rect 109788 263468 109794 263532
rect 113357 263530 113423 263533
rect 115933 263532 115999 263533
rect 113582 263530 113588 263532
rect 113357 263528 113588 263530
rect 113357 263472 113362 263528
rect 113418 263472 113588 263528
rect 113357 263470 113588 263472
rect 113357 263467 113423 263470
rect 113582 263468 113588 263470
rect 113652 263468 113658 263532
rect 115933 263528 115980 263532
rect 116044 263530 116050 263532
rect 116209 263530 116275 263533
rect 116894 263530 116900 263532
rect 115933 263472 115938 263528
rect 115933 263468 115980 263472
rect 116044 263470 116090 263530
rect 116209 263528 116900 263530
rect 116209 263472 116214 263528
rect 116270 263472 116900 263528
rect 116209 263470 116900 263472
rect 116044 263468 116050 263470
rect 115933 263467 115999 263468
rect 116209 263467 116275 263470
rect 116894 263468 116900 263470
rect 116964 263468 116970 263532
rect 118049 263530 118115 263533
rect 120901 263532 120967 263533
rect 123477 263532 123543 263533
rect 150985 263532 151051 263533
rect 155953 263532 156019 263533
rect 158529 263532 158595 263533
rect 118366 263530 118372 263532
rect 118049 263528 118372 263530
rect 118049 263472 118054 263528
rect 118110 263472 118372 263528
rect 118049 263470 118372 263472
rect 118049 263467 118115 263470
rect 118366 263468 118372 263470
rect 118436 263468 118442 263532
rect 120901 263528 120948 263532
rect 121012 263530 121018 263532
rect 120901 263472 120906 263528
rect 120901 263468 120948 263472
rect 121012 263470 121058 263530
rect 123477 263528 123524 263532
rect 123588 263530 123594 263532
rect 150934 263530 150940 263532
rect 123477 263472 123482 263528
rect 121012 263468 121018 263470
rect 123477 263468 123524 263472
rect 123588 263470 123634 263530
rect 150894 263470 150940 263530
rect 151004 263528 151051 263532
rect 155902 263530 155908 263532
rect 151046 263472 151051 263528
rect 123588 263468 123594 263470
rect 150934 263468 150940 263470
rect 151004 263468 151051 263472
rect 155862 263470 155908 263530
rect 155972 263528 156019 263532
rect 158478 263530 158484 263532
rect 156014 263472 156019 263528
rect 155902 263468 155908 263470
rect 155972 263468 156019 263472
rect 158438 263470 158484 263530
rect 158548 263528 158595 263532
rect 158590 263472 158595 263528
rect 158478 263468 158484 263470
rect 158548 263468 158595 263472
rect 160870 263468 160876 263532
rect 160940 263530 160946 263532
rect 161105 263530 161171 263533
rect 163497 263532 163563 263533
rect 166073 263532 166139 263533
rect 235993 263532 236059 263533
rect 163446 263530 163452 263532
rect 160940 263528 161171 263530
rect 160940 263472 161110 263528
rect 161166 263472 161171 263528
rect 160940 263470 161171 263472
rect 163406 263470 163452 263530
rect 163516 263528 163563 263532
rect 166022 263530 166028 263532
rect 163558 263472 163563 263528
rect 160940 263468 160946 263470
rect 120901 263467 120967 263468
rect 123477 263467 123543 263468
rect 150985 263467 151051 263468
rect 155953 263467 156019 263468
rect 158529 263467 158595 263468
rect 161105 263467 161171 263470
rect 163446 263468 163452 263470
rect 163516 263468 163563 263472
rect 165982 263470 166028 263530
rect 166092 263528 166139 263532
rect 235942 263530 235948 263532
rect 166134 263472 166139 263528
rect 166022 263468 166028 263470
rect 166092 263468 166139 263472
rect 235902 263470 235948 263530
rect 236012 263528 236059 263532
rect 236054 263472 236059 263528
rect 235942 263468 235948 263470
rect 236012 263468 236059 263472
rect 163497 263467 163563 263468
rect 166073 263467 166139 263468
rect 235993 263467 236059 263468
rect 238753 263530 238819 263533
rect 243077 263532 243143 263533
rect 239622 263530 239628 263532
rect 238753 263528 239628 263530
rect 238753 263472 238758 263528
rect 238814 263472 239628 263528
rect 238753 263470 239628 263472
rect 238753 263467 238819 263470
rect 239622 263468 239628 263470
rect 239692 263468 239698 263532
rect 243077 263528 243124 263532
rect 243188 263530 243194 263532
rect 247125 263530 247191 263533
rect 247534 263530 247540 263532
rect 243077 263472 243082 263528
rect 243077 263468 243124 263472
rect 243188 263470 243234 263530
rect 247125 263528 247540 263530
rect 247125 263472 247130 263528
rect 247186 263472 247540 263528
rect 247125 263470 247540 263472
rect 243188 263468 243194 263470
rect 243077 263467 243143 263468
rect 247125 263467 247191 263470
rect 247534 263468 247540 263470
rect 247604 263468 247610 263532
rect 247677 263530 247743 263533
rect 253565 263532 253631 263533
rect 256141 263532 256207 263533
rect 258165 263532 258231 263533
rect 248270 263530 248276 263532
rect 247677 263528 248276 263530
rect 247677 263472 247682 263528
rect 247738 263472 248276 263528
rect 247677 263470 248276 263472
rect 247677 263467 247743 263470
rect 248270 263468 248276 263470
rect 248340 263468 248346 263532
rect 253565 263528 253612 263532
rect 253676 263530 253682 263532
rect 253565 263472 253570 263528
rect 253565 263468 253612 263472
rect 253676 263470 253722 263530
rect 256141 263528 256188 263532
rect 256252 263530 256258 263532
rect 256141 263472 256146 263528
rect 253676 263468 253682 263470
rect 256141 263468 256188 263472
rect 256252 263470 256298 263530
rect 258165 263528 258212 263532
rect 258276 263530 258282 263532
rect 260833 263530 260899 263533
rect 261702 263530 261708 263532
rect 258165 263472 258170 263528
rect 256252 263468 256258 263470
rect 258165 263468 258212 263472
rect 258276 263470 258322 263530
rect 260833 263528 261708 263530
rect 260833 263472 260838 263528
rect 260894 263472 261708 263528
rect 260833 263470 261708 263472
rect 258276 263468 258282 263470
rect 253565 263467 253631 263468
rect 256141 263467 256207 263468
rect 258165 263467 258231 263468
rect 260833 263467 260899 263470
rect 261702 263468 261708 263470
rect 261772 263468 261778 263532
rect 262213 263530 262279 263533
rect 263593 263532 263659 263533
rect 262806 263530 262812 263532
rect 262213 263528 262812 263530
rect 262213 263472 262218 263528
rect 262274 263472 262812 263528
rect 262213 263470 262812 263472
rect 262213 263467 262279 263470
rect 262806 263468 262812 263470
rect 262876 263468 262882 263532
rect 263542 263530 263548 263532
rect 263502 263470 263548 263530
rect 263612 263528 263659 263532
rect 263654 263472 263659 263528
rect 263542 263468 263548 263470
rect 263612 263468 263659 263472
rect 263593 263467 263659 263468
rect 264973 263530 265039 263533
rect 265893 263532 265959 263533
rect 268285 263532 268351 263533
rect 269757 263532 269823 263533
rect 270861 263532 270927 263533
rect 271229 263532 271295 263533
rect 265198 263530 265204 263532
rect 264973 263528 265204 263530
rect 264973 263472 264978 263528
rect 265034 263472 265204 263528
rect 264973 263470 265204 263472
rect 264973 263467 265039 263470
rect 265198 263468 265204 263470
rect 265268 263468 265274 263532
rect 265893 263528 265940 263532
rect 266004 263530 266010 263532
rect 265893 263472 265898 263528
rect 265893 263468 265940 263472
rect 266004 263470 266050 263530
rect 268285 263528 268332 263532
rect 268396 263530 268402 263532
rect 268285 263472 268290 263528
rect 266004 263468 266010 263470
rect 268285 263468 268332 263472
rect 268396 263470 268442 263530
rect 269757 263528 269804 263532
rect 269868 263530 269874 263532
rect 269757 263472 269762 263528
rect 268396 263468 268402 263470
rect 269757 263468 269804 263472
rect 269868 263470 269914 263530
rect 270861 263528 270908 263532
rect 270972 263530 270978 263532
rect 270861 263472 270866 263528
rect 269868 263468 269874 263470
rect 270861 263468 270908 263472
rect 270972 263470 271018 263530
rect 271229 263528 271276 263532
rect 271340 263530 271346 263532
rect 272057 263530 272123 263533
rect 273253 263532 273319 263533
rect 275921 263532 275987 263533
rect 276105 263532 276171 263533
rect 279233 263532 279299 263533
rect 272190 263530 272196 263532
rect 271229 263472 271234 263528
rect 270972 263468 270978 263470
rect 271229 263468 271276 263472
rect 271340 263470 271386 263530
rect 272057 263528 272196 263530
rect 272057 263472 272062 263528
rect 272118 263472 272196 263528
rect 272057 263470 272196 263472
rect 271340 263468 271346 263470
rect 265893 263467 265959 263468
rect 268285 263467 268351 263468
rect 269757 263467 269823 263468
rect 270861 263467 270927 263468
rect 271229 263467 271295 263468
rect 272057 263467 272123 263470
rect 272190 263468 272196 263470
rect 272260 263468 272266 263532
rect 273253 263528 273300 263532
rect 273364 263530 273370 263532
rect 275870 263530 275876 263532
rect 273253 263472 273258 263528
rect 273253 263468 273300 263472
rect 273364 263470 273410 263530
rect 275830 263470 275876 263530
rect 275940 263528 275987 263532
rect 275982 263472 275987 263528
rect 273364 263468 273370 263470
rect 275870 263468 275876 263470
rect 275940 263468 275987 263472
rect 276054 263468 276060 263532
rect 276124 263530 276171 263532
rect 279182 263530 279188 263532
rect 276124 263528 276216 263530
rect 276166 263472 276216 263528
rect 276124 263470 276216 263472
rect 279142 263470 279188 263530
rect 279252 263528 279299 263532
rect 279294 263472 279299 263528
rect 276124 263468 276171 263470
rect 279182 263468 279188 263470
rect 279252 263468 279299 263472
rect 273253 263467 273319 263468
rect 275921 263467 275987 263468
rect 276105 263467 276171 263468
rect 279233 263467 279299 263468
rect 305821 263532 305887 263533
rect 308397 263532 308463 263533
rect 305821 263528 305868 263532
rect 305932 263530 305938 263532
rect 305821 263472 305826 263528
rect 305821 263468 305868 263472
rect 305932 263470 305978 263530
rect 308397 263528 308444 263532
rect 308508 263530 308514 263532
rect 323025 263530 323091 263533
rect 323342 263530 323348 263532
rect 308397 263472 308402 263528
rect 305932 263468 305938 263470
rect 308397 263468 308444 263472
rect 308508 263470 308554 263530
rect 323025 263528 323348 263530
rect 323025 263472 323030 263528
rect 323086 263472 323348 263528
rect 323025 263470 323348 263472
rect 308508 263468 308514 263470
rect 305821 263467 305887 263468
rect 308397 263467 308463 263468
rect 323025 263467 323091 263470
rect 323342 263468 323348 263470
rect 323412 263468 323418 263532
rect 325785 263530 325851 263533
rect 325918 263530 325924 263532
rect 325785 263528 325924 263530
rect 325785 263472 325790 263528
rect 325846 263472 325924 263528
rect 325785 263470 325924 263472
rect 325785 263467 325851 263470
rect 325918 263468 325924 263470
rect 325988 263468 325994 263532
rect 343214 263468 343220 263532
rect 343284 263530 343290 263532
rect 343449 263530 343515 263533
rect 343284 263528 343515 263530
rect 343284 263472 343454 263528
rect 343510 263472 343515 263528
rect 343284 263470 343515 263472
rect 343284 263468 343290 263470
rect 343449 263467 343515 263470
rect 397453 263530 397519 263533
rect 398230 263530 398236 263532
rect 397453 263528 398236 263530
rect 397453 263472 397458 263528
rect 397514 263472 398236 263528
rect 397453 263470 398236 263472
rect 397453 263467 397519 263470
rect 398230 263468 398236 263470
rect 398300 263468 398306 263532
rect 401593 263530 401659 263533
rect 401726 263530 401732 263532
rect 401593 263528 401732 263530
rect 401593 263472 401598 263528
rect 401654 263472 401732 263528
rect 401593 263470 401732 263472
rect 401593 263467 401659 263470
rect 401726 263468 401732 263470
rect 401796 263468 401802 263532
rect 404353 263530 404419 263533
rect 408309 263532 408375 263533
rect 410701 263532 410767 263533
rect 413645 263532 413711 263533
rect 405406 263530 405412 263532
rect 404353 263528 405412 263530
rect 404353 263472 404358 263528
rect 404414 263472 405412 263528
rect 404353 263470 405412 263472
rect 404353 263467 404419 263470
rect 405406 263468 405412 263470
rect 405476 263468 405482 263532
rect 408309 263528 408356 263532
rect 408420 263530 408426 263532
rect 408309 263472 408314 263528
rect 408309 263468 408356 263472
rect 408420 263470 408466 263530
rect 410701 263528 410748 263532
rect 410812 263530 410818 263532
rect 410701 263472 410706 263528
rect 408420 263468 408426 263470
rect 410701 263468 410748 263472
rect 410812 263470 410858 263530
rect 413645 263528 413692 263532
rect 413756 263530 413762 263532
rect 415761 263530 415827 263533
rect 419349 263532 419415 263533
rect 425237 263532 425303 263533
rect 426433 263532 426499 263533
rect 416078 263530 416084 263532
rect 413645 263472 413650 263528
rect 410812 263468 410818 263470
rect 413645 263468 413692 263472
rect 413756 263470 413802 263530
rect 415761 263528 416084 263530
rect 415761 263472 415766 263528
rect 415822 263472 416084 263528
rect 415761 263470 416084 263472
rect 413756 263468 413762 263470
rect 408309 263467 408375 263468
rect 410701 263467 410767 263468
rect 413645 263467 413711 263468
rect 415761 263467 415827 263470
rect 416078 263468 416084 263470
rect 416148 263468 416154 263532
rect 419349 263528 419396 263532
rect 419460 263530 419466 263532
rect 419349 263472 419354 263528
rect 419349 263468 419396 263472
rect 419460 263470 419506 263530
rect 425237 263528 425284 263532
rect 425348 263530 425354 263532
rect 426382 263530 426388 263532
rect 425237 263472 425242 263528
rect 419460 263468 419466 263470
rect 425237 263468 425284 263472
rect 425348 263470 425394 263530
rect 426342 263470 426388 263530
rect 426452 263528 426499 263532
rect 426494 263472 426499 263528
rect 425348 263468 425354 263470
rect 426382 263468 426388 263470
rect 426452 263468 426499 263472
rect 419349 263467 419415 263468
rect 425237 263467 425303 263468
rect 426433 263467 426499 263468
rect 427445 263532 427511 263533
rect 428181 263532 428247 263533
rect 430941 263532 431007 263533
rect 432229 263532 432295 263533
rect 433333 263532 433399 263533
rect 427445 263528 427492 263532
rect 427556 263530 427562 263532
rect 427445 263472 427450 263528
rect 427445 263468 427492 263472
rect 427556 263470 427602 263530
rect 428181 263528 428228 263532
rect 428292 263530 428298 263532
rect 428181 263472 428186 263528
rect 427556 263468 427562 263470
rect 428181 263468 428228 263472
rect 428292 263470 428338 263530
rect 430941 263528 430988 263532
rect 431052 263530 431058 263532
rect 430941 263472 430946 263528
rect 428292 263468 428298 263470
rect 430941 263468 430988 263472
rect 431052 263470 431098 263530
rect 432229 263528 432276 263532
rect 432340 263530 432346 263532
rect 432229 263472 432234 263528
rect 431052 263468 431058 263470
rect 432229 263468 432276 263472
rect 432340 263470 432386 263530
rect 433333 263528 433380 263532
rect 433444 263530 433450 263532
rect 433333 263472 433338 263528
rect 432340 263468 432346 263470
rect 433333 263468 433380 263472
rect 433444 263470 433490 263530
rect 433444 263468 433450 263470
rect 434478 263468 434484 263532
rect 434548 263530 434554 263532
rect 434621 263530 434687 263533
rect 434548 263528 434687 263530
rect 434548 263472 434626 263528
rect 434682 263472 434687 263528
rect 434548 263470 434687 263472
rect 434548 263468 434554 263470
rect 427445 263467 427511 263468
rect 428181 263467 428247 263468
rect 430941 263467 431007 263468
rect 432229 263467 432295 263468
rect 433333 263467 433399 263468
rect 434621 263467 434687 263470
rect 435909 263532 435975 263533
rect 435909 263528 435956 263532
rect 436020 263530 436026 263532
rect 435909 263472 435914 263528
rect 435909 263468 435956 263472
rect 436020 263470 436066 263530
rect 436020 263468 436026 263470
rect 438158 263468 438164 263532
rect 438228 263530 438234 263532
rect 438761 263530 438827 263533
rect 438228 263528 438827 263530
rect 438228 263472 438766 263528
rect 438822 263472 438827 263528
rect 438228 263470 438827 263472
rect 438228 263468 438234 263470
rect 435909 263467 435975 263468
rect 438761 263467 438827 263470
rect 440877 263532 440943 263533
rect 443453 263532 443519 263533
rect 448237 263532 448303 263533
rect 450997 263532 451063 263533
rect 453389 263532 453455 263533
rect 455781 263532 455847 263533
rect 503529 263532 503595 263533
rect 440877 263528 440924 263532
rect 440988 263530 440994 263532
rect 440877 263472 440882 263528
rect 440877 263468 440924 263472
rect 440988 263470 441034 263530
rect 443453 263528 443500 263532
rect 443564 263530 443570 263532
rect 443453 263472 443458 263528
rect 440988 263468 440994 263470
rect 443453 263468 443500 263472
rect 443564 263470 443610 263530
rect 448237 263528 448284 263532
rect 448348 263530 448354 263532
rect 448237 263472 448242 263528
rect 443564 263468 443570 263470
rect 448237 263468 448284 263472
rect 448348 263470 448394 263530
rect 450997 263528 451044 263532
rect 451108 263530 451114 263532
rect 450997 263472 451002 263528
rect 448348 263468 448354 263470
rect 450997 263468 451044 263472
rect 451108 263470 451154 263530
rect 453389 263528 453436 263532
rect 453500 263530 453506 263532
rect 453389 263472 453394 263528
rect 451108 263468 451114 263470
rect 453389 263468 453436 263472
rect 453500 263470 453546 263530
rect 455781 263528 455828 263532
rect 455892 263530 455898 263532
rect 503478 263530 503484 263532
rect 455781 263472 455786 263528
rect 453500 263468 453506 263470
rect 455781 263468 455828 263472
rect 455892 263470 455938 263530
rect 503438 263470 503484 263530
rect 503548 263528 503595 263532
rect 503590 263472 503595 263528
rect 455892 263468 455898 263470
rect 503478 263468 503484 263470
rect 503548 263468 503595 263472
rect 440877 263467 440943 263468
rect 443453 263467 443519 263468
rect 448237 263467 448303 263468
rect 450997 263467 451063 263468
rect 453389 263467 453455 263468
rect 455781 263467 455847 263468
rect 503529 263467 503595 263468
rect 48957 263394 49023 263397
rect 83038 263394 83044 263396
rect 48957 263392 83044 263394
rect 48957 263336 48962 263392
rect 49018 263336 83044 263392
rect 48957 263334 83044 263336
rect 48957 263331 49023 263334
rect 83038 263332 83044 263334
rect 83108 263332 83114 263396
rect 113398 263332 113404 263396
rect 113468 263394 113474 263396
rect 114369 263394 114435 263397
rect 113468 263392 114435 263394
rect 113468 263336 114374 263392
rect 114430 263336 114435 263392
rect 113468 263334 114435 263336
rect 113468 263332 113474 263334
rect 114369 263331 114435 263334
rect 153510 263332 153516 263396
rect 153580 263394 153586 263396
rect 198774 263394 198780 263396
rect 153580 263334 198780 263394
rect 153580 263332 153586 263334
rect 198774 263332 198780 263334
rect 198844 263332 198850 263396
rect 213453 263394 213519 263397
rect 320950 263394 320956 263396
rect 213453 263392 320956 263394
rect 213453 263336 213458 263392
rect 213514 263336 320956 263392
rect 213453 263334 320956 263336
rect 213453 263331 213519 263334
rect 320950 263332 320956 263334
rect 321020 263332 321026 263396
rect 373441 263394 373507 263397
rect 463550 263394 463556 263396
rect 373441 263392 463556 263394
rect 373441 263336 373446 263392
rect 373502 263336 463556 263392
rect 373441 263334 463556 263336
rect 373441 263331 373507 263334
rect 463550 263332 463556 263334
rect 463620 263332 463626 263396
rect 46565 263258 46631 263261
rect 77150 263258 77156 263260
rect 46565 263256 77156 263258
rect 46565 263200 46570 263256
rect 46626 263200 77156 263256
rect 46565 263198 77156 263200
rect 46565 263195 46631 263198
rect 77150 263196 77156 263198
rect 77220 263196 77226 263260
rect 81433 263258 81499 263261
rect 81750 263258 81756 263260
rect 81433 263256 81756 263258
rect 81433 263200 81438 263256
rect 81494 263200 81756 263256
rect 81433 263198 81756 263200
rect 81433 263195 81499 263198
rect 81750 263196 81756 263198
rect 81820 263196 81826 263260
rect 84745 263258 84811 263261
rect 85430 263258 85436 263260
rect 84745 263256 85436 263258
rect 84745 263200 84750 263256
rect 84806 263200 85436 263256
rect 84745 263198 85436 263200
rect 84745 263195 84811 263198
rect 85430 263196 85436 263198
rect 85500 263196 85506 263260
rect 95918 263196 95924 263260
rect 95988 263258 95994 263260
rect 96521 263258 96587 263261
rect 99465 263260 99531 263261
rect 99414 263258 99420 263260
rect 95988 263256 96587 263258
rect 95988 263200 96526 263256
rect 96582 263200 96587 263256
rect 95988 263198 96587 263200
rect 99374 263198 99420 263258
rect 99484 263256 99531 263260
rect 99526 263200 99531 263256
rect 95988 263196 95994 263198
rect 96521 263195 96587 263198
rect 99414 263196 99420 263198
rect 99484 263196 99531 263200
rect 99465 263195 99531 263196
rect 213269 263258 213335 263261
rect 313406 263258 313412 263260
rect 213269 263256 313412 263258
rect 213269 263200 213274 263256
rect 213330 263200 313412 263256
rect 213269 263198 313412 263200
rect 213269 263195 213335 263198
rect 313406 263196 313412 263198
rect 313476 263196 313482 263260
rect 315798 263196 315804 263260
rect 315868 263196 315874 263260
rect 379237 263258 379303 263261
rect 465942 263258 465948 263260
rect 379237 263256 465948 263258
rect 379237 263200 379242 263256
rect 379298 263200 465948 263256
rect 379237 263198 465948 263200
rect 48221 263122 48287 263125
rect 76046 263122 76052 263124
rect 48221 263120 76052 263122
rect 48221 263064 48226 263120
rect 48282 263064 76052 263120
rect 48221 263062 76052 263064
rect 48221 263059 48287 263062
rect 76046 263060 76052 263062
rect 76116 263060 76122 263124
rect 82077 263122 82143 263125
rect 103830 263122 103836 263124
rect 82077 263120 103836 263122
rect 82077 263064 82082 263120
rect 82138 263064 103836 263120
rect 82077 263062 103836 263064
rect 82077 263059 82143 263062
rect 103830 263060 103836 263062
rect 103900 263060 103906 263124
rect 217174 263060 217180 263124
rect 217244 263122 217250 263124
rect 278446 263122 278452 263124
rect 217244 263062 278452 263122
rect 217244 263060 217250 263062
rect 278446 263060 278452 263062
rect 278516 263060 278522 263124
rect 315806 263122 315866 263196
rect 379237 263195 379303 263198
rect 465942 263196 465948 263198
rect 466012 263196 466018 263260
rect 296670 263062 315866 263122
rect 83958 262924 83964 262988
rect 84028 262986 84034 262988
rect 84193 262986 84259 262989
rect 84028 262984 84259 262986
rect 84028 262928 84198 262984
rect 84254 262928 84259 262984
rect 84028 262926 84259 262928
rect 84028 262924 84034 262926
rect 84193 262923 84259 262926
rect 87597 262988 87663 262989
rect 87597 262984 87644 262988
rect 87708 262986 87714 262988
rect 88609 262986 88675 262989
rect 100753 262988 100819 262989
rect 88742 262986 88748 262988
rect 87597 262928 87602 262984
rect 87597 262924 87644 262928
rect 87708 262926 87754 262986
rect 88609 262984 88748 262986
rect 88609 262928 88614 262984
rect 88670 262928 88748 262984
rect 88609 262926 88748 262928
rect 87708 262924 87714 262926
rect 87597 262923 87663 262924
rect 88609 262923 88675 262926
rect 88742 262924 88748 262926
rect 88812 262924 88818 262988
rect 100702 262986 100708 262988
rect 100662 262926 100708 262986
rect 100772 262984 100819 262988
rect 100814 262928 100819 262984
rect 100702 262924 100708 262926
rect 100772 262924 100819 262928
rect 100753 262923 100819 262924
rect 118693 262986 118759 262989
rect 119102 262986 119108 262988
rect 118693 262984 119108 262986
rect 118693 262928 118698 262984
rect 118754 262928 119108 262984
rect 118693 262926 119108 262928
rect 118693 262923 118759 262926
rect 119102 262924 119108 262926
rect 119172 262924 119178 262988
rect 215753 262986 215819 262989
rect 216489 262986 216555 262989
rect 237046 262986 237052 262988
rect 215753 262984 237052 262986
rect 215753 262928 215758 262984
rect 215814 262928 216494 262984
rect 216550 262928 237052 262984
rect 215753 262926 237052 262928
rect 215753 262923 215819 262926
rect 216489 262923 216555 262926
rect 237046 262924 237052 262926
rect 237116 262924 237122 262988
rect 244222 262924 244228 262988
rect 244292 262986 244298 262988
rect 244365 262986 244431 262989
rect 244292 262984 244431 262986
rect 244292 262928 244370 262984
rect 244426 262928 244431 262984
rect 244292 262926 244431 262928
rect 244292 262924 244298 262926
rect 244365 262923 244431 262926
rect 258349 262988 258415 262989
rect 260925 262988 260991 262989
rect 258349 262984 258396 262988
rect 258460 262986 258466 262988
rect 258349 262928 258354 262984
rect 258349 262924 258396 262928
rect 258460 262926 258506 262986
rect 260925 262984 260972 262988
rect 261036 262986 261042 262988
rect 273345 262986 273411 262989
rect 273478 262986 273484 262988
rect 260925 262928 260930 262984
rect 258460 262924 258466 262926
rect 260925 262924 260972 262928
rect 261036 262926 261082 262986
rect 273345 262984 273484 262986
rect 273345 262928 273350 262984
rect 273406 262928 273484 262984
rect 273345 262926 273484 262928
rect 261036 262924 261042 262926
rect 258349 262923 258415 262924
rect 260925 262923 260991 262924
rect 273345 262923 273411 262926
rect 273478 262924 273484 262926
rect 273548 262924 273554 262988
rect 49049 262850 49115 262853
rect 66253 262850 66319 262853
rect 49049 262848 66319 262850
rect 49049 262792 49054 262848
rect 49110 262792 66258 262848
rect 66314 262792 66319 262848
rect 49049 262790 66319 262792
rect 49049 262787 49115 262790
rect 66253 262787 66319 262790
rect 78673 262850 78739 262853
rect 79542 262850 79548 262852
rect 78673 262848 79548 262850
rect 78673 262792 78678 262848
rect 78734 262792 79548 262848
rect 78673 262790 79548 262792
rect 78673 262787 78739 262790
rect 79542 262788 79548 262790
rect 79612 262788 79618 262852
rect 80145 262850 80211 262853
rect 112110 262850 112116 262852
rect 80145 262848 112116 262850
rect 80145 262792 80150 262848
rect 80206 262792 112116 262848
rect 80145 262790 112116 262792
rect 80145 262787 80211 262790
rect 112110 262788 112116 262790
rect 112180 262788 112186 262852
rect 59813 262714 59879 262717
rect 101765 262716 101831 262717
rect 94446 262714 94452 262716
rect 59813 262712 94452 262714
rect 59813 262656 59818 262712
rect 59874 262656 94452 262712
rect 59813 262654 94452 262656
rect 59813 262651 59879 262654
rect 94446 262652 94452 262654
rect 94516 262652 94522 262716
rect 101765 262712 101812 262716
rect 101876 262714 101882 262716
rect 102317 262714 102383 262717
rect 102726 262714 102732 262716
rect 101765 262656 101770 262712
rect 101765 262652 101812 262656
rect 101876 262654 101922 262714
rect 102317 262712 102732 262714
rect 102317 262656 102322 262712
rect 102378 262656 102732 262712
rect 102317 262654 102732 262656
rect 101876 262652 101882 262654
rect 101765 262651 101831 262652
rect 102317 262651 102383 262654
rect 102726 262652 102732 262654
rect 102796 262652 102802 262716
rect 105077 262714 105143 262717
rect 105302 262714 105308 262716
rect 105077 262712 105308 262714
rect 105077 262656 105082 262712
rect 105138 262656 105308 262712
rect 105077 262654 105308 262656
rect 105077 262651 105143 262654
rect 105302 262652 105308 262654
rect 105372 262652 105378 262716
rect 108021 262714 108087 262717
rect 108614 262714 108620 262716
rect 108021 262712 108620 262714
rect 108021 262656 108026 262712
rect 108082 262656 108620 262712
rect 108021 262654 108620 262656
rect 108021 262651 108087 262654
rect 108614 262652 108620 262654
rect 108684 262652 108690 262716
rect 205265 262714 205331 262717
rect 296670 262714 296730 263062
rect 343398 263060 343404 263124
rect 343468 263122 343474 263124
rect 343541 263122 343607 263125
rect 343468 263120 343607 263122
rect 343468 263064 343546 263120
rect 343602 263064 343607 263120
rect 343468 263062 343607 263064
rect 343468 263060 343474 263062
rect 343541 263059 343607 263062
rect 376385 263122 376451 263125
rect 460974 263122 460980 263124
rect 376385 263120 460980 263122
rect 376385 263064 376390 263120
rect 376446 263064 460980 263120
rect 376385 263062 460980 263064
rect 376385 263059 376451 263062
rect 460974 263060 460980 263062
rect 461044 263060 461050 263124
rect 378174 262924 378180 262988
rect 378244 262986 378250 262988
rect 378501 262986 378567 262989
rect 378244 262984 378567 262986
rect 378244 262928 378506 262984
rect 378562 262928 378567 262984
rect 378244 262926 378567 262928
rect 378244 262924 378250 262926
rect 378501 262923 378567 262926
rect 419809 262986 419875 262989
rect 421741 262988 421807 262989
rect 433517 262988 433583 262989
rect 420678 262986 420684 262988
rect 419809 262984 420684 262986
rect 419809 262928 419814 262984
rect 419870 262928 420684 262984
rect 419809 262926 420684 262928
rect 419809 262923 419875 262926
rect 420678 262924 420684 262926
rect 420748 262924 420754 262988
rect 421741 262984 421788 262988
rect 421852 262986 421858 262988
rect 421741 262928 421746 262984
rect 421741 262924 421788 262928
rect 421852 262926 421898 262986
rect 433517 262984 433564 262988
rect 433628 262986 433634 262988
rect 435173 262986 435239 262989
rect 435766 262986 435772 262988
rect 433517 262928 433522 262984
rect 421852 262924 421858 262926
rect 433517 262924 433564 262928
rect 433628 262926 433674 262986
rect 435173 262984 435772 262986
rect 435173 262928 435178 262984
rect 435234 262928 435772 262984
rect 435173 262926 435772 262928
rect 433628 262924 433634 262926
rect 421741 262923 421807 262924
rect 433517 262923 433583 262924
rect 435173 262923 435239 262926
rect 435766 262924 435772 262926
rect 435836 262924 435842 262988
rect 438393 262986 438459 262989
rect 438526 262986 438532 262988
rect 438393 262984 438532 262986
rect 438393 262928 438398 262984
rect 438454 262928 438532 262984
rect 438393 262926 438532 262928
rect 438393 262923 438459 262926
rect 438526 262924 438532 262926
rect 438596 262924 438602 262988
rect 396073 262850 396139 262853
rect 397126 262850 397132 262852
rect 396073 262848 397132 262850
rect 396073 262792 396078 262848
rect 396134 262792 397132 262848
rect 396073 262790 397132 262792
rect 396073 262787 396139 262790
rect 397126 262788 397132 262790
rect 397196 262788 397202 262852
rect 412725 262850 412791 262853
rect 418153 262852 418219 262853
rect 413318 262850 413324 262852
rect 412725 262848 413324 262850
rect 412725 262792 412730 262848
rect 412786 262792 413324 262848
rect 412725 262790 413324 262792
rect 412725 262787 412791 262790
rect 413318 262788 413324 262790
rect 413388 262788 413394 262852
rect 418102 262850 418108 262852
rect 418062 262790 418108 262850
rect 418172 262848 418219 262852
rect 418214 262792 418219 262848
rect 418102 262788 418108 262790
rect 418172 262788 418219 262792
rect 418153 262787 418219 262788
rect 205265 262712 296730 262714
rect 205265 262656 205270 262712
rect 205326 262656 296730 262712
rect 205265 262654 296730 262656
rect 366725 262714 366791 262717
rect 458398 262714 458404 262716
rect 366725 262712 458404 262714
rect 366725 262656 366730 262712
rect 366786 262656 458404 262712
rect 366725 262654 458404 262656
rect 205265 262651 205331 262654
rect 366725 262651 366791 262654
rect 458398 262652 458404 262654
rect 458468 262652 458474 262716
rect 85941 262578 86007 262581
rect 86534 262578 86540 262580
rect 85941 262576 86540 262578
rect 85941 262520 85946 262576
rect 86002 262520 86540 262576
rect 85941 262518 86540 262520
rect 85941 262515 86007 262518
rect 86534 262516 86540 262518
rect 86604 262516 86610 262580
rect 114645 262578 114711 262581
rect 423949 262580 424015 262581
rect 115790 262578 115796 262580
rect 114645 262576 115796 262578
rect 114645 262520 114650 262576
rect 114706 262520 115796 262576
rect 114645 262518 115796 262520
rect 114645 262515 114711 262518
rect 115790 262516 115796 262518
rect 115860 262516 115866 262580
rect 423949 262576 423996 262580
rect 424060 262578 424066 262580
rect 423949 262520 423954 262576
rect 423949 262516 423996 262520
rect 424060 262518 424106 262578
rect 424060 262516 424066 262518
rect 423949 262515 424015 262516
rect 106406 262380 106412 262444
rect 106476 262442 106482 262444
rect 107561 262442 107627 262445
rect 106476 262440 107627 262442
rect 106476 262384 107566 262440
rect 107622 262384 107627 262440
rect 106476 262382 107627 262384
rect 106476 262380 106482 262382
rect 107561 262379 107627 262382
rect 183134 262380 183140 262444
rect 183204 262442 183210 262444
rect 183461 262442 183527 262445
rect 183204 262440 183527 262442
rect 183204 262384 183466 262440
rect 183522 262384 183527 262440
rect 183204 262382 183527 262384
rect 183204 262380 183210 262382
rect 183461 262379 183527 262382
rect 251173 262442 251239 262445
rect 252318 262442 252324 262444
rect 251173 262440 252324 262442
rect 251173 262384 251178 262440
rect 251234 262384 252324 262440
rect 251173 262382 252324 262384
rect 251173 262379 251239 262382
rect 252318 262380 252324 262382
rect 252388 262380 252394 262444
rect 259545 262442 259611 262445
rect 260598 262442 260604 262444
rect 259545 262440 260604 262442
rect 259545 262384 259550 262440
rect 259606 262384 260604 262440
rect 259545 262382 260604 262384
rect 259545 262379 259611 262382
rect 260598 262380 260604 262382
rect 260668 262380 260674 262444
rect 266353 262442 266419 262445
rect 267590 262442 267596 262444
rect 266353 262440 267596 262442
rect 266353 262384 266358 262440
rect 266414 262384 267596 262440
rect 266353 262382 267596 262384
rect 266353 262379 266419 262382
rect 267590 262380 267596 262382
rect 267660 262380 267666 262444
rect 403065 262442 403131 262445
rect 404118 262442 404124 262444
rect 403065 262440 404124 262442
rect 403065 262384 403070 262440
rect 403126 262384 404124 262440
rect 403065 262382 404124 262384
rect 403065 262379 403131 262382
rect 404118 262380 404124 262382
rect 404188 262380 404194 262444
rect 411253 262442 411319 262445
rect 412398 262442 412404 262444
rect 411253 262440 412404 262442
rect 411253 262384 411258 262440
rect 411314 262384 412404 262440
rect 411253 262382 412404 262384
rect 411253 262379 411319 262382
rect 412398 262380 412404 262382
rect 412468 262380 412474 262444
rect 580901 262442 580967 262445
rect 583520 262442 584960 262532
rect 580901 262440 584960 262442
rect 580901 262384 580906 262440
rect 580962 262384 584960 262440
rect 580901 262382 584960 262384
rect 580901 262379 580967 262382
rect 77293 262306 77359 262309
rect 78254 262306 78260 262308
rect 77293 262304 78260 262306
rect 77293 262248 77298 262304
rect 77354 262248 78260 262304
rect 77293 262246 78260 262248
rect 77293 262243 77359 262246
rect 78254 262244 78260 262246
rect 78324 262244 78330 262308
rect 97022 262244 97028 262308
rect 97092 262306 97098 262308
rect 97901 262306 97967 262309
rect 97092 262304 97967 262306
rect 97092 262248 97906 262304
rect 97962 262248 97967 262304
rect 97092 262246 97967 262248
rect 97092 262244 97098 262246
rect 97901 262243 97967 262246
rect 98126 262244 98132 262308
rect 98196 262306 98202 262308
rect 99281 262306 99347 262309
rect 107561 262308 107627 262309
rect 107510 262306 107516 262308
rect 98196 262304 99347 262306
rect 98196 262248 99286 262304
rect 99342 262248 99347 262304
rect 98196 262246 99347 262248
rect 107470 262246 107516 262306
rect 107580 262304 107627 262308
rect 107622 262248 107627 262304
rect 98196 262244 98202 262246
rect 99281 262243 99347 262246
rect 107510 262244 107516 262246
rect 107580 262244 107627 262248
rect 107561 262243 107627 262244
rect 110413 262306 110479 262309
rect 111190 262306 111196 262308
rect 110413 262304 111196 262306
rect 110413 262248 110418 262304
rect 110474 262248 111196 262304
rect 110413 262246 111196 262248
rect 110413 262243 110479 262246
rect 111190 262244 111196 262246
rect 111260 262244 111266 262308
rect 113173 262306 113239 262309
rect 114318 262306 114324 262308
rect 113173 262304 114324 262306
rect 113173 262248 113178 262304
rect 113234 262248 114324 262304
rect 113173 262246 114324 262248
rect 113173 262243 113239 262246
rect 114318 262244 114324 262246
rect 114388 262244 114394 262308
rect 183369 262306 183435 262309
rect 183502 262306 183508 262308
rect 183369 262304 183508 262306
rect 183369 262248 183374 262304
rect 183430 262248 183508 262304
rect 183369 262246 183508 262248
rect 183369 262243 183435 262246
rect 183502 262244 183508 262246
rect 183572 262244 183578 262308
rect 237373 262306 237439 262309
rect 238150 262306 238156 262308
rect 237373 262304 238156 262306
rect 237373 262248 237378 262304
rect 237434 262248 238156 262304
rect 237373 262246 238156 262248
rect 237373 262243 237439 262246
rect 238150 262244 238156 262246
rect 238220 262244 238226 262308
rect 240133 262306 240199 262309
rect 240542 262306 240548 262308
rect 240133 262304 240548 262306
rect 240133 262248 240138 262304
rect 240194 262248 240548 262304
rect 240133 262246 240548 262248
rect 240133 262243 240199 262246
rect 240542 262244 240548 262246
rect 240612 262244 240618 262308
rect 241513 262306 241579 262309
rect 241646 262306 241652 262308
rect 241513 262304 241652 262306
rect 241513 262248 241518 262304
rect 241574 262248 241652 262304
rect 241513 262246 241652 262248
rect 241513 262243 241579 262246
rect 241646 262244 241652 262246
rect 241716 262244 241722 262308
rect 244273 262306 244339 262309
rect 245326 262306 245332 262308
rect 244273 262304 245332 262306
rect 244273 262248 244278 262304
rect 244334 262248 245332 262304
rect 244273 262246 245332 262248
rect 244273 262243 244339 262246
rect 245326 262244 245332 262246
rect 245396 262244 245402 262308
rect 245653 262306 245719 262309
rect 246430 262306 246436 262308
rect 245653 262304 246436 262306
rect 245653 262248 245658 262304
rect 245714 262248 246436 262304
rect 245653 262246 246436 262248
rect 245653 262243 245719 262246
rect 246430 262244 246436 262246
rect 246500 262244 246506 262308
rect 248413 262306 248479 262309
rect 248638 262306 248644 262308
rect 248413 262304 248644 262306
rect 248413 262248 248418 262304
rect 248474 262248 248644 262304
rect 248413 262246 248644 262248
rect 248413 262243 248479 262246
rect 248638 262244 248644 262246
rect 248708 262244 248714 262308
rect 249793 262306 249859 262309
rect 251265 262308 251331 262309
rect 250110 262306 250116 262308
rect 249793 262304 250116 262306
rect 249793 262248 249798 262304
rect 249854 262248 250116 262304
rect 249793 262246 250116 262248
rect 249793 262243 249859 262246
rect 250110 262244 250116 262246
rect 250180 262244 250186 262308
rect 251214 262306 251220 262308
rect 251174 262246 251220 262306
rect 251284 262304 251331 262308
rect 251326 262248 251331 262304
rect 251214 262244 251220 262246
rect 251284 262244 251331 262248
rect 251265 262243 251331 262244
rect 252645 262306 252711 262309
rect 253422 262306 253428 262308
rect 252645 262304 253428 262306
rect 252645 262248 252650 262304
rect 252706 262248 253428 262304
rect 252645 262246 253428 262248
rect 252645 262243 252711 262246
rect 253422 262244 253428 262246
rect 253492 262244 253498 262308
rect 253933 262306 253999 262309
rect 254526 262306 254532 262308
rect 253933 262304 254532 262306
rect 253933 262248 253938 262304
rect 253994 262248 254532 262304
rect 253933 262246 254532 262248
rect 253933 262243 253999 262246
rect 254526 262244 254532 262246
rect 254596 262244 254602 262308
rect 255313 262306 255379 262309
rect 255814 262306 255820 262308
rect 255313 262304 255820 262306
rect 255313 262248 255318 262304
rect 255374 262248 255820 262304
rect 255313 262246 255820 262248
rect 255313 262243 255379 262246
rect 255814 262244 255820 262246
rect 255884 262244 255890 262308
rect 256693 262306 256759 262309
rect 259453 262308 259519 262309
rect 256918 262306 256924 262308
rect 256693 262304 256924 262306
rect 256693 262248 256698 262304
rect 256754 262248 256924 262304
rect 256693 262246 256924 262248
rect 256693 262243 256759 262246
rect 256918 262244 256924 262246
rect 256988 262244 256994 262308
rect 259453 262304 259500 262308
rect 259564 262306 259570 262308
rect 263593 262306 263659 262309
rect 263910 262306 263916 262308
rect 259453 262248 259458 262304
rect 259453 262244 259500 262248
rect 259564 262246 259610 262306
rect 263593 262304 263916 262306
rect 263593 262248 263598 262304
rect 263654 262248 263916 262304
rect 263593 262246 263916 262248
rect 259564 262244 259570 262246
rect 259453 262243 259519 262244
rect 263593 262243 263659 262246
rect 263910 262244 263916 262246
rect 263980 262244 263986 262308
rect 266302 262244 266308 262308
rect 266372 262306 266378 262308
rect 266445 262306 266511 262309
rect 266372 262304 266511 262306
rect 266372 262248 266450 262304
rect 266506 262248 266511 262304
rect 266372 262246 266511 262248
rect 266372 262244 266378 262246
rect 266445 262243 266511 262246
rect 267733 262306 267799 262309
rect 268694 262306 268700 262308
rect 267733 262304 268700 262306
rect 267733 262248 267738 262304
rect 267794 262248 268700 262304
rect 267733 262246 268700 262248
rect 267733 262243 267799 262246
rect 268694 262244 268700 262246
rect 268764 262244 268770 262308
rect 276974 262244 276980 262308
rect 277044 262306 277050 262308
rect 277301 262306 277367 262309
rect 277044 262304 277367 262306
rect 277044 262248 277306 262304
rect 277362 262248 277367 262304
rect 277044 262246 277367 262248
rect 277044 262244 277050 262246
rect 277301 262243 277367 262246
rect 278078 262244 278084 262308
rect 278148 262306 278154 262308
rect 278681 262306 278747 262309
rect 278148 262304 278747 262306
rect 278148 262248 278686 262304
rect 278742 262248 278747 262304
rect 278148 262246 278747 262248
rect 278148 262244 278154 262246
rect 278681 262243 278747 262246
rect 303470 262244 303476 262308
rect 303540 262244 303546 262308
rect 396022 262244 396028 262308
rect 396092 262306 396098 262308
rect 396165 262306 396231 262309
rect 396092 262304 396231 262306
rect 396092 262248 396170 262304
rect 396226 262248 396231 262304
rect 396092 262246 396231 262248
rect 396092 262244 396098 262246
rect 199326 262108 199332 262172
rect 199396 262170 199402 262172
rect 303478 262170 303538 262244
rect 396165 262243 396231 262246
rect 398833 262306 398899 262309
rect 399518 262306 399524 262308
rect 398833 262304 399524 262306
rect 398833 262248 398838 262304
rect 398894 262248 399524 262304
rect 398833 262246 399524 262248
rect 398833 262243 398899 262246
rect 399518 262244 399524 262246
rect 399588 262244 399594 262308
rect 400213 262306 400279 262309
rect 402973 262308 403039 262309
rect 400438 262306 400444 262308
rect 400213 262304 400444 262306
rect 400213 262248 400218 262304
rect 400274 262248 400444 262304
rect 400213 262246 400444 262248
rect 400213 262243 400279 262246
rect 400438 262244 400444 262246
rect 400508 262244 400514 262308
rect 402973 262304 403020 262308
rect 403084 262306 403090 262308
rect 405733 262306 405799 262309
rect 406510 262306 406516 262308
rect 402973 262248 402978 262304
rect 402973 262244 403020 262248
rect 403084 262246 403130 262306
rect 405733 262304 406516 262306
rect 405733 262248 405738 262304
rect 405794 262248 406516 262304
rect 405733 262246 406516 262248
rect 403084 262244 403090 262246
rect 402973 262243 403039 262244
rect 405733 262243 405799 262246
rect 406510 262244 406516 262246
rect 406580 262244 406586 262308
rect 407205 262306 407271 262309
rect 407614 262306 407620 262308
rect 407205 262304 407620 262306
rect 407205 262248 407210 262304
rect 407266 262248 407620 262304
rect 407205 262246 407620 262248
rect 407205 262243 407271 262246
rect 407614 262244 407620 262246
rect 407684 262244 407690 262308
rect 408493 262306 408559 262309
rect 408718 262306 408724 262308
rect 408493 262304 408724 262306
rect 408493 262248 408498 262304
rect 408554 262248 408724 262304
rect 408493 262246 408724 262248
rect 408493 262243 408559 262246
rect 408718 262244 408724 262246
rect 408788 262244 408794 262308
rect 409873 262306 409939 262309
rect 411345 262308 411411 262309
rect 410006 262306 410012 262308
rect 409873 262304 410012 262306
rect 409873 262248 409878 262304
rect 409934 262248 410012 262304
rect 409873 262246 410012 262248
rect 409873 262243 409939 262246
rect 410006 262244 410012 262246
rect 410076 262244 410082 262308
rect 411294 262306 411300 262308
rect 411254 262246 411300 262306
rect 411364 262304 411411 262308
rect 411406 262248 411411 262304
rect 411294 262244 411300 262246
rect 411364 262244 411411 262248
rect 411345 262243 411411 262244
rect 414013 262306 414079 262309
rect 414606 262306 414612 262308
rect 414013 262304 414612 262306
rect 414013 262248 414018 262304
rect 414074 262248 414612 262304
rect 414013 262246 414612 262248
rect 414013 262243 414079 262246
rect 414606 262244 414612 262246
rect 414676 262244 414682 262308
rect 416773 262306 416839 262309
rect 416998 262306 417004 262308
rect 416773 262304 417004 262306
rect 416773 262248 416778 262304
rect 416834 262248 417004 262304
rect 416773 262246 417004 262248
rect 416773 262243 416839 262246
rect 416998 262244 417004 262246
rect 417068 262244 417074 262308
rect 422886 262244 422892 262308
rect 422956 262306 422962 262308
rect 423581 262306 423647 262309
rect 422956 262304 423647 262306
rect 422956 262248 423586 262304
rect 423642 262248 423647 262304
rect 422956 262246 423647 262248
rect 422956 262244 422962 262246
rect 423581 262243 423647 262246
rect 428273 262306 428339 262309
rect 428590 262306 428596 262308
rect 428273 262304 428596 262306
rect 428273 262248 428278 262304
rect 428334 262248 428596 262304
rect 428273 262246 428596 262248
rect 428273 262243 428339 262246
rect 428590 262244 428596 262246
rect 428660 262244 428666 262308
rect 430665 262306 430731 262309
rect 431166 262306 431172 262308
rect 430665 262304 431172 262306
rect 430665 262248 430670 262304
rect 430726 262248 431172 262304
rect 430665 262246 431172 262248
rect 430665 262243 430731 262246
rect 431166 262244 431172 262246
rect 431236 262244 431242 262308
rect 436093 262306 436159 262309
rect 436870 262306 436876 262308
rect 436093 262304 436876 262306
rect 436093 262248 436098 262304
rect 436154 262248 436876 262304
rect 436093 262246 436876 262248
rect 436093 262243 436159 262246
rect 436870 262244 436876 262246
rect 436940 262244 436946 262308
rect 439262 262244 439268 262308
rect 439332 262306 439338 262308
rect 440141 262306 440207 262309
rect 439332 262304 440207 262306
rect 439332 262248 440146 262304
rect 440202 262248 440207 262304
rect 439332 262246 440207 262248
rect 439332 262244 439338 262246
rect 440141 262243 440207 262246
rect 503110 262244 503116 262308
rect 503180 262306 503186 262308
rect 503621 262306 503687 262309
rect 503180 262304 503687 262306
rect 503180 262248 503626 262304
rect 503682 262248 503687 262304
rect 583520 262292 584960 262382
rect 503180 262246 503687 262248
rect 503180 262244 503186 262246
rect 503621 262243 503687 262246
rect 199396 262110 303538 262170
rect 199396 262108 199402 262110
rect 377990 260884 377996 260948
rect 378060 260946 378066 260948
rect 380341 260946 380407 260949
rect 378060 260944 380407 260946
rect 378060 260888 380346 260944
rect 380402 260888 380407 260944
rect 378060 260886 380407 260888
rect 378060 260884 378066 260886
rect 47710 260748 47716 260812
rect 47780 260810 47786 260812
rect 50429 260810 50495 260813
rect 47780 260808 50495 260810
rect 47780 260752 50434 260808
rect 50490 260752 50495 260808
rect 47780 260750 50495 260752
rect 47780 260748 47786 260750
rect 50429 260747 50495 260750
rect 379470 260677 379530 260886
rect 380341 260883 380407 260886
rect 379470 260672 379579 260677
rect 379470 260616 379518 260672
rect 379574 260616 379579 260672
rect 379470 260614 379579 260616
rect 379513 260611 379579 260614
rect 44950 260340 44956 260404
rect 45020 260402 45026 260404
rect 46473 260402 46539 260405
rect 80145 260402 80211 260405
rect 45020 260400 80211 260402
rect 45020 260344 46478 260400
rect 46534 260344 80150 260400
rect 80206 260344 80211 260400
rect 45020 260342 80211 260344
rect 45020 260340 45026 260342
rect 46473 260339 46539 260342
rect 80145 260339 80211 260342
rect 50429 260266 50495 260269
rect 96521 260266 96587 260269
rect 50429 260264 96587 260266
rect 50429 260208 50434 260264
rect 50490 260208 96526 260264
rect 96582 260208 96587 260264
rect 50429 260206 96587 260208
rect 50429 260203 50495 260206
rect 96521 260203 96587 260206
rect 44766 260068 44772 260132
rect 44836 260130 44842 260132
rect 46381 260130 46447 260133
rect 114645 260130 114711 260133
rect 44836 260128 114711 260130
rect 44836 260072 46386 260128
rect 46442 260072 114650 260128
rect 114706 260072 114711 260128
rect 44836 260070 114711 260072
rect 44836 260068 44842 260070
rect 46381 260067 46447 260070
rect 114645 260067 114711 260070
rect 377806 260068 377812 260132
rect 377876 260130 377882 260132
rect 393957 260130 394023 260133
rect 377876 260128 394023 260130
rect 377876 260072 393962 260128
rect 394018 260072 394023 260128
rect 377876 260070 394023 260072
rect 377876 260068 377882 260070
rect 393957 260067 394023 260070
rect -960 257682 480 257772
rect 2773 257682 2839 257685
rect -960 257680 2839 257682
rect -960 257624 2778 257680
rect 2834 257624 2839 257680
rect -960 257622 2839 257624
rect -960 257532 480 257622
rect 2773 257619 2839 257622
rect 583520 249508 584960 249748
rect -960 245020 480 245260
rect 510838 241436 510844 241500
rect 510908 241498 510914 241500
rect 511901 241498 511967 241501
rect 510908 241496 511967 241498
rect 510908 241440 511906 241496
rect 511962 241440 511967 241496
rect 510908 241438 511967 241440
rect 510908 241436 510914 241438
rect 511901 241435 511967 241438
rect 393957 240818 394023 240821
rect 416773 240818 416839 240821
rect 393957 240816 416839 240818
rect 393957 240760 393962 240816
rect 394018 240760 416778 240816
rect 416834 240760 416839 240816
rect 393957 240758 416839 240760
rect 393957 240755 394023 240758
rect 416773 240755 416839 240758
rect 178534 240212 178540 240276
rect 178604 240274 178610 240276
rect 179321 240274 179387 240277
rect 178604 240272 179387 240274
rect 178604 240216 179326 240272
rect 179382 240216 179387 240272
rect 178604 240214 179387 240216
rect 178604 240212 178610 240214
rect 179321 240211 179387 240214
rect 179638 240212 179644 240276
rect 179708 240274 179714 240276
rect 180149 240274 180215 240277
rect 190913 240276 190979 240277
rect 190862 240274 190868 240276
rect 179708 240272 180215 240274
rect 179708 240216 180154 240272
rect 180210 240216 180215 240272
rect 179708 240214 180215 240216
rect 190822 240214 190868 240274
rect 190932 240272 190979 240276
rect 190974 240216 190979 240272
rect 179708 240212 179714 240214
rect 180149 240211 180215 240214
rect 190862 240212 190868 240214
rect 190932 240212 190979 240216
rect 217542 240212 217548 240276
rect 217612 240274 217618 240276
rect 220077 240274 220143 240277
rect 217612 240272 220143 240274
rect 217612 240216 220082 240272
rect 220138 240216 220143 240272
rect 217612 240214 220143 240216
rect 217612 240212 217618 240214
rect 190913 240211 190979 240212
rect 220077 240211 220143 240214
rect 338430 240212 338436 240276
rect 338500 240274 338506 240276
rect 339401 240274 339467 240277
rect 338500 240272 339467 240274
rect 338500 240216 339406 240272
rect 339462 240216 339467 240272
rect 338500 240214 339467 240216
rect 338500 240212 338506 240214
rect 339401 240211 339467 240214
rect 339718 240212 339724 240276
rect 339788 240274 339794 240276
rect 340045 240274 340111 240277
rect 339788 240272 340111 240274
rect 339788 240216 340050 240272
rect 340106 240216 340111 240272
rect 339788 240214 340111 240216
rect 339788 240212 339794 240214
rect 340045 240211 340111 240214
rect 350942 240212 350948 240276
rect 351012 240274 351018 240276
rect 351545 240274 351611 240277
rect 351012 240272 351611 240274
rect 351012 240216 351550 240272
rect 351606 240216 351611 240272
rect 351012 240214 351611 240216
rect 351012 240212 351018 240214
rect 351545 240211 351611 240214
rect 379646 240212 379652 240276
rect 379716 240274 379722 240276
rect 379881 240274 379947 240277
rect 379716 240272 379947 240274
rect 379716 240216 379886 240272
rect 379942 240216 379947 240272
rect 379716 240214 379947 240216
rect 379716 240212 379722 240214
rect 379881 240211 379947 240214
rect 498510 240212 498516 240276
rect 498580 240274 498586 240276
rect 499021 240274 499087 240277
rect 498580 240272 499087 240274
rect 498580 240216 499026 240272
rect 499082 240216 499087 240272
rect 498580 240214 499087 240216
rect 498580 240212 498586 240214
rect 499021 240211 499087 240214
rect 499798 240212 499804 240276
rect 499868 240274 499874 240276
rect 500769 240274 500835 240277
rect 499868 240272 500835 240274
rect 499868 240216 500774 240272
rect 500830 240216 500835 240272
rect 499868 240214 500835 240216
rect 499868 240212 499874 240214
rect 500769 240211 500835 240214
rect 375833 239866 375899 239869
rect 377254 239866 377260 239868
rect 375833 239864 377260 239866
rect 375833 239808 375838 239864
rect 375894 239808 377260 239864
rect 375833 239806 377260 239808
rect 375833 239803 375899 239806
rect 377254 239804 377260 239806
rect 377324 239866 377330 239868
rect 378041 239866 378107 239869
rect 377324 239864 378107 239866
rect 377324 239808 378046 239864
rect 378102 239808 378107 239864
rect 377324 239806 378107 239808
rect 377324 239804 377330 239806
rect 378041 239803 378107 239806
rect 379697 239596 379763 239597
rect 379646 239594 379652 239596
rect 379606 239534 379652 239594
rect 379716 239592 379763 239596
rect 379758 239536 379763 239592
rect 379646 239532 379652 239534
rect 379716 239532 379763 239536
rect 379697 239531 379763 239532
rect 377990 239396 377996 239460
rect 378060 239458 378066 239460
rect 393957 239458 394023 239461
rect 378060 239456 394023 239458
rect 378060 239400 393962 239456
rect 394018 239400 394023 239456
rect 378060 239398 394023 239400
rect 378060 239396 378066 239398
rect 393957 239395 394023 239398
rect 47894 238580 47900 238644
rect 47964 238642 47970 238644
rect 58893 238642 58959 238645
rect 47964 238640 58959 238642
rect 47964 238584 58898 238640
rect 58954 238584 58959 238640
rect 47964 238582 58959 238584
rect 47964 238580 47970 238582
rect 58893 238579 58959 238582
rect 57145 237420 57211 237421
rect 57094 237356 57100 237420
rect 57164 237418 57211 237420
rect 58617 237418 58683 237421
rect 58893 237418 58959 237421
rect 57164 237416 57256 237418
rect 57206 237360 57256 237416
rect 57164 237358 57256 237360
rect 58617 237416 58959 237418
rect 58617 237360 58622 237416
rect 58678 237360 58898 237416
rect 58954 237360 58959 237416
rect 58617 237358 58959 237360
rect 57164 237356 57211 237358
rect 57145 237355 57211 237356
rect 58617 237355 58683 237358
rect 58893 237355 58959 237358
rect 583520 236588 584960 236828
rect 518985 234562 519051 234565
rect 519353 234562 519419 234565
rect 516558 234560 519419 234562
rect 516558 234504 518990 234560
rect 519046 234504 519358 234560
rect 519414 234504 519419 234560
rect 516558 234502 519419 234504
rect 516558 234190 516618 234502
rect 518985 234499 519051 234502
rect 519353 234499 519419 234502
rect 196558 234018 196618 234190
rect 198825 234018 198891 234021
rect 199193 234018 199259 234021
rect 196558 234016 199259 234018
rect 196558 233960 198830 234016
rect 198886 233960 199198 234016
rect 199254 233960 199259 234016
rect 196558 233958 199259 233960
rect 356562 234018 356622 234190
rect 358905 234018 358971 234021
rect 359273 234018 359339 234021
rect 356562 234016 359339 234018
rect 356562 233960 358910 234016
rect 358966 233960 359278 234016
rect 359334 233960 359339 234016
rect 356562 233958 359339 233960
rect 198825 233955 198891 233958
rect 199193 233955 199259 233958
rect 358905 233955 358971 233958
rect 359273 233955 359339 233958
rect -960 232372 480 232612
rect 580901 223954 580967 223957
rect 583520 223954 584960 224044
rect 580901 223952 584960 223954
rect 580901 223896 580906 223952
rect 580962 223896 584960 223952
rect 580901 223894 584960 223896
rect 580901 223891 580967 223894
rect 583520 223804 584960 223894
rect -960 220010 480 220100
rect -960 219950 674 220010
rect -960 219874 480 219950
rect 614 219874 674 219950
rect -960 219860 674 219874
rect 246 219814 674 219860
rect 246 219466 306 219814
rect 51574 219466 51580 219468
rect 246 219406 51580 219466
rect 51574 219404 51580 219406
rect 51644 219404 51650 219468
rect 583520 211020 584960 211260
rect -960 207362 480 207452
rect 2773 207362 2839 207365
rect -960 207360 2839 207362
rect -960 207304 2778 207360
rect 2834 207304 2839 207360
rect -960 207302 2839 207304
rect -960 207212 480 207302
rect 2773 207299 2839 207302
rect 583520 198236 584960 198476
rect -960 194700 480 194940
rect 56777 193218 56843 193221
rect 57605 193218 57671 193221
rect 56777 193216 57671 193218
rect 56777 193160 56782 193216
rect 56838 193160 57610 193216
rect 57666 193160 57671 193216
rect 56777 193158 57671 193160
rect 56777 193155 56843 193158
rect 57605 193155 57671 193158
rect 216765 193218 216831 193221
rect 217133 193218 217199 193221
rect 216765 193216 217199 193218
rect 216765 193160 216770 193216
rect 216826 193160 217138 193216
rect 217194 193160 217199 193216
rect 216765 193158 217199 193160
rect 216765 193155 216831 193158
rect 217133 193155 217199 193158
rect 377213 193218 377279 193221
rect 377949 193218 378015 193221
rect 377213 193216 378015 193218
rect 377213 193160 377218 193216
rect 377274 193160 377954 193216
rect 378010 193160 378015 193216
rect 377213 193158 378015 193160
rect 377213 193155 377279 193158
rect 377949 193155 378015 193158
rect 57605 191858 57671 191861
rect 60002 191858 60062 191894
rect 219390 191864 220064 191924
rect 379838 191864 380052 191924
rect 57605 191856 60062 191858
rect 57605 191800 57610 191856
rect 57666 191800 60062 191856
rect 57605 191798 60062 191800
rect 216765 191858 216831 191861
rect 219390 191858 219450 191864
rect 216765 191856 219450 191858
rect 216765 191800 216770 191856
rect 216826 191800 219450 191856
rect 216765 191798 219450 191800
rect 377949 191858 378015 191861
rect 379838 191858 379898 191864
rect 377949 191856 379898 191858
rect 377949 191800 377954 191856
rect 378010 191800 379898 191856
rect 377949 191798 379898 191800
rect 57605 191795 57671 191798
rect 216765 191795 216831 191798
rect 377949 191795 378015 191798
rect 56593 191722 56659 191725
rect 56777 191722 56843 191725
rect 56593 191720 56843 191722
rect 56593 191664 56598 191720
rect 56654 191664 56782 191720
rect 56838 191664 56843 191720
rect 56593 191662 56843 191664
rect 56593 191659 56659 191662
rect 56777 191659 56843 191662
rect 216857 191722 216923 191725
rect 217685 191722 217751 191725
rect 216857 191720 217751 191722
rect 216857 191664 216862 191720
rect 216918 191664 217690 191720
rect 217746 191664 217751 191720
rect 216857 191662 217751 191664
rect 216857 191659 216923 191662
rect 217685 191659 217751 191662
rect 376845 191722 376911 191725
rect 377857 191722 377923 191725
rect 376845 191720 377923 191722
rect 376845 191664 376850 191720
rect 376906 191664 377862 191720
rect 377918 191664 377923 191720
rect 376845 191662 377923 191664
rect 376845 191659 376911 191662
rect 377857 191659 377923 191662
rect 217685 191042 217751 191045
rect 217685 191040 219450 191042
rect 217685 190984 217690 191040
rect 217746 190984 219450 191040
rect 217685 190982 219450 190984
rect 217685 190979 217751 190982
rect 219390 190972 219450 190982
rect 56777 190906 56843 190909
rect 60002 190906 60062 190942
rect 219390 190912 220064 190972
rect 379838 190912 380052 190972
rect 56777 190904 60062 190906
rect 56777 190848 56782 190904
rect 56838 190848 60062 190904
rect 56777 190846 60062 190848
rect 377857 190906 377923 190909
rect 379838 190906 379898 190912
rect 377857 190904 379898 190906
rect 377857 190848 377862 190904
rect 377918 190848 379898 190904
rect 377857 190846 379898 190848
rect 56777 190843 56843 190846
rect 377857 190843 377923 190846
rect 57697 188730 57763 188733
rect 60002 188730 60062 188766
rect 219390 188736 220064 188796
rect 379838 188736 380052 188796
rect 57697 188728 60062 188730
rect 57697 188672 57702 188728
rect 57758 188672 60062 188728
rect 57697 188670 60062 188672
rect 217777 188730 217843 188733
rect 219390 188730 219450 188736
rect 217777 188728 219450 188730
rect 217777 188672 217782 188728
rect 217838 188672 219450 188728
rect 217777 188670 219450 188672
rect 376937 188730 377003 188733
rect 379838 188730 379898 188736
rect 376937 188728 379898 188730
rect 376937 188672 376942 188728
rect 376998 188672 379898 188728
rect 376937 188670 379898 188672
rect 57697 188667 57763 188670
rect 217777 188667 217843 188670
rect 376937 188667 377003 188670
rect 56869 187914 56935 187917
rect 57421 187914 57487 187917
rect 376937 187914 377003 187917
rect 377213 187914 377279 187917
rect 56869 187912 59554 187914
rect 56869 187856 56874 187912
rect 56930 187856 57426 187912
rect 57482 187856 59554 187912
rect 56869 187854 59554 187856
rect 56869 187851 56935 187854
rect 57421 187851 57487 187854
rect 59494 187844 59554 187854
rect 376937 187912 377279 187914
rect 376937 187856 376942 187912
rect 376998 187856 377218 187912
rect 377274 187856 377279 187912
rect 376937 187854 377279 187856
rect 376937 187851 377003 187854
rect 377213 187851 377279 187854
rect 59494 187784 60032 187844
rect 219390 187784 220064 187844
rect 379838 187784 380052 187844
rect 57329 187778 57395 187781
rect 57697 187778 57763 187781
rect 57329 187776 57763 187778
rect 57329 187720 57334 187776
rect 57390 187720 57702 187776
rect 57758 187720 57763 187776
rect 57329 187718 57763 187720
rect 57329 187715 57395 187718
rect 57697 187715 57763 187718
rect 216673 187778 216739 187781
rect 217961 187778 218027 187781
rect 219390 187778 219450 187784
rect 216673 187776 219450 187778
rect 216673 187720 216678 187776
rect 216734 187720 217966 187776
rect 218022 187720 219450 187776
rect 216673 187718 219450 187720
rect 377305 187778 377371 187781
rect 378041 187778 378107 187781
rect 379838 187778 379898 187784
rect 377305 187776 379898 187778
rect 377305 187720 377310 187776
rect 377366 187720 378046 187776
rect 378102 187720 379898 187776
rect 377305 187718 379898 187720
rect 216673 187715 216739 187718
rect 217961 187715 218027 187718
rect 377305 187715 377371 187718
rect 378041 187715 378107 187718
rect 57145 185738 57211 185741
rect 57513 185738 57579 185741
rect 60002 185738 60062 186046
rect 219390 186016 220064 186076
rect 379838 186016 380052 186076
rect 217501 186010 217567 186013
rect 219390 186010 219450 186016
rect 217501 186008 219450 186010
rect 217501 185952 217506 186008
rect 217562 185952 219450 186008
rect 217501 185950 219450 185952
rect 376937 186010 377003 186013
rect 379838 186010 379898 186016
rect 376937 186008 379898 186010
rect 376937 185952 376942 186008
rect 376998 185952 379898 186008
rect 376937 185950 379898 185952
rect 217501 185947 217567 185950
rect 376937 185947 377003 185950
rect 57145 185736 60062 185738
rect 57145 185680 57150 185736
rect 57206 185680 57518 185736
rect 57574 185680 60062 185736
rect 57145 185678 60062 185680
rect 57145 185675 57211 185678
rect 57513 185675 57579 185678
rect 580901 185602 580967 185605
rect 583520 185602 584960 185692
rect 580901 185600 584960 185602
rect 580901 185544 580906 185600
rect 580962 185544 584960 185600
rect 580901 185542 584960 185544
rect 580901 185539 580967 185542
rect 56685 185466 56751 185469
rect 57697 185466 57763 185469
rect 56685 185464 60062 185466
rect 56685 185408 56690 185464
rect 56746 185408 57702 185464
rect 57758 185408 60062 185464
rect 583520 185452 584960 185542
rect 56685 185406 60062 185408
rect 56685 185403 56751 185406
rect 57697 185403 57763 185406
rect 60002 184958 60062 185406
rect 216949 185058 217015 185061
rect 217409 185058 217475 185061
rect 377121 185058 377187 185061
rect 216949 185056 219450 185058
rect 216949 185000 216954 185056
rect 217010 185000 217414 185056
rect 217470 185000 219450 185056
rect 216949 184998 219450 185000
rect 216949 184995 217015 184998
rect 217409 184995 217475 184998
rect 219390 184988 219450 184998
rect 377121 185056 379898 185058
rect 377121 185000 377126 185056
rect 377182 185000 379898 185056
rect 377121 184998 379898 185000
rect 377121 184995 377187 184998
rect 379838 184988 379898 184998
rect 219390 184928 220064 184988
rect 379838 184928 380052 184988
rect 57053 183562 57119 183565
rect 57421 183562 57487 183565
rect 377489 183562 377555 183565
rect 377765 183562 377831 183565
rect 57053 183560 60062 183562
rect 57053 183504 57058 183560
rect 57114 183504 57426 183560
rect 57482 183504 60062 183560
rect 57053 183502 60062 183504
rect 57053 183499 57119 183502
rect 57421 183499 57487 183502
rect 60002 183190 60062 183502
rect 377489 183560 379530 183562
rect 377489 183504 377494 183560
rect 377550 183504 377770 183560
rect 377826 183504 379530 183560
rect 377489 183502 379530 183504
rect 377489 183499 377555 183502
rect 377765 183499 377831 183502
rect 217409 183290 217475 183293
rect 217869 183290 217935 183293
rect 217409 183288 219450 183290
rect 217409 183232 217414 183288
rect 217470 183232 217874 183288
rect 217930 183232 219450 183288
rect 217409 183230 219450 183232
rect 217409 183227 217475 183230
rect 217869 183227 217935 183230
rect 219390 183220 219450 183230
rect 379470 183220 379530 183502
rect 219390 183160 220064 183220
rect 379470 183160 380052 183220
rect -960 182188 480 182428
rect 198733 174994 198799 174997
rect 199377 174994 199443 174997
rect 358813 174994 358879 174997
rect 359549 174994 359615 174997
rect 196558 174992 199443 174994
rect 196558 174936 198738 174992
rect 198794 174936 199382 174992
rect 199438 174936 199443 174992
rect 196558 174934 199443 174936
rect 196558 174350 196618 174934
rect 198733 174931 198799 174934
rect 199377 174931 199443 174934
rect 356562 174992 359615 174994
rect 356562 174936 358818 174992
rect 358874 174936 359554 174992
rect 359610 174936 359615 174992
rect 356562 174934 359615 174936
rect 356562 174350 356622 174934
rect 358813 174931 358879 174934
rect 359549 174931 359615 174934
rect 516558 174314 516618 174350
rect 518893 174314 518959 174317
rect 516558 174312 518959 174314
rect 516558 174256 518898 174312
rect 518954 174256 518959 174312
rect 516558 174254 518959 174256
rect 518893 174251 518959 174254
rect 196558 172682 196618 172718
rect 199285 172682 199351 172685
rect 196558 172680 199351 172682
rect 196558 172624 199290 172680
rect 199346 172624 199351 172680
rect 196558 172622 199351 172624
rect 356562 172682 356622 172718
rect 359181 172682 359247 172685
rect 356562 172680 359247 172682
rect 356562 172624 359186 172680
rect 359242 172624 359247 172680
rect 356562 172622 359247 172624
rect 516558 172682 516618 172718
rect 519445 172682 519511 172685
rect 516558 172680 519511 172682
rect 516558 172624 519450 172680
rect 519506 172624 519511 172680
rect 583520 172668 584960 172908
rect 516558 172622 519511 172624
rect 199285 172619 199351 172622
rect 359181 172619 359247 172622
rect 519445 172619 519511 172622
rect 358813 172410 358879 172413
rect 359641 172410 359707 172413
rect 358813 172408 359707 172410
rect 358813 172352 358818 172408
rect 358874 172352 359646 172408
rect 359702 172352 359707 172408
rect 358813 172350 359707 172352
rect 358813 172347 358879 172350
rect 359641 172347 359707 172350
rect 196558 171322 196618 171358
rect 199101 171322 199167 171325
rect 196558 171320 199167 171322
rect 196558 171264 199106 171320
rect 199162 171264 199167 171320
rect 196558 171262 199167 171264
rect 356562 171322 356622 171358
rect 358813 171322 358879 171325
rect 356562 171320 358879 171322
rect 356562 171264 358818 171320
rect 358874 171264 358879 171320
rect 356562 171262 358879 171264
rect 516558 171322 516618 171358
rect 519077 171322 519143 171325
rect 516558 171320 519143 171322
rect 516558 171264 519082 171320
rect 519138 171264 519143 171320
rect 516558 171262 519143 171264
rect 199101 171259 199167 171262
rect 358813 171259 358879 171262
rect 519077 171259 519143 171262
rect 196558 169826 196618 169862
rect 198825 169826 198891 169829
rect 196558 169824 198891 169826
rect -960 169690 480 169780
rect 196558 169768 198830 169824
rect 198886 169768 198891 169824
rect 196558 169766 198891 169768
rect 356562 169826 356622 169862
rect 358905 169826 358971 169829
rect 359365 169826 359431 169829
rect 356562 169824 359431 169826
rect 356562 169768 358910 169824
rect 358966 169768 359370 169824
rect 359426 169768 359431 169824
rect 356562 169766 359431 169768
rect 516558 169826 516618 169862
rect 519077 169826 519143 169829
rect 516558 169824 519143 169826
rect 516558 169768 519082 169824
rect 519138 169768 519143 169824
rect 516558 169766 519143 169768
rect 198825 169763 198891 169766
rect 358905 169763 358971 169766
rect 359365 169763 359431 169766
rect 519077 169763 519143 169766
rect 2865 169690 2931 169693
rect -960 169688 2931 169690
rect -960 169632 2870 169688
rect 2926 169632 2931 169688
rect -960 169630 2931 169632
rect -960 169540 480 169630
rect 2865 169627 2931 169630
rect 519261 169010 519327 169013
rect 516558 169008 519327 169010
rect 516558 168952 519266 169008
rect 519322 168952 519327 169008
rect 516558 168950 519327 168952
rect 516558 168638 516618 168950
rect 519261 168947 519327 168950
rect 196558 168466 196618 168638
rect 356562 168602 356622 168638
rect 358997 168602 359063 168605
rect 356562 168600 359063 168602
rect 356562 168544 359002 168600
rect 359058 168544 359063 168600
rect 356562 168542 359063 168544
rect 358997 168539 359063 168542
rect 198733 168466 198799 168469
rect 199009 168466 199075 168469
rect 196558 168464 199075 168466
rect 196558 168408 198738 168464
rect 198794 168408 199014 168464
rect 199070 168408 199075 168464
rect 196558 168406 199075 168408
rect 198733 168403 198799 168406
rect 199009 168403 199075 168406
rect 59077 165610 59143 165613
rect 59077 165608 60062 165610
rect 59077 165552 59082 165608
rect 59138 165552 60062 165608
rect 59077 165550 60062 165552
rect 59077 165547 59143 165550
rect 60002 164966 60062 165550
rect 216673 165066 216739 165069
rect 376937 165066 377003 165069
rect 216673 165064 219450 165066
rect 216673 165008 216678 165064
rect 216734 165008 219450 165064
rect 216673 165006 219450 165008
rect 216673 165003 216739 165006
rect 219390 164996 219450 165006
rect 376937 165064 379530 165066
rect 376937 165008 376942 165064
rect 376998 165008 379530 165064
rect 376937 165006 379530 165008
rect 376937 165003 377003 165006
rect 379470 164996 379530 165006
rect 219390 164936 220064 164996
rect 379470 164936 380052 164996
rect 216673 163434 216739 163437
rect 376937 163434 377003 163437
rect 216673 163432 219450 163434
rect 216673 163376 216678 163432
rect 216734 163376 219450 163432
rect 216673 163374 219450 163376
rect 216673 163371 216739 163374
rect 219390 163364 219450 163374
rect 376937 163432 379530 163434
rect 376937 163376 376942 163432
rect 376998 163376 379530 163432
rect 376937 163374 379530 163376
rect 376937 163371 377003 163374
rect 379470 163364 379530 163374
rect 59862 163304 60032 163364
rect 219390 163304 220064 163364
rect 379470 163304 380052 163364
rect 57881 163298 57947 163301
rect 59862 163298 59922 163304
rect 57881 163296 59922 163298
rect 57881 163240 57886 163296
rect 57942 163240 59922 163296
rect 57881 163238 59922 163240
rect 57881 163235 57947 163238
rect 217041 163162 217107 163165
rect 376753 163162 376819 163165
rect 217041 163160 219450 163162
rect 217041 163104 217046 163160
rect 217102 163104 219450 163160
rect 217041 163102 219450 163104
rect 217041 163099 217107 163102
rect 219390 163092 219450 163102
rect 376753 163160 379530 163162
rect 376753 163104 376758 163160
rect 376814 163104 379530 163160
rect 376753 163102 379530 163104
rect 376753 163099 376819 163102
rect 379470 163092 379530 163102
rect 57462 162964 57468 163028
rect 57532 163026 57538 163028
rect 60002 163026 60062 163062
rect 219390 163032 220064 163092
rect 379470 163032 380052 163092
rect 57532 162966 60062 163026
rect 57532 162964 57538 162966
rect 583520 159884 584960 160124
rect -960 157178 480 157268
rect 2773 157178 2839 157181
rect -960 157176 2839 157178
rect -960 157120 2778 157176
rect 2834 157120 2839 157176
rect -960 157118 2839 157120
rect -960 157028 480 157118
rect 2773 157115 2839 157118
rect 96061 154732 96127 154733
rect 113357 154732 113423 154733
rect 96040 154668 96046 154732
rect 96110 154730 96127 154732
rect 113312 154730 113318 154732
rect 96110 154728 96202 154730
rect 96122 154672 96202 154728
rect 96110 154670 96202 154672
rect 113266 154670 113318 154730
rect 113382 154728 113423 154732
rect 163313 154732 163379 154733
rect 165889 154732 165955 154733
rect 163313 154730 163366 154732
rect 113418 154672 113423 154728
rect 96110 154668 96127 154670
rect 113312 154668 113318 154670
rect 113382 154668 113423 154672
rect 163274 154728 163366 154730
rect 163274 154672 163318 154728
rect 163274 154670 163366 154672
rect 96061 154667 96127 154668
rect 113357 154667 113423 154668
rect 163313 154668 163366 154670
rect 163430 154668 163436 154732
rect 165889 154730 165950 154732
rect 165858 154728 165950 154730
rect 165858 154672 165894 154728
rect 165858 154670 165950 154672
rect 165889 154668 165950 154670
rect 166014 154668 166020 154732
rect 163313 154667 163379 154668
rect 165889 154667 165955 154668
rect 261017 154596 261083 154597
rect 273529 154596 273595 154597
rect 261017 154594 261078 154596
rect 260986 154592 261078 154594
rect 260986 154536 261022 154592
rect 260986 154534 261078 154536
rect 261017 154532 261078 154534
rect 261142 154532 261148 154596
rect 273529 154594 273590 154596
rect 273498 154592 273590 154594
rect 273498 154536 273534 154592
rect 273498 154534 273590 154536
rect 273529 154532 273590 154534
rect 273654 154532 273660 154596
rect 261017 154531 261083 154532
rect 273529 154531 273595 154532
rect 418429 154460 418495 154461
rect 421005 154460 421071 154461
rect 425973 154460 426039 154461
rect 443453 154460 443519 154461
rect 57646 154396 57652 154460
rect 57716 154458 57722 154460
rect 148542 154458 148548 154460
rect 57716 154398 148548 154458
rect 57716 154396 57722 154398
rect 148542 154396 148548 154398
rect 148612 154396 148618 154460
rect 202454 154396 202460 154460
rect 202524 154458 202530 154460
rect 315798 154458 315804 154460
rect 202524 154398 315804 154458
rect 202524 154396 202530 154398
rect 315798 154396 315804 154398
rect 315868 154396 315874 154460
rect 418429 154458 418476 154460
rect 418384 154456 418476 154458
rect 418384 154400 418434 154456
rect 418384 154398 418476 154400
rect 418429 154396 418476 154398
rect 418540 154396 418546 154460
rect 421005 154458 421052 154460
rect 420960 154456 421052 154458
rect 420960 154400 421010 154456
rect 420960 154398 421052 154400
rect 421005 154396 421052 154398
rect 421116 154396 421122 154460
rect 425973 154458 426020 154460
rect 425928 154456 426020 154458
rect 425928 154400 425978 154456
rect 425928 154398 426020 154400
rect 425973 154396 426020 154398
rect 426084 154396 426090 154460
rect 443453 154458 443500 154460
rect 443408 154456 443500 154458
rect 443408 154400 443458 154456
rect 443408 154398 443500 154400
rect 443453 154396 443500 154398
rect 443564 154396 443570 154460
rect 418429 154395 418495 154396
rect 421005 154395 421071 154396
rect 425973 154395 426039 154396
rect 443453 154395 443519 154396
rect 138381 154324 138447 154325
rect 475837 154324 475903 154325
rect 478413 154324 478479 154325
rect 57830 154260 57836 154324
rect 57900 154322 57906 154324
rect 138381 154322 138428 154324
rect 57900 154262 122850 154322
rect 138336 154320 138428 154322
rect 138336 154264 138386 154320
rect 138336 154262 138428 154264
rect 57900 154260 57906 154262
rect 98453 154188 98519 154189
rect 101029 154188 101095 154189
rect 105813 154188 105879 154189
rect 108205 154188 108271 154189
rect 98453 154186 98500 154188
rect 98408 154184 98500 154186
rect 98408 154128 98458 154184
rect 98408 154126 98500 154128
rect 98453 154124 98500 154126
rect 98564 154124 98570 154188
rect 101029 154186 101076 154188
rect 100984 154184 101076 154186
rect 100984 154128 101034 154184
rect 100984 154126 101076 154128
rect 101029 154124 101076 154126
rect 101140 154124 101146 154188
rect 105813 154186 105860 154188
rect 105768 154184 105860 154186
rect 105768 154128 105818 154184
rect 105768 154126 105860 154128
rect 105813 154124 105860 154126
rect 105924 154124 105930 154188
rect 108205 154186 108252 154188
rect 108160 154184 108252 154186
rect 108160 154128 108210 154184
rect 108160 154126 108252 154128
rect 108205 154124 108252 154126
rect 108316 154124 108322 154188
rect 122790 154186 122850 154262
rect 138381 154260 138428 154262
rect 138492 154260 138498 154324
rect 208158 154260 208164 154324
rect 208228 154322 208234 154324
rect 313406 154322 313412 154324
rect 208228 154262 313412 154322
rect 208228 154260 208234 154262
rect 313406 154260 313412 154262
rect 313476 154260 313482 154324
rect 475837 154322 475884 154324
rect 475792 154320 475884 154322
rect 475792 154264 475842 154320
rect 475792 154262 475884 154264
rect 475837 154260 475884 154262
rect 475948 154260 475954 154324
rect 478413 154322 478460 154324
rect 478368 154320 478460 154322
rect 478368 154264 478418 154320
rect 478368 154262 478460 154264
rect 478413 154260 478460 154262
rect 478524 154260 478530 154324
rect 138381 154259 138447 154260
rect 475837 154259 475903 154260
rect 478413 154259 478479 154260
rect 143533 154188 143599 154189
rect 140814 154186 140820 154188
rect 122790 154126 140820 154186
rect 140814 154124 140820 154126
rect 140884 154124 140890 154188
rect 143533 154186 143580 154188
rect 143488 154184 143580 154186
rect 143488 154128 143538 154184
rect 143488 154126 143580 154128
rect 143533 154124 143580 154126
rect 143644 154124 143650 154188
rect 203006 154124 203012 154188
rect 203076 154186 203082 154188
rect 287973 154186 288039 154189
rect 288157 154188 288223 154189
rect 293309 154188 293375 154189
rect 473445 154188 473511 154189
rect 480805 154188 480871 154189
rect 288157 154186 288204 154188
rect 203076 154184 288039 154186
rect 203076 154128 287978 154184
rect 288034 154128 288039 154184
rect 203076 154126 288039 154128
rect 288112 154184 288204 154186
rect 288112 154128 288162 154184
rect 288112 154126 288204 154128
rect 203076 154124 203082 154126
rect 98453 154123 98519 154124
rect 101029 154123 101095 154124
rect 105813 154123 105879 154124
rect 108205 154123 108271 154124
rect 143533 154123 143599 154124
rect 287973 154123 288039 154126
rect 288157 154124 288204 154126
rect 288268 154124 288274 154188
rect 293309 154186 293356 154188
rect 293264 154184 293356 154186
rect 293264 154128 293314 154184
rect 293264 154126 293356 154128
rect 293309 154124 293356 154126
rect 293420 154124 293426 154188
rect 305862 154186 305868 154188
rect 296670 154126 305868 154186
rect 288157 154123 288223 154124
rect 293309 154123 293375 154124
rect 145925 154052 145991 154053
rect 150893 154052 150959 154053
rect 145925 154050 145972 154052
rect 145880 154048 145972 154050
rect 145880 153992 145930 154048
rect 145880 153990 145972 153992
rect 145925 153988 145972 153990
rect 146036 153988 146042 154052
rect 150893 154050 150940 154052
rect 150848 154048 150940 154050
rect 150848 153992 150898 154048
rect 150848 153990 150940 153992
rect 150893 153988 150940 153990
rect 151004 153988 151010 154052
rect 216070 153988 216076 154052
rect 216140 154050 216146 154052
rect 296670 154050 296730 154126
rect 305862 154124 305868 154126
rect 305932 154124 305938 154188
rect 473445 154186 473492 154188
rect 473400 154184 473492 154186
rect 473400 154128 473450 154184
rect 473400 154126 473492 154128
rect 473445 154124 473492 154126
rect 473556 154124 473562 154188
rect 480805 154186 480852 154188
rect 480760 154184 480852 154186
rect 480760 154128 480810 154184
rect 480760 154126 480852 154128
rect 480805 154124 480852 154126
rect 480916 154124 480922 154188
rect 473445 154123 473511 154124
rect 480805 154123 480871 154124
rect 298461 154052 298527 154053
rect 303429 154052 303495 154053
rect 470869 154052 470935 154053
rect 483197 154052 483263 154053
rect 298461 154050 298508 154052
rect 216140 153990 296730 154050
rect 298416 154048 298508 154050
rect 298416 153992 298466 154048
rect 298416 153990 298508 153992
rect 216140 153988 216146 153990
rect 298461 153988 298508 153990
rect 298572 153988 298578 154052
rect 303429 154050 303476 154052
rect 303384 154048 303476 154050
rect 303384 153992 303434 154048
rect 303384 153990 303476 153992
rect 303429 153988 303476 153990
rect 303540 153988 303546 154052
rect 470869 154050 470916 154052
rect 470824 154048 470916 154050
rect 470824 153992 470874 154048
rect 470824 153990 470916 153992
rect 470869 153988 470916 153990
rect 470980 153988 470986 154052
rect 483197 154050 483244 154052
rect 483152 154048 483244 154050
rect 483152 153992 483202 154048
rect 483152 153990 483244 153992
rect 483197 153988 483244 153990
rect 483308 153988 483314 154052
rect 145925 153987 145991 153988
rect 150893 153987 150959 153988
rect 298461 153987 298527 153988
rect 303429 153987 303495 153988
rect 470869 153987 470935 153988
rect 483197 153987 483263 153988
rect 153285 153916 153351 153917
rect 153285 153914 153332 153916
rect 153240 153912 153332 153914
rect 153240 153856 153290 153912
rect 153240 153854 153332 153856
rect 153285 153852 153332 153854
rect 153396 153852 153402 153916
rect 213126 153852 213132 153916
rect 213196 153914 213202 153916
rect 270902 153914 270908 153916
rect 213196 153854 270908 153914
rect 213196 153852 213202 153854
rect 270902 153852 270908 153854
rect 270972 153852 270978 153916
rect 287973 153914 288039 153917
rect 308397 153916 308463 153917
rect 423397 153916 423463 153917
rect 485957 153916 486023 153917
rect 295926 153914 295932 153916
rect 287973 153912 295932 153914
rect 287973 153856 287978 153912
rect 288034 153856 295932 153912
rect 287973 153854 295932 153856
rect 153285 153851 153351 153852
rect 287973 153851 288039 153854
rect 295926 153852 295932 153854
rect 295996 153852 296002 153916
rect 308397 153914 308444 153916
rect 308352 153912 308444 153914
rect 308352 153856 308402 153912
rect 308352 153854 308444 153856
rect 308397 153852 308444 153854
rect 308508 153852 308514 153916
rect 423397 153914 423444 153916
rect 423352 153912 423444 153914
rect 423352 153856 423402 153912
rect 423352 153854 423444 153856
rect 423397 153852 423444 153854
rect 423508 153852 423514 153916
rect 485957 153914 486004 153916
rect 485912 153912 486004 153914
rect 485912 153856 485962 153912
rect 485912 153854 486004 153856
rect 485957 153852 486004 153854
rect 486068 153852 486074 153916
rect 308397 153851 308463 153852
rect 423397 153851 423463 153852
rect 485957 153851 486023 153852
rect 85430 153172 85436 153236
rect 85500 153172 85506 153236
rect 95918 153172 95924 153236
rect 95988 153172 95994 153236
rect 99414 153172 99420 153236
rect 99484 153172 99490 153236
rect 236126 153172 236132 153236
rect 236196 153172 236202 153236
rect 261702 153172 261708 153236
rect 261772 153172 261778 153236
rect 265198 153172 265204 153236
rect 265268 153172 265274 153236
rect 272190 153172 272196 153236
rect 272260 153172 272266 153236
rect 300894 153172 300900 153236
rect 300964 153172 300970 153236
rect 398230 153172 398236 153236
rect 398300 153172 398306 153236
rect 401726 153172 401732 153236
rect 401796 153172 401802 153236
rect 416078 153172 416084 153236
rect 416148 153172 416154 153236
rect 455822 153172 455828 153236
rect 455892 153172 455898 153236
rect 463550 153172 463556 153236
rect 463620 153172 463626 153236
rect 75913 153098 75979 153101
rect 76046 153098 76052 153100
rect 75913 153096 76052 153098
rect 75913 153040 75918 153096
rect 75974 153040 76052 153096
rect 75913 153038 76052 153040
rect 75913 153035 75979 153038
rect 76046 153036 76052 153038
rect 76116 153036 76122 153100
rect 77293 153098 77359 153101
rect 78254 153098 78260 153100
rect 77293 153096 78260 153098
rect 77293 153040 77298 153096
rect 77354 153040 78260 153096
rect 77293 153038 78260 153040
rect 77293 153035 77359 153038
rect 78254 153036 78260 153038
rect 78324 153036 78330 153100
rect 78673 153098 78739 153101
rect 79542 153098 79548 153100
rect 78673 153096 79548 153098
rect 78673 153040 78678 153096
rect 78734 153040 79548 153096
rect 78673 153038 79548 153040
rect 78673 153035 78739 153038
rect 79542 153036 79548 153038
rect 79612 153036 79618 153100
rect 81433 153098 81499 153101
rect 81934 153098 81940 153100
rect 81433 153096 81940 153098
rect 81433 153040 81438 153096
rect 81494 153040 81940 153096
rect 81433 153038 81940 153040
rect 81433 153035 81499 153038
rect 81934 153036 81940 153038
rect 82004 153036 82010 153100
rect 82813 153098 82879 153101
rect 83038 153098 83044 153100
rect 82813 153096 83044 153098
rect 82813 153040 82818 153096
rect 82874 153040 83044 153096
rect 82813 153038 83044 153040
rect 82813 153035 82879 153038
rect 83038 153036 83044 153038
rect 83108 153036 83114 153100
rect 84193 153098 84259 153101
rect 85438 153098 85498 153172
rect 84193 153096 85498 153098
rect 84193 153040 84198 153096
rect 84254 153040 85498 153096
rect 84193 153038 85498 153040
rect 85573 153098 85639 153101
rect 86534 153098 86540 153100
rect 85573 153096 86540 153098
rect 85573 153040 85578 153096
rect 85634 153040 86540 153096
rect 85573 153038 86540 153040
rect 84193 153035 84259 153038
rect 85573 153035 85639 153038
rect 86534 153036 86540 153038
rect 86604 153036 86610 153100
rect 86953 153098 87019 153101
rect 87638 153098 87644 153100
rect 86953 153096 87644 153098
rect 86953 153040 86958 153096
rect 87014 153040 87644 153096
rect 86953 153038 87644 153040
rect 86953 153035 87019 153038
rect 87638 153036 87644 153038
rect 87708 153036 87714 153100
rect 88425 153098 88491 153101
rect 88742 153098 88748 153100
rect 88425 153096 88748 153098
rect 88425 153040 88430 153096
rect 88486 153040 88748 153096
rect 88425 153038 88748 153040
rect 88425 153035 88491 153038
rect 88742 153036 88748 153038
rect 88812 153036 88818 153100
rect 89805 153098 89871 153101
rect 90030 153098 90036 153100
rect 89805 153096 90036 153098
rect 89805 153040 89810 153096
rect 89866 153040 90036 153096
rect 89805 153038 90036 153040
rect 89805 153035 89871 153038
rect 90030 153036 90036 153038
rect 90100 153036 90106 153100
rect 91093 153098 91159 153101
rect 91318 153098 91324 153100
rect 91093 153096 91324 153098
rect 91093 153040 91098 153096
rect 91154 153040 91324 153096
rect 91093 153038 91324 153040
rect 91093 153035 91159 153038
rect 91318 153036 91324 153038
rect 91388 153036 91394 153100
rect 92473 153098 92539 153101
rect 93342 153098 93348 153100
rect 92473 153096 93348 153098
rect 92473 153040 92478 153096
rect 92534 153040 93348 153096
rect 92473 153038 93348 153040
rect 92473 153035 92539 153038
rect 93342 153036 93348 153038
rect 93412 153036 93418 153100
rect 93853 153098 93919 153101
rect 94446 153098 94452 153100
rect 93853 153096 94452 153098
rect 93853 153040 93858 153096
rect 93914 153040 94452 153096
rect 93853 153038 94452 153040
rect 93853 153035 93919 153038
rect 94446 153036 94452 153038
rect 94516 153036 94522 153100
rect 95233 153098 95299 153101
rect 95926 153098 95986 153172
rect 99422 153101 99482 153172
rect 236134 153101 236194 153172
rect 95233 153096 95986 153098
rect 95233 153040 95238 153096
rect 95294 153040 95986 153096
rect 95233 153038 95986 153040
rect 96613 153098 96679 153101
rect 97022 153098 97028 153100
rect 96613 153096 97028 153098
rect 96613 153040 96618 153096
rect 96674 153040 97028 153096
rect 96613 153038 97028 153040
rect 95233 153035 95299 153038
rect 96613 153035 96679 153038
rect 97022 153036 97028 153038
rect 97092 153036 97098 153100
rect 97993 153098 98059 153101
rect 98126 153098 98132 153100
rect 97993 153096 98132 153098
rect 97993 153040 97998 153096
rect 98054 153040 98132 153096
rect 97993 153038 98132 153040
rect 97993 153035 98059 153038
rect 98126 153036 98132 153038
rect 98196 153036 98202 153100
rect 99373 153096 99482 153101
rect 99373 153040 99378 153096
rect 99434 153040 99482 153096
rect 99373 153038 99482 153040
rect 99373 153035 99439 153038
rect 100702 153036 100708 153100
rect 100772 153098 100778 153100
rect 100845 153098 100911 153101
rect 100772 153096 100911 153098
rect 100772 153040 100850 153096
rect 100906 153040 100911 153096
rect 100772 153038 100911 153040
rect 100772 153036 100778 153038
rect 100845 153035 100911 153038
rect 102133 153098 102199 153101
rect 102726 153098 102732 153100
rect 102133 153096 102732 153098
rect 102133 153040 102138 153096
rect 102194 153040 102732 153096
rect 102133 153038 102732 153040
rect 102133 153035 102199 153038
rect 102726 153036 102732 153038
rect 102796 153036 102802 153100
rect 103605 153098 103671 153101
rect 106365 153100 106431 153101
rect 103830 153098 103836 153100
rect 103605 153096 103836 153098
rect 103605 153040 103610 153096
rect 103666 153040 103836 153096
rect 103605 153038 103836 153040
rect 103605 153035 103671 153038
rect 103830 153036 103836 153038
rect 103900 153036 103906 153100
rect 106365 153098 106412 153100
rect 106320 153096 106412 153098
rect 106320 153040 106370 153096
rect 106320 153038 106412 153040
rect 106365 153036 106412 153038
rect 106476 153036 106482 153100
rect 108798 153036 108804 153100
rect 108868 153098 108874 153100
rect 109033 153098 109099 153101
rect 108868 153096 109099 153098
rect 108868 153040 109038 153096
rect 109094 153040 109099 153096
rect 108868 153038 109099 153040
rect 108868 153036 108874 153038
rect 106365 153035 106431 153036
rect 109033 153035 109099 153038
rect 110413 153098 110479 153101
rect 111149 153100 111215 153101
rect 111006 153098 111012 153100
rect 110413 153096 111012 153098
rect 110413 153040 110418 153096
rect 110474 153040 111012 153096
rect 110413 153038 111012 153040
rect 110413 153035 110479 153038
rect 111006 153036 111012 153038
rect 111076 153036 111082 153100
rect 111149 153096 111196 153100
rect 111260 153098 111266 153100
rect 111793 153098 111859 153101
rect 114553 153100 114619 153101
rect 112110 153098 112116 153100
rect 111149 153040 111154 153096
rect 111149 153036 111196 153040
rect 111260 153038 111306 153098
rect 111793 153096 112116 153098
rect 111793 153040 111798 153096
rect 111854 153040 112116 153096
rect 111793 153038 112116 153040
rect 111260 153036 111266 153038
rect 111149 153035 111215 153036
rect 111793 153035 111859 153038
rect 112110 153036 112116 153038
rect 112180 153036 112186 153100
rect 114502 153036 114508 153100
rect 114572 153098 114619 153100
rect 114737 153098 114803 153101
rect 115790 153098 115796 153100
rect 114572 153096 114664 153098
rect 114614 153040 114664 153096
rect 114572 153038 114664 153040
rect 114737 153096 115796 153098
rect 114737 153040 114742 153096
rect 114798 153040 115796 153096
rect 114737 153038 115796 153040
rect 114572 153036 114619 153038
rect 114553 153035 114619 153036
rect 114737 153035 114803 153038
rect 115790 153036 115796 153038
rect 115860 153036 115866 153100
rect 117078 153036 117084 153100
rect 117148 153098 117154 153100
rect 117313 153098 117379 153101
rect 117148 153096 117379 153098
rect 117148 153040 117318 153096
rect 117374 153040 117379 153096
rect 117148 153038 117379 153040
rect 117148 153036 117154 153038
rect 117313 153035 117379 153038
rect 117497 153098 117563 153101
rect 118366 153098 118372 153100
rect 117497 153096 118372 153098
rect 117497 153040 117502 153096
rect 117558 153040 118372 153096
rect 117497 153038 118372 153040
rect 117497 153035 117563 153038
rect 118366 153036 118372 153038
rect 118436 153036 118442 153100
rect 118693 153098 118759 153101
rect 119102 153098 119108 153100
rect 118693 153096 119108 153098
rect 118693 153040 118698 153096
rect 118754 153040 119108 153096
rect 118693 153038 119108 153040
rect 118693 153035 118759 153038
rect 119102 153036 119108 153038
rect 119172 153036 119178 153100
rect 125593 153098 125659 153101
rect 125910 153098 125916 153100
rect 125593 153096 125916 153098
rect 125593 153040 125598 153096
rect 125654 153040 125916 153096
rect 125593 153038 125916 153040
rect 125593 153035 125659 153038
rect 125910 153036 125916 153038
rect 125980 153036 125986 153100
rect 128353 153098 128419 153101
rect 128486 153098 128492 153100
rect 128353 153096 128492 153098
rect 128353 153040 128358 153096
rect 128414 153040 128492 153096
rect 128353 153038 128492 153040
rect 128353 153035 128419 153038
rect 128486 153036 128492 153038
rect 128556 153036 128562 153100
rect 129733 153098 129799 153101
rect 130878 153098 130884 153100
rect 129733 153096 130884 153098
rect 129733 153040 129738 153096
rect 129794 153040 130884 153096
rect 129733 153038 130884 153040
rect 129733 153035 129799 153038
rect 130878 153036 130884 153038
rect 130948 153036 130954 153100
rect 132769 153098 132835 153101
rect 133454 153098 133460 153100
rect 132769 153096 133460 153098
rect 132769 153040 132774 153096
rect 132830 153040 133460 153096
rect 132769 153038 133460 153040
rect 132769 153035 132835 153038
rect 133454 153036 133460 153038
rect 133524 153036 133530 153100
rect 135253 153098 135319 153101
rect 155953 153100 156019 153101
rect 136030 153098 136036 153100
rect 135253 153096 136036 153098
rect 135253 153040 135258 153096
rect 135314 153040 136036 153096
rect 135253 153038 136036 153040
rect 135253 153035 135319 153038
rect 136030 153036 136036 153038
rect 136100 153036 136106 153100
rect 155902 153036 155908 153100
rect 155972 153098 156019 153100
rect 218237 153098 218303 153101
rect 218646 153098 218652 153100
rect 155972 153096 156064 153098
rect 156014 153040 156064 153096
rect 155972 153038 156064 153040
rect 218237 153096 218652 153098
rect 218237 153040 218242 153096
rect 218298 153040 218652 153096
rect 218237 153038 218652 153040
rect 155972 153036 156019 153038
rect 155953 153035 156019 153036
rect 218237 153035 218303 153038
rect 218646 153036 218652 153038
rect 218716 153036 218722 153100
rect 236085 153096 236194 153101
rect 236085 153040 236090 153096
rect 236146 153040 236194 153096
rect 236085 153038 236194 153040
rect 237373 153098 237439 153101
rect 238150 153098 238156 153100
rect 237373 153096 238156 153098
rect 237373 153040 237378 153096
rect 237434 153040 238156 153096
rect 237373 153038 238156 153040
rect 236085 153035 236151 153038
rect 237373 153035 237439 153038
rect 238150 153036 238156 153038
rect 238220 153036 238226 153100
rect 240133 153098 240199 153101
rect 240542 153098 240548 153100
rect 240133 153096 240548 153098
rect 240133 153040 240138 153096
rect 240194 153040 240548 153096
rect 240133 153038 240548 153040
rect 240133 153035 240199 153038
rect 240542 153036 240548 153038
rect 240612 153036 240618 153100
rect 241513 153098 241579 153101
rect 242893 153100 242959 153101
rect 244273 153100 244339 153101
rect 241646 153098 241652 153100
rect 241513 153096 241652 153098
rect 241513 153040 241518 153096
rect 241574 153040 241652 153096
rect 241513 153038 241652 153040
rect 241513 153035 241579 153038
rect 241646 153036 241652 153038
rect 241716 153036 241722 153100
rect 242893 153098 242940 153100
rect 242848 153096 242940 153098
rect 242848 153040 242898 153096
rect 242848 153038 242940 153040
rect 242893 153036 242940 153038
rect 243004 153036 243010 153100
rect 244222 153036 244228 153100
rect 244292 153098 244339 153100
rect 245653 153098 245719 153101
rect 246430 153098 246436 153100
rect 244292 153096 244384 153098
rect 244334 153040 244384 153096
rect 244292 153038 244384 153040
rect 245653 153096 246436 153098
rect 245653 153040 245658 153096
rect 245714 153040 246436 153096
rect 245653 153038 246436 153040
rect 244292 153036 244339 153038
rect 242893 153035 242959 153036
rect 244273 153035 244339 153036
rect 245653 153035 245719 153038
rect 246430 153036 246436 153038
rect 246500 153036 246506 153100
rect 247033 153098 247099 153101
rect 247718 153098 247724 153100
rect 247033 153096 247724 153098
rect 247033 153040 247038 153096
rect 247094 153040 247724 153096
rect 247033 153038 247724 153040
rect 247033 153035 247099 153038
rect 247718 153036 247724 153038
rect 247788 153036 247794 153100
rect 248413 153098 248479 153101
rect 248638 153098 248644 153100
rect 248413 153096 248644 153098
rect 248413 153040 248418 153096
rect 248474 153040 248644 153096
rect 248413 153038 248644 153040
rect 248413 153035 248479 153038
rect 248638 153036 248644 153038
rect 248708 153036 248714 153100
rect 249793 153098 249859 153101
rect 250110 153098 250116 153100
rect 249793 153096 250116 153098
rect 249793 153040 249798 153096
rect 249854 153040 250116 153096
rect 249793 153038 250116 153040
rect 249793 153035 249859 153038
rect 250110 153036 250116 153038
rect 250180 153036 250186 153100
rect 250253 153098 250319 153101
rect 251173 153100 251239 153101
rect 250662 153098 250668 153100
rect 250253 153096 250668 153098
rect 250253 153040 250258 153096
rect 250314 153040 250668 153096
rect 250253 153038 250668 153040
rect 250253 153035 250319 153038
rect 250662 153036 250668 153038
rect 250732 153036 250738 153100
rect 251173 153098 251220 153100
rect 251128 153096 251220 153098
rect 251128 153040 251178 153096
rect 251128 153038 251220 153040
rect 251173 153036 251220 153038
rect 251284 153036 251290 153100
rect 252553 153098 252619 153101
rect 253565 153100 253631 153101
rect 253422 153098 253428 153100
rect 252553 153096 253428 153098
rect 252553 153040 252558 153096
rect 252614 153040 253428 153096
rect 252553 153038 253428 153040
rect 251173 153035 251239 153036
rect 252553 153035 252619 153038
rect 253422 153036 253428 153038
rect 253492 153036 253498 153100
rect 253565 153096 253612 153100
rect 253676 153098 253682 153100
rect 253933 153098 253999 153101
rect 254526 153098 254532 153100
rect 253565 153040 253570 153096
rect 253565 153036 253612 153040
rect 253676 153038 253722 153098
rect 253933 153096 254532 153098
rect 253933 153040 253938 153096
rect 253994 153040 254532 153096
rect 253933 153038 254532 153040
rect 253676 153036 253682 153038
rect 253565 153035 253631 153036
rect 253933 153035 253999 153038
rect 254526 153036 254532 153038
rect 254596 153036 254602 153100
rect 255313 153098 255379 153101
rect 255814 153098 255820 153100
rect 255313 153096 255820 153098
rect 255313 153040 255318 153096
rect 255374 153040 255820 153096
rect 255313 153038 255820 153040
rect 255313 153035 255379 153038
rect 255814 153036 255820 153038
rect 255884 153036 255890 153100
rect 255957 153098 256023 153101
rect 256182 153098 256188 153100
rect 255957 153096 256188 153098
rect 255957 153040 255962 153096
rect 256018 153040 256188 153096
rect 255957 153038 256188 153040
rect 255957 153035 256023 153038
rect 256182 153036 256188 153038
rect 256252 153036 256258 153100
rect 256693 153098 256759 153101
rect 256918 153098 256924 153100
rect 256693 153096 256924 153098
rect 256693 153040 256698 153096
rect 256754 153040 256924 153096
rect 256693 153038 256924 153040
rect 256693 153035 256759 153038
rect 256918 153036 256924 153038
rect 256988 153036 256994 153100
rect 258073 153098 258139 153101
rect 259545 153100 259611 153101
rect 258206 153098 258212 153100
rect 258073 153096 258212 153098
rect 258073 153040 258078 153096
rect 258134 153040 258212 153096
rect 258073 153038 258212 153040
rect 258073 153035 258139 153038
rect 258206 153036 258212 153038
rect 258276 153036 258282 153100
rect 259494 153036 259500 153100
rect 259564 153098 259611 153100
rect 261201 153098 261267 153101
rect 261710 153098 261770 153172
rect 259564 153096 259656 153098
rect 259606 153040 259656 153096
rect 259564 153038 259656 153040
rect 261201 153096 261770 153098
rect 261201 153040 261206 153096
rect 261262 153040 261770 153096
rect 261201 153038 261770 153040
rect 262213 153098 262279 153101
rect 262806 153098 262812 153100
rect 262213 153096 262812 153098
rect 262213 153040 262218 153096
rect 262274 153040 262812 153096
rect 262213 153038 262812 153040
rect 259564 153036 259611 153038
rect 259545 153035 259611 153036
rect 261201 153035 261267 153038
rect 262213 153035 262279 153038
rect 262806 153036 262812 153038
rect 262876 153036 262882 153100
rect 263593 153098 263659 153101
rect 263910 153098 263916 153100
rect 263593 153096 263916 153098
rect 263593 153040 263598 153096
rect 263654 153040 263916 153096
rect 263593 153038 263916 153040
rect 263593 153035 263659 153038
rect 263910 153036 263916 153038
rect 263980 153036 263986 153100
rect 264973 153098 265039 153101
rect 265206 153098 265266 153172
rect 266353 153100 266419 153101
rect 264973 153096 265266 153098
rect 264973 153040 264978 153096
rect 265034 153040 265266 153096
rect 264973 153038 265266 153040
rect 264973 153035 265039 153038
rect 266302 153036 266308 153100
rect 266372 153098 266419 153100
rect 267733 153098 267799 153101
rect 268694 153098 268700 153100
rect 266372 153096 266464 153098
rect 266414 153040 266464 153096
rect 266372 153038 266464 153040
rect 267733 153096 268700 153098
rect 267733 153040 267738 153096
rect 267794 153040 268700 153096
rect 267733 153038 268700 153040
rect 266372 153036 266419 153038
rect 266353 153035 266419 153036
rect 267733 153035 267799 153038
rect 268694 153036 268700 153038
rect 268764 153036 268770 153100
rect 269113 153098 269179 153101
rect 269798 153098 269804 153100
rect 269113 153096 269804 153098
rect 269113 153040 269118 153096
rect 269174 153040 269804 153096
rect 269113 153038 269804 153040
rect 269113 153035 269179 153038
rect 269798 153036 269804 153038
rect 269868 153036 269874 153100
rect 270493 153098 270559 153101
rect 271086 153098 271092 153100
rect 270493 153096 271092 153098
rect 270493 153040 270498 153096
rect 270554 153040 271092 153096
rect 270493 153038 271092 153040
rect 270493 153035 270559 153038
rect 271086 153036 271092 153038
rect 271156 153036 271162 153100
rect 271873 153098 271939 153101
rect 272198 153098 272258 153172
rect 300902 153101 300962 153172
rect 271873 153096 272258 153098
rect 271873 153040 271878 153096
rect 271934 153040 272258 153096
rect 271873 153038 272258 153040
rect 273253 153098 273319 153101
rect 274398 153098 274404 153100
rect 273253 153096 274404 153098
rect 273253 153040 273258 153096
rect 273314 153040 274404 153096
rect 273253 153038 274404 153040
rect 271873 153035 271939 153038
rect 273253 153035 273319 153038
rect 274398 153036 274404 153038
rect 274468 153036 274474 153100
rect 274725 153098 274791 153101
rect 275318 153098 275324 153100
rect 274725 153096 275324 153098
rect 274725 153040 274730 153096
rect 274786 153040 275324 153096
rect 274725 153038 275324 153040
rect 274725 153035 274791 153038
rect 275318 153036 275324 153038
rect 275388 153036 275394 153100
rect 277945 153098 278011 153101
rect 278446 153098 278452 153100
rect 277945 153096 278452 153098
rect 277945 153040 277950 153096
rect 278006 153040 278452 153096
rect 277945 153038 278452 153040
rect 277945 153035 278011 153038
rect 278446 153036 278452 153038
rect 278516 153036 278522 153100
rect 278998 153036 279004 153100
rect 279068 153098 279074 153100
rect 280061 153098 280127 153101
rect 279068 153096 280127 153098
rect 279068 153040 280066 153096
rect 280122 153040 280127 153096
rect 279068 153038 280127 153040
rect 279068 153036 279074 153038
rect 280061 153035 280127 153038
rect 280245 153098 280311 153101
rect 280838 153098 280844 153100
rect 280245 153096 280844 153098
rect 280245 153040 280250 153096
rect 280306 153040 280844 153096
rect 280245 153038 280844 153040
rect 280245 153035 280311 153038
rect 280838 153036 280844 153038
rect 280908 153036 280914 153100
rect 282913 153098 282979 153101
rect 283782 153098 283788 153100
rect 282913 153096 283788 153098
rect 282913 153040 282918 153096
rect 282974 153040 283788 153096
rect 282913 153038 283788 153040
rect 282913 153035 282979 153038
rect 283782 153036 283788 153038
rect 283852 153036 283858 153100
rect 285673 153098 285739 153101
rect 285990 153098 285996 153100
rect 285673 153096 285996 153098
rect 285673 153040 285678 153096
rect 285734 153040 285996 153096
rect 285673 153038 285996 153040
rect 285673 153035 285739 153038
rect 285990 153036 285996 153038
rect 286060 153036 286066 153100
rect 289813 153098 289879 153101
rect 290958 153098 290964 153100
rect 289813 153096 290964 153098
rect 289813 153040 289818 153096
rect 289874 153040 290964 153096
rect 289813 153038 290964 153040
rect 289813 153035 289879 153038
rect 290958 153036 290964 153038
rect 291028 153036 291034 153100
rect 300853 153096 300962 153101
rect 300853 153040 300858 153096
rect 300914 153040 300962 153096
rect 300853 153038 300962 153040
rect 320173 153098 320239 153101
rect 396073 153100 396139 153101
rect 320950 153098 320956 153100
rect 320173 153096 320956 153098
rect 320173 153040 320178 153096
rect 320234 153040 320956 153096
rect 320173 153038 320956 153040
rect 300853 153035 300919 153038
rect 320173 153035 320239 153038
rect 320950 153036 320956 153038
rect 321020 153036 321026 153100
rect 396022 153036 396028 153100
rect 396092 153098 396139 153100
rect 397453 153098 397519 153101
rect 398238 153098 398298 153172
rect 396092 153096 396184 153098
rect 396134 153040 396184 153096
rect 396092 153038 396184 153040
rect 397453 153096 398298 153098
rect 397453 153040 397458 153096
rect 397514 153040 398298 153096
rect 397453 153038 398298 153040
rect 398833 153098 398899 153101
rect 399518 153098 399524 153100
rect 398833 153096 399524 153098
rect 398833 153040 398838 153096
rect 398894 153040 399524 153096
rect 398833 153038 399524 153040
rect 396092 153036 396139 153038
rect 396073 153035 396139 153036
rect 397453 153035 397519 153038
rect 398833 153035 398899 153038
rect 399518 153036 399524 153038
rect 399588 153036 399594 153100
rect 400213 153098 400279 153101
rect 400438 153098 400444 153100
rect 400213 153096 400444 153098
rect 400213 153040 400218 153096
rect 400274 153040 400444 153096
rect 400213 153038 400444 153040
rect 400213 153035 400279 153038
rect 400438 153036 400444 153038
rect 400508 153036 400514 153100
rect 401593 153098 401659 153101
rect 401734 153098 401794 153172
rect 403065 153100 403131 153101
rect 401593 153096 401794 153098
rect 401593 153040 401598 153096
rect 401654 153040 401794 153096
rect 401593 153038 401794 153040
rect 401593 153035 401659 153038
rect 403014 153036 403020 153100
rect 403084 153098 403131 153100
rect 404353 153098 404419 153101
rect 405038 153098 405044 153100
rect 403084 153096 403176 153098
rect 403126 153040 403176 153096
rect 403084 153038 403176 153040
rect 404353 153096 405044 153098
rect 404353 153040 404358 153096
rect 404414 153040 405044 153096
rect 404353 153038 405044 153040
rect 403084 153036 403131 153038
rect 403065 153035 403131 153036
rect 404353 153035 404419 153038
rect 405038 153036 405044 153038
rect 405108 153036 405114 153100
rect 405733 153098 405799 153101
rect 406510 153098 406516 153100
rect 405733 153096 406516 153098
rect 405733 153040 405738 153096
rect 405794 153040 406516 153096
rect 405733 153038 406516 153040
rect 405733 153035 405799 153038
rect 406510 153036 406516 153038
rect 406580 153036 406586 153100
rect 407205 153098 407271 153101
rect 407614 153098 407620 153100
rect 407205 153096 407620 153098
rect 407205 153040 407210 153096
rect 407266 153040 407620 153096
rect 407205 153038 407620 153040
rect 407205 153035 407271 153038
rect 407614 153036 407620 153038
rect 407684 153036 407690 153100
rect 408493 153098 408559 153101
rect 409965 153100 410031 153101
rect 411345 153100 411411 153101
rect 408718 153098 408724 153100
rect 408493 153096 408724 153098
rect 408493 153040 408498 153096
rect 408554 153040 408724 153096
rect 408493 153038 408724 153040
rect 408493 153035 408559 153038
rect 408718 153036 408724 153038
rect 408788 153036 408794 153100
rect 409965 153098 410012 153100
rect 409920 153096 410012 153098
rect 409920 153040 409970 153096
rect 409920 153038 410012 153040
rect 409965 153036 410012 153038
rect 410076 153036 410082 153100
rect 411294 153036 411300 153100
rect 411364 153098 411411 153100
rect 412725 153098 412791 153101
rect 413502 153098 413508 153100
rect 411364 153096 411456 153098
rect 411406 153040 411456 153096
rect 411364 153038 411456 153040
rect 412725 153096 413508 153098
rect 412725 153040 412730 153096
rect 412786 153040 413508 153096
rect 412725 153038 413508 153040
rect 411364 153036 411411 153038
rect 409965 153035 410031 153036
rect 411345 153035 411411 153036
rect 412725 153035 412791 153038
rect 413502 153036 413508 153038
rect 413572 153036 413578 153100
rect 414013 153098 414079 153101
rect 415485 153100 415551 153101
rect 414422 153098 414428 153100
rect 414013 153096 414428 153098
rect 414013 153040 414018 153096
rect 414074 153040 414428 153096
rect 414013 153038 414428 153040
rect 414013 153035 414079 153038
rect 414422 153036 414428 153038
rect 414492 153036 414498 153100
rect 415485 153098 415532 153100
rect 415440 153096 415532 153098
rect 415440 153040 415490 153096
rect 415440 153038 415532 153040
rect 415485 153036 415532 153038
rect 415596 153036 415602 153100
rect 415669 153098 415735 153101
rect 416086 153098 416146 153172
rect 415669 153096 416146 153098
rect 415669 153040 415674 153096
rect 415730 153040 416146 153096
rect 415669 153038 416146 153040
rect 416773 153098 416839 153101
rect 416998 153098 417004 153100
rect 416773 153096 417004 153098
rect 416773 153040 416778 153096
rect 416834 153040 417004 153096
rect 416773 153038 417004 153040
rect 415485 153035 415551 153036
rect 415669 153035 415735 153038
rect 416773 153035 416839 153038
rect 416998 153036 417004 153038
rect 417068 153036 417074 153100
rect 418102 153036 418108 153100
rect 418172 153098 418178 153100
rect 418245 153098 418311 153101
rect 418172 153096 418311 153098
rect 418172 153040 418250 153096
rect 418306 153040 418311 153096
rect 418172 153038 418311 153040
rect 418172 153036 418178 153038
rect 418245 153035 418311 153038
rect 419533 153098 419599 153101
rect 420678 153098 420684 153100
rect 419533 153096 420684 153098
rect 419533 153040 419538 153096
rect 419594 153040 420684 153096
rect 419533 153038 420684 153040
rect 419533 153035 419599 153038
rect 420678 153036 420684 153038
rect 420748 153036 420754 153100
rect 420913 153098 420979 153101
rect 421782 153098 421788 153100
rect 420913 153096 421788 153098
rect 420913 153040 420918 153096
rect 420974 153040 421788 153096
rect 420913 153038 421788 153040
rect 420913 153035 420979 153038
rect 421782 153036 421788 153038
rect 421852 153036 421858 153100
rect 422293 153098 422359 153101
rect 422886 153098 422892 153100
rect 422293 153096 422892 153098
rect 422293 153040 422298 153096
rect 422354 153040 422892 153096
rect 422293 153038 422892 153040
rect 422293 153035 422359 153038
rect 422886 153036 422892 153038
rect 422956 153036 422962 153100
rect 423673 153098 423739 153101
rect 423990 153098 423996 153100
rect 423673 153096 423996 153098
rect 423673 153040 423678 153096
rect 423734 153040 423996 153096
rect 423673 153038 423996 153040
rect 423673 153035 423739 153038
rect 423990 153036 423996 153038
rect 424060 153036 424066 153100
rect 425053 153098 425119 153101
rect 425278 153098 425284 153100
rect 425053 153096 425284 153098
rect 425053 153040 425058 153096
rect 425114 153040 425284 153096
rect 425053 153038 425284 153040
rect 425053 153035 425119 153038
rect 425278 153036 425284 153038
rect 425348 153036 425354 153100
rect 426382 153036 426388 153100
rect 426452 153098 426458 153100
rect 426525 153098 426591 153101
rect 426452 153096 426591 153098
rect 426452 153040 426530 153096
rect 426586 153040 426591 153096
rect 426452 153038 426591 153040
rect 426452 153036 426458 153038
rect 426525 153035 426591 153038
rect 427813 153098 427879 153101
rect 428590 153098 428596 153100
rect 427813 153096 428596 153098
rect 427813 153040 427818 153096
rect 427874 153040 428596 153096
rect 427813 153038 428596 153040
rect 427813 153035 427879 153038
rect 428590 153036 428596 153038
rect 428660 153036 428666 153100
rect 429193 153098 429259 153101
rect 429694 153098 429700 153100
rect 429193 153096 429700 153098
rect 429193 153040 429198 153096
rect 429254 153040 429700 153096
rect 429193 153038 429700 153040
rect 429193 153035 429259 153038
rect 429694 153036 429700 153038
rect 429764 153036 429770 153100
rect 430573 153098 430639 153101
rect 431166 153098 431172 153100
rect 430573 153096 431172 153098
rect 430573 153040 430578 153096
rect 430634 153040 431172 153096
rect 430573 153038 431172 153040
rect 430573 153035 430639 153038
rect 431166 153036 431172 153038
rect 431236 153036 431242 153100
rect 431718 153036 431724 153100
rect 431788 153098 431794 153100
rect 431953 153098 432019 153101
rect 431788 153096 432019 153098
rect 431788 153040 431958 153096
rect 432014 153040 432019 153096
rect 431788 153038 432019 153040
rect 431788 153036 431794 153038
rect 431953 153035 432019 153038
rect 433333 153098 433399 153101
rect 433558 153098 433564 153100
rect 433333 153096 433564 153098
rect 433333 153040 433338 153096
rect 433394 153040 433564 153096
rect 433333 153038 433564 153040
rect 433333 153035 433399 153038
rect 433558 153036 433564 153038
rect 433628 153036 433634 153100
rect 433977 153098 434043 153101
rect 434662 153098 434668 153100
rect 433977 153096 434668 153098
rect 433977 153040 433982 153096
rect 434038 153040 434668 153096
rect 433977 153038 434668 153040
rect 433977 153035 434043 153038
rect 434662 153036 434668 153038
rect 434732 153036 434738 153100
rect 434805 153098 434871 153101
rect 435950 153098 435956 153100
rect 434805 153096 435956 153098
rect 434805 153040 434810 153096
rect 434866 153040 435956 153096
rect 434805 153038 435956 153040
rect 434805 153035 434871 153038
rect 435950 153036 435956 153038
rect 436020 153036 436026 153100
rect 436185 153098 436251 153101
rect 436870 153098 436876 153100
rect 436185 153096 436876 153098
rect 436185 153040 436190 153096
rect 436246 153040 436876 153096
rect 436185 153038 436876 153040
rect 436185 153035 436251 153038
rect 436870 153036 436876 153038
rect 436940 153036 436946 153100
rect 438342 153036 438348 153100
rect 438412 153098 438418 153100
rect 438853 153098 438919 153101
rect 438412 153096 438919 153098
rect 438412 153040 438858 153096
rect 438914 153040 438919 153096
rect 438412 153038 438919 153040
rect 438412 153036 438418 153038
rect 438853 153035 438919 153038
rect 439262 153036 439268 153100
rect 439332 153098 439338 153100
rect 440141 153098 440207 153101
rect 439332 153096 440207 153098
rect 439332 153040 440146 153096
rect 440202 153040 440207 153096
rect 439332 153038 440207 153040
rect 439332 153036 439338 153038
rect 440141 153035 440207 153038
rect 440325 153098 440391 153101
rect 440918 153098 440924 153100
rect 440325 153096 440924 153098
rect 440325 153040 440330 153096
rect 440386 153040 440924 153096
rect 440325 153038 440924 153040
rect 440325 153035 440391 153038
rect 440918 153036 440924 153038
rect 440988 153036 440994 153100
rect 445753 153098 445819 153101
rect 445886 153098 445892 153100
rect 445753 153096 445892 153098
rect 445753 153040 445758 153096
rect 445814 153040 445892 153096
rect 445753 153038 445892 153040
rect 445753 153035 445819 153038
rect 445886 153036 445892 153038
rect 445956 153036 445962 153100
rect 447133 153098 447199 153101
rect 448278 153098 448284 153100
rect 447133 153096 448284 153098
rect 447133 153040 447138 153096
rect 447194 153040 448284 153096
rect 447133 153038 448284 153040
rect 447133 153035 447199 153038
rect 448278 153036 448284 153038
rect 448348 153036 448354 153100
rect 449893 153098 449959 153101
rect 451038 153098 451044 153100
rect 449893 153096 451044 153098
rect 449893 153040 449898 153096
rect 449954 153040 451044 153096
rect 449893 153038 451044 153040
rect 449893 153035 449959 153038
rect 451038 153036 451044 153038
rect 451108 153036 451114 153100
rect 452653 153098 452719 153101
rect 453430 153098 453436 153100
rect 452653 153096 453436 153098
rect 452653 153040 452658 153096
rect 452714 153040 453436 153096
rect 452653 153038 453436 153040
rect 452653 153035 452719 153038
rect 453430 153036 453436 153038
rect 453500 153036 453506 153100
rect 455413 153098 455479 153101
rect 455830 153098 455890 153172
rect 455413 153096 455890 153098
rect 455413 153040 455418 153096
rect 455474 153040 455890 153096
rect 455413 153038 455890 153040
rect 458173 153098 458239 153101
rect 458398 153098 458404 153100
rect 458173 153096 458404 153098
rect 458173 153040 458178 153096
rect 458234 153040 458404 153096
rect 458173 153038 458404 153040
rect 455413 153035 455479 153038
rect 458173 153035 458239 153038
rect 458398 153036 458404 153038
rect 458468 153036 458474 153100
rect 49417 152962 49483 152965
rect 158478 152962 158484 152964
rect 49417 152960 158484 152962
rect 49417 152904 49422 152960
rect 49478 152904 158484 152960
rect 49417 152902 158484 152904
rect 49417 152899 49483 152902
rect 158478 152900 158484 152902
rect 158548 152900 158554 152964
rect 206502 152900 206508 152964
rect 206572 152962 206578 152964
rect 318374 152962 318380 152964
rect 206572 152902 318380 152962
rect 206572 152900 206578 152902
rect 318374 152900 318380 152902
rect 318444 152900 318450 152964
rect 370589 152962 370655 152965
rect 463558 152962 463618 153172
rect 370589 152960 463618 152962
rect 370589 152904 370594 152960
rect 370650 152904 463618 152960
rect 370589 152902 463618 152904
rect 370589 152899 370655 152902
rect 48078 152764 48084 152828
rect 48148 152826 48154 152828
rect 88885 152826 88951 152829
rect 48148 152824 88951 152826
rect 48148 152768 88890 152824
rect 88946 152768 88951 152824
rect 48148 152766 88951 152768
rect 48148 152764 48154 152766
rect 88885 152763 88951 152766
rect 91185 152826 91251 152829
rect 91502 152826 91508 152828
rect 91185 152824 91508 152826
rect 91185 152768 91190 152824
rect 91246 152768 91508 152824
rect 91185 152766 91508 152768
rect 91185 152763 91251 152766
rect 91502 152764 91508 152766
rect 91572 152764 91578 152828
rect 100753 152826 100819 152829
rect 101806 152826 101812 152828
rect 100753 152824 101812 152826
rect 100753 152768 100758 152824
rect 100814 152768 101812 152824
rect 100753 152766 101812 152768
rect 100753 152763 100819 152766
rect 101806 152764 101812 152766
rect 101876 152764 101882 152828
rect 103513 152826 103579 152829
rect 103830 152826 103836 152828
rect 103513 152824 103836 152826
rect 103513 152768 103518 152824
rect 103574 152768 103836 152824
rect 103513 152766 103836 152768
rect 103513 152763 103579 152766
rect 103830 152764 103836 152766
rect 103900 152764 103906 152828
rect 106273 152826 106339 152829
rect 107510 152826 107516 152828
rect 106273 152824 107516 152826
rect 106273 152768 106278 152824
rect 106334 152768 107516 152824
rect 106273 152766 107516 152768
rect 106273 152763 106339 152766
rect 107510 152764 107516 152766
rect 107580 152764 107586 152828
rect 109125 152826 109191 152829
rect 113173 152828 113239 152829
rect 109534 152826 109540 152828
rect 109125 152824 109540 152826
rect 109125 152768 109130 152824
rect 109186 152768 109540 152824
rect 109125 152766 109540 152768
rect 109125 152763 109191 152766
rect 109534 152764 109540 152766
rect 109604 152764 109610 152828
rect 113173 152824 113220 152828
rect 113284 152826 113290 152828
rect 117405 152826 117471 152829
rect 117998 152826 118004 152828
rect 113173 152768 113178 152824
rect 113173 152764 113220 152768
rect 113284 152766 113330 152826
rect 117405 152824 118004 152826
rect 117405 152768 117410 152824
rect 117466 152768 118004 152824
rect 117405 152766 118004 152768
rect 113284 152764 113290 152766
rect 113173 152763 113239 152764
rect 117405 152763 117471 152766
rect 117998 152764 118004 152766
rect 118068 152764 118074 152828
rect 120073 152826 120139 152829
rect 120758 152826 120764 152828
rect 120073 152824 120764 152826
rect 120073 152768 120078 152824
rect 120134 152768 120764 152824
rect 120073 152766 120764 152768
rect 120073 152763 120139 152766
rect 120758 152764 120764 152766
rect 120828 152764 120834 152828
rect 122598 152764 122604 152828
rect 122668 152826 122674 152828
rect 122833 152826 122899 152829
rect 122668 152824 122899 152826
rect 122668 152768 122838 152824
rect 122894 152768 122899 152824
rect 122668 152766 122899 152768
rect 122668 152764 122674 152766
rect 122833 152763 122899 152766
rect 183134 152764 183140 152828
rect 183204 152826 183210 152828
rect 183461 152826 183527 152829
rect 183204 152824 183527 152826
rect 183204 152768 183466 152824
rect 183522 152768 183527 152824
rect 183204 152766 183527 152768
rect 183204 152764 183210 152766
rect 183461 152763 183527 152766
rect 207657 152826 207723 152829
rect 311014 152826 311020 152828
rect 207657 152824 311020 152826
rect 207657 152768 207662 152824
rect 207718 152768 311020 152824
rect 207657 152766 311020 152768
rect 207657 152763 207723 152766
rect 311014 152764 311020 152766
rect 311084 152764 311090 152828
rect 343214 152764 343220 152828
rect 343284 152826 343290 152828
rect 343541 152826 343607 152829
rect 343284 152824 343607 152826
rect 343284 152768 343546 152824
rect 343602 152768 343607 152824
rect 343284 152766 343607 152768
rect 343284 152764 343290 152766
rect 343541 152763 343607 152766
rect 378961 152826 379027 152829
rect 468518 152826 468524 152828
rect 378961 152824 468524 152826
rect 378961 152768 378966 152824
rect 379022 152768 468524 152824
rect 378961 152766 468524 152768
rect 378961 152763 379027 152766
rect 468518 152764 468524 152766
rect 468588 152764 468594 152828
rect 49325 152690 49391 152693
rect 160870 152690 160876 152692
rect 49325 152688 160876 152690
rect 49325 152632 49330 152688
rect 49386 152632 160876 152688
rect 49325 152630 160876 152632
rect 49325 152627 49391 152630
rect 160870 152628 160876 152630
rect 160940 152628 160946 152692
rect 214598 152628 214604 152692
rect 214668 152690 214674 152692
rect 259453 152690 259519 152693
rect 260598 152690 260604 152692
rect 214668 152630 259378 152690
rect 214668 152628 214674 152630
rect 76005 152554 76071 152557
rect 77150 152554 77156 152556
rect 76005 152552 77156 152554
rect 76005 152496 76010 152552
rect 76066 152496 77156 152552
rect 76005 152494 77156 152496
rect 76005 152491 76071 152494
rect 77150 152492 77156 152494
rect 77220 152492 77226 152556
rect 88885 152554 88951 152557
rect 115933 152556 115999 152557
rect 183461 152556 183527 152557
rect 93710 152554 93716 152556
rect 88885 152552 93716 152554
rect 88885 152496 88890 152552
rect 88946 152496 93716 152552
rect 88885 152494 93716 152496
rect 88885 152491 88951 152494
rect 93710 152492 93716 152494
rect 93780 152492 93786 152556
rect 115933 152554 115980 152556
rect 115888 152552 115980 152554
rect 115888 152496 115938 152552
rect 115888 152494 115980 152496
rect 115933 152492 115980 152494
rect 116044 152492 116050 152556
rect 183461 152552 183508 152556
rect 183572 152554 183578 152556
rect 183461 152496 183466 152552
rect 183461 152492 183508 152496
rect 183572 152494 183618 152554
rect 183572 152492 183578 152494
rect 203190 152492 203196 152556
rect 203260 152554 203266 152556
rect 258257 152554 258323 152557
rect 258390 152554 258396 152556
rect 203260 152494 258090 152554
rect 203260 152492 203266 152494
rect 115933 152491 115999 152492
rect 183461 152491 183527 152492
rect 88333 152420 88399 152421
rect 88333 152418 88380 152420
rect 88288 152416 88380 152418
rect 88288 152360 88338 152416
rect 88288 152358 88380 152360
rect 88333 152356 88380 152358
rect 88444 152356 88450 152420
rect 89713 152418 89779 152421
rect 90766 152418 90772 152420
rect 89713 152416 90772 152418
rect 89713 152360 89718 152416
rect 89774 152360 90772 152416
rect 89713 152358 90772 152360
rect 88333 152355 88399 152356
rect 89713 152355 89779 152358
rect 90766 152356 90772 152358
rect 90836 152356 90842 152420
rect 235993 152418 236059 152421
rect 237046 152418 237052 152420
rect 235993 152416 237052 152418
rect 235993 152360 235998 152416
rect 236054 152360 237052 152416
rect 235993 152358 237052 152360
rect 235993 152355 236059 152358
rect 237046 152356 237052 152358
rect 237116 152356 237122 152420
rect 244365 152418 244431 152421
rect 245326 152418 245332 152420
rect 244365 152416 245332 152418
rect 244365 152360 244370 152416
rect 244426 152360 245332 152416
rect 244365 152358 245332 152360
rect 244365 152355 244431 152358
rect 245326 152356 245332 152358
rect 245396 152356 245402 152420
rect 247125 152418 247191 152421
rect 248270 152418 248276 152420
rect 247125 152416 248276 152418
rect 247125 152360 247130 152416
rect 247186 152360 248276 152416
rect 247125 152358 248276 152360
rect 247125 152355 247191 152358
rect 248270 152356 248276 152358
rect 248340 152356 248346 152420
rect 251265 152418 251331 152421
rect 252318 152418 252324 152420
rect 251265 152416 252324 152418
rect 251265 152360 251270 152416
rect 251326 152360 252324 152416
rect 251265 152358 252324 152360
rect 251265 152355 251331 152358
rect 252318 152356 252324 152358
rect 252388 152356 252394 152420
rect 258030 152418 258090 152494
rect 258257 152552 258396 152554
rect 258257 152496 258262 152552
rect 258318 152496 258396 152552
rect 258257 152494 258396 152496
rect 258257 152491 258323 152494
rect 258390 152492 258396 152494
rect 258460 152492 258466 152556
rect 259318 152554 259378 152630
rect 259453 152688 260604 152690
rect 259453 152632 259458 152688
rect 259514 152632 260604 152688
rect 259453 152630 260604 152632
rect 259453 152627 259519 152630
rect 260598 152628 260604 152630
rect 260668 152628 260674 152692
rect 265065 152690 265131 152693
rect 265934 152690 265940 152692
rect 265065 152688 265940 152690
rect 265065 152632 265070 152688
rect 265126 152632 265940 152688
rect 265065 152630 265940 152632
rect 265065 152627 265131 152630
rect 265934 152628 265940 152630
rect 266004 152628 266010 152692
rect 266445 152690 266511 152693
rect 267590 152690 267596 152692
rect 266445 152688 267596 152690
rect 266445 152632 266450 152688
rect 266506 152632 267596 152688
rect 266445 152630 267596 152632
rect 266445 152627 266511 152630
rect 267590 152628 267596 152630
rect 267660 152628 267666 152692
rect 268009 152690 268075 152693
rect 268326 152690 268332 152692
rect 268009 152688 268332 152690
rect 268009 152632 268014 152688
rect 268070 152632 268332 152688
rect 268009 152630 268332 152632
rect 268009 152627 268075 152630
rect 268326 152628 268332 152630
rect 268396 152628 268402 152692
rect 273294 152628 273300 152692
rect 273364 152690 273370 152692
rect 274633 152690 274699 152693
rect 273364 152688 274699 152690
rect 273364 152632 274638 152688
rect 274694 152632 274699 152688
rect 273364 152630 274699 152632
rect 273364 152628 273370 152630
rect 274633 152627 274699 152630
rect 379145 152690 379211 152693
rect 460974 152690 460980 152692
rect 379145 152688 460980 152690
rect 379145 152632 379150 152688
rect 379206 152632 460980 152688
rect 379145 152630 460980 152632
rect 379145 152627 379211 152630
rect 460974 152628 460980 152630
rect 461044 152628 461050 152692
rect 503478 152628 503484 152692
rect 503548 152690 503554 152692
rect 503621 152690 503687 152693
rect 503548 152688 503687 152690
rect 503548 152632 503626 152688
rect 503682 152632 503687 152688
rect 503548 152630 503687 152632
rect 503548 152628 503554 152630
rect 503621 152627 503687 152630
rect 276238 152554 276244 152556
rect 259318 152494 276244 152554
rect 276238 152492 276244 152494
rect 276308 152492 276314 152556
rect 343398 152492 343404 152556
rect 343468 152554 343474 152556
rect 343541 152554 343607 152557
rect 343468 152552 343607 152554
rect 343468 152496 343546 152552
rect 343602 152496 343607 152552
rect 343468 152494 343607 152496
rect 343468 152492 343474 152494
rect 343541 152491 343607 152494
rect 396165 152554 396231 152557
rect 397126 152554 397132 152556
rect 396165 152552 397132 152554
rect 396165 152496 396170 152552
rect 396226 152496 397132 152552
rect 396165 152494 397132 152496
rect 396165 152491 396231 152494
rect 397126 152492 397132 152494
rect 397196 152492 397202 152556
rect 402973 152554 403039 152557
rect 404118 152554 404124 152556
rect 402973 152552 404124 152554
rect 402973 152496 402978 152552
rect 403034 152496 404124 152552
rect 402973 152494 404124 152496
rect 402973 152491 403039 152494
rect 404118 152492 404124 152494
rect 404188 152492 404194 152556
rect 409873 152554 409939 152557
rect 410742 152554 410748 152556
rect 409873 152552 410748 152554
rect 409873 152496 409878 152552
rect 409934 152496 410748 152552
rect 409873 152494 410748 152496
rect 409873 152491 409939 152494
rect 410742 152492 410748 152494
rect 410812 152492 410818 152556
rect 411253 152554 411319 152557
rect 412398 152554 412404 152556
rect 411253 152552 412404 152554
rect 411253 152496 411258 152552
rect 411314 152496 412404 152552
rect 411253 152494 412404 152496
rect 411253 152491 411319 152494
rect 412398 152492 412404 152494
rect 412468 152492 412474 152556
rect 413093 152554 413159 152557
rect 413686 152554 413692 152556
rect 413093 152552 413692 152554
rect 413093 152496 413098 152552
rect 413154 152496 413692 152552
rect 413093 152494 413692 152496
rect 413093 152491 413159 152494
rect 413686 152492 413692 152494
rect 413756 152492 413762 152556
rect 418153 152554 418219 152557
rect 419206 152554 419212 152556
rect 418153 152552 419212 152554
rect 418153 152496 418158 152552
rect 418214 152496 419212 152552
rect 418153 152494 419212 152496
rect 418153 152491 418219 152494
rect 419206 152492 419212 152494
rect 419276 152492 419282 152556
rect 426433 152554 426499 152557
rect 427670 152554 427676 152556
rect 426433 152552 427676 152554
rect 426433 152496 426438 152552
rect 426494 152496 427676 152552
rect 426433 152494 427676 152496
rect 426433 152491 426499 152494
rect 427670 152492 427676 152494
rect 427740 152492 427746 152556
rect 433374 152492 433380 152556
rect 433444 152554 433450 152556
rect 434713 152554 434779 152557
rect 433444 152552 434779 152554
rect 433444 152496 434718 152552
rect 434774 152496 434779 152552
rect 433444 152494 434779 152496
rect 433444 152492 433450 152494
rect 434713 152491 434779 152494
rect 435766 152492 435772 152556
rect 435836 152554 435842 152556
rect 436093 152554 436159 152557
rect 435836 152552 436159 152554
rect 435836 152496 436098 152552
rect 436154 152496 436159 152552
rect 435836 152494 436159 152496
rect 435836 152492 435842 152494
rect 436093 152491 436159 152494
rect 437473 152554 437539 152557
rect 438526 152554 438532 152556
rect 437473 152552 438532 152554
rect 437473 152496 437478 152552
rect 437534 152496 438532 152552
rect 437473 152494 438532 152496
rect 437473 152491 437539 152494
rect 438526 152492 438532 152494
rect 438596 152492 438602 152556
rect 503110 152492 503116 152556
rect 503180 152554 503186 152556
rect 503621 152554 503687 152557
rect 503180 152552 503687 152554
rect 503180 152496 503626 152552
rect 503682 152496 503687 152552
rect 503180 152494 503687 152496
rect 503180 152492 503186 152494
rect 503621 152491 503687 152494
rect 263542 152418 263548 152420
rect 258030 152358 263548 152418
rect 263542 152356 263548 152358
rect 263612 152356 263618 152420
rect 407113 152418 407179 152421
rect 408166 152418 408172 152420
rect 407113 152416 408172 152418
rect 407113 152360 407118 152416
rect 407174 152360 408172 152416
rect 407113 152358 408172 152360
rect 407113 152355 407179 152358
rect 408166 152356 408172 152358
rect 408236 152356 408242 152420
rect 367921 152282 367987 152285
rect 465942 152282 465948 152284
rect 367921 152280 465948 152282
rect 367921 152224 367926 152280
rect 367982 152224 465948 152280
rect 367921 152222 465948 152224
rect 367921 152219 367987 152222
rect 465942 152220 465948 152222
rect 466012 152220 466018 152284
rect 104893 152146 104959 152149
rect 105302 152146 105308 152148
rect 104893 152144 105308 152146
rect 104893 152088 104898 152144
rect 104954 152088 105308 152144
rect 104893 152086 105308 152088
rect 104893 152083 104959 152086
rect 105302 152084 105308 152086
rect 105372 152084 105378 152148
rect 202270 152084 202276 152148
rect 202340 152146 202346 152148
rect 325550 152146 325556 152148
rect 202340 152086 325556 152146
rect 202340 152084 202346 152086
rect 325550 152084 325556 152086
rect 325620 152084 325626 152148
rect 80053 152010 80119 152013
rect 80462 152010 80468 152012
rect 80053 152008 80468 152010
rect 80053 151952 80058 152008
rect 80114 151952 80468 152008
rect 80053 151950 80468 151952
rect 80053 151947 80119 151950
rect 80462 151948 80468 151950
rect 80532 151948 80538 152012
rect 84142 151948 84148 152012
rect 84212 152010 84218 152012
rect 84285 152010 84351 152013
rect 238753 152012 238819 152013
rect 84212 152008 84351 152010
rect 84212 151952 84290 152008
rect 84346 151952 84351 152008
rect 84212 151950 84351 151952
rect 84212 151948 84218 151950
rect 84285 151947 84351 151950
rect 238702 151948 238708 152012
rect 238772 152010 238819 152012
rect 238772 152008 238864 152010
rect 238814 151952 238864 152008
rect 238772 151950 238864 151952
rect 238772 151948 238819 151950
rect 276974 151948 276980 152012
rect 277044 152010 277050 152012
rect 277393 152010 277459 152013
rect 277044 152008 277459 152010
rect 277044 151952 277398 152008
rect 277454 151952 277459 152008
rect 277044 151950 277459 151952
rect 277044 151948 277050 151950
rect 238753 151947 238819 151948
rect 277393 151947 277459 151950
rect 277342 151812 277348 151876
rect 277412 151874 277418 151876
rect 278681 151874 278747 151877
rect 277412 151872 278747 151874
rect 277412 151816 278686 151872
rect 278742 151816 278747 151872
rect 277412 151814 278747 151816
rect 277412 151812 277418 151814
rect 278681 151811 278747 151814
rect 205398 151676 205404 151740
rect 205468 151738 205474 151740
rect 322974 151738 322980 151740
rect 205468 151678 322980 151738
rect 205468 151676 205474 151678
rect 322974 151676 322980 151678
rect 323044 151676 323050 151740
rect 358537 151738 358603 151741
rect 430614 151738 430620 151740
rect 358537 151736 430620 151738
rect 358537 151680 358542 151736
rect 358598 151680 430620 151736
rect 358537 151678 430620 151680
rect 358537 151675 358603 151678
rect 430614 151676 430620 151678
rect 430684 151676 430690 151740
rect 361205 151602 361271 151605
rect 427854 151602 427860 151604
rect 361205 151600 427860 151602
rect 361205 151544 361210 151600
rect 361266 151544 427860 151600
rect 361205 151542 427860 151544
rect 361205 151539 361271 151542
rect 427854 151540 427860 151542
rect 427924 151540 427930 151604
rect 379462 151268 379468 151332
rect 379532 151330 379538 151332
rect 380801 151330 380867 151333
rect 379532 151328 380867 151330
rect 379532 151272 380806 151328
rect 380862 151272 380867 151328
rect 379532 151270 380867 151272
rect 379532 151268 379538 151270
rect 380801 151267 380867 151270
rect 57789 150516 57855 150517
rect 57789 150512 57836 150516
rect 57900 150514 57906 150516
rect 57789 150456 57794 150512
rect 57789 150452 57836 150456
rect 57900 150454 57946 150514
rect 57900 150452 57906 150454
rect 57789 150451 57855 150452
rect 580901 147250 580967 147253
rect 583520 147250 584960 147340
rect 580901 147248 584960 147250
rect 580901 147192 580906 147248
rect 580962 147192 584960 147248
rect 580901 147190 584960 147192
rect 580901 147187 580967 147190
rect 583520 147100 584960 147190
rect -960 144380 480 144620
rect 583520 134316 584960 134556
rect 56961 133786 57027 133789
rect 57094 133786 57100 133788
rect 56961 133784 57100 133786
rect 56961 133728 56966 133784
rect 57022 133728 57100 133784
rect 56961 133726 57100 133728
rect 56961 133723 57027 133726
rect 57094 133724 57100 133726
rect 57164 133724 57170 133788
rect 374361 133786 374427 133789
rect 377254 133786 377260 133788
rect 374361 133784 377260 133786
rect 374361 133728 374366 133784
rect 374422 133728 377260 133784
rect 374361 133726 377260 133728
rect 374361 133723 374427 133726
rect 377254 133724 377260 133726
rect 377324 133786 377330 133788
rect 377673 133786 377739 133789
rect 377324 133784 377739 133786
rect 377324 133728 377678 133784
rect 377734 133728 377739 133784
rect 377324 133726 377739 133728
rect 377324 133724 377330 133726
rect 377673 133723 377739 133726
rect 98637 133106 98703 133109
rect 56550 133104 98703 133106
rect 56550 133048 98642 133104
rect 98698 133048 98703 133104
rect 56550 133046 98703 133048
rect 51625 132426 51691 132429
rect 56550 132426 56610 133046
rect 98637 133043 98703 133046
rect 377806 133044 377812 133108
rect 377876 133106 377882 133108
rect 438853 133106 438919 133109
rect 377876 133104 438919 133106
rect 377876 133048 438858 133104
rect 438914 133048 438919 133104
rect 377876 133046 438919 133048
rect 377876 133044 377882 133046
rect 438853 133043 438919 133046
rect 57094 132426 57100 132428
rect 51625 132424 57100 132426
rect 51625 132368 51630 132424
rect 51686 132368 57100 132424
rect 51625 132366 57100 132368
rect 51625 132363 51691 132366
rect 57094 132364 57100 132366
rect 57164 132364 57170 132428
rect -960 131868 480 132108
rect 56041 131066 56107 131069
rect 57973 131066 58039 131069
rect 102133 131066 102199 131069
rect 56041 131064 102199 131066
rect 56041 131008 56046 131064
rect 56102 131008 57978 131064
rect 58034 131008 102138 131064
rect 102194 131008 102199 131064
rect 56041 131006 102199 131008
rect 56041 131003 56107 131006
rect 57973 131003 58039 131006
rect 102133 131003 102199 131006
rect 214373 131066 214439 131069
rect 274633 131066 274699 131069
rect 214373 131064 274699 131066
rect 214373 131008 214378 131064
rect 214434 131008 274638 131064
rect 274694 131008 274699 131064
rect 214373 131006 274699 131008
rect 214373 131003 214439 131006
rect 274633 131003 274699 131006
rect 379605 131066 379671 131069
rect 426433 131066 426499 131069
rect 379605 131064 426499 131066
rect 379605 131008 379610 131064
rect 379666 131008 426438 131064
rect 426494 131008 426499 131064
rect 379605 131006 426499 131008
rect 379605 131003 379671 131006
rect 426433 131003 426499 131006
rect 53005 130930 53071 130933
rect 56133 130930 56199 130933
rect 53005 130928 56199 130930
rect 53005 130872 53010 130928
rect 53066 130872 56138 130928
rect 56194 130872 56199 130928
rect 53005 130870 56199 130872
rect 53005 130867 53071 130870
rect 56133 130867 56199 130870
rect 217542 130868 217548 130932
rect 217612 130930 217618 130932
rect 249793 130930 249859 130933
rect 217612 130928 249859 130930
rect 217612 130872 249798 130928
rect 249854 130872 249859 130928
rect 217612 130870 249859 130872
rect 217612 130868 217618 130870
rect 249793 130867 249859 130870
rect 377990 130868 377996 130932
rect 378060 130930 378066 130932
rect 416773 130930 416839 130933
rect 378060 130928 416839 130930
rect 378060 130872 416778 130928
rect 416834 130872 416839 130928
rect 378060 130870 416839 130872
rect 378060 130868 378066 130870
rect 416773 130867 416839 130870
rect 379881 130794 379947 130797
rect 414013 130794 414079 130797
rect 379881 130792 414079 130794
rect 379881 130736 379886 130792
rect 379942 130736 414018 130792
rect 414074 130736 414079 130792
rect 379881 130734 414079 130736
rect 379881 130731 379947 130734
rect 414013 130731 414079 130734
rect 50429 130658 50495 130661
rect 58985 130658 59051 130661
rect 97257 130658 97323 130661
rect 50429 130656 97323 130658
rect 50429 130600 50434 130656
rect 50490 130600 58990 130656
rect 59046 130600 97262 130656
rect 97318 130600 97323 130656
rect 50429 130598 97323 130600
rect 50429 130595 50495 130598
rect 58985 130595 59051 130598
rect 97257 130595 97323 130598
rect 56133 130522 56199 130525
rect 95233 130522 95299 130525
rect 56133 130520 95299 130522
rect 56133 130464 56138 130520
rect 56194 130464 95238 130520
rect 95294 130464 95299 130520
rect 56133 130462 95299 130464
rect 56133 130459 56199 130462
rect 95233 130459 95299 130462
rect 210877 130522 210943 130525
rect 214833 130522 214899 130525
rect 237373 130522 237439 130525
rect 210877 130520 237439 130522
rect 210877 130464 210882 130520
rect 210938 130464 214838 130520
rect 214894 130464 237378 130520
rect 237434 130464 237439 130520
rect 210877 130462 237439 130464
rect 210877 130459 210943 130462
rect 214833 130459 214899 130462
rect 237373 130459 237439 130462
rect 57278 130324 57284 130388
rect 57348 130386 57354 130388
rect 99373 130386 99439 130389
rect 57348 130384 99439 130386
rect 57348 130328 99378 130384
rect 99434 130328 99439 130384
rect 57348 130326 99439 130328
rect 57348 130324 57354 130326
rect 99373 130323 99439 130326
rect 190862 130324 190868 130388
rect 190932 130386 190938 130388
rect 191741 130386 191807 130389
rect 190932 130384 191807 130386
rect 190932 130328 191746 130384
rect 191802 130328 191807 130384
rect 190932 130326 191807 130328
rect 190932 130324 190938 130326
rect 191741 130323 191807 130326
rect 215845 130386 215911 130389
rect 269113 130386 269179 130389
rect 215845 130384 269179 130386
rect 215845 130328 215850 130384
rect 215906 130328 269118 130384
rect 269174 130328 269179 130384
rect 215845 130326 269179 130328
rect 215845 130323 215911 130326
rect 269113 130323 269179 130326
rect 376569 130386 376635 130389
rect 429193 130386 429259 130389
rect 376569 130384 429259 130386
rect 376569 130328 376574 130384
rect 376630 130328 429198 130384
rect 429254 130328 429259 130384
rect 376569 130326 429259 130328
rect 376569 130323 376635 130326
rect 429193 130323 429259 130326
rect 510613 130386 510679 130389
rect 510838 130386 510844 130388
rect 510613 130384 510844 130386
rect 510613 130328 510618 130384
rect 510674 130328 510844 130384
rect 510613 130326 510844 130328
rect 510613 130323 510679 130326
rect 510838 130324 510844 130326
rect 510908 130324 510914 130388
rect 178534 129780 178540 129844
rect 178604 129842 178610 129844
rect 179045 129842 179111 129845
rect 178604 129840 179111 129842
rect 178604 129784 179050 129840
rect 179106 129784 179111 129840
rect 178604 129782 179111 129784
rect 178604 129780 178610 129782
rect 179045 129779 179111 129782
rect 179638 129780 179644 129844
rect 179708 129842 179714 129844
rect 179781 129842 179847 129845
rect 338481 129844 338547 129845
rect 338430 129842 338436 129844
rect 179708 129840 179847 129842
rect 179708 129784 179786 129840
rect 179842 129784 179847 129840
rect 179708 129782 179847 129784
rect 338390 129782 338436 129842
rect 338500 129840 338547 129844
rect 338542 129784 338547 129840
rect 179708 129780 179714 129782
rect 179781 129779 179847 129782
rect 338430 129780 338436 129782
rect 338500 129780 338547 129784
rect 339718 129780 339724 129844
rect 339788 129842 339794 129844
rect 340597 129842 340663 129845
rect 339788 129840 340663 129842
rect 339788 129784 340602 129840
rect 340658 129784 340663 129840
rect 339788 129782 340663 129784
rect 339788 129780 339794 129782
rect 338481 129779 338547 129780
rect 340597 129779 340663 129782
rect 350942 129780 350948 129844
rect 351012 129842 351018 129844
rect 351729 129842 351795 129845
rect 351012 129840 351795 129842
rect 351012 129784 351734 129840
rect 351790 129784 351795 129840
rect 351012 129782 351795 129784
rect 351012 129780 351018 129782
rect 351729 129779 351795 129782
rect 377213 129842 377279 129845
rect 377990 129842 377996 129844
rect 377213 129840 377996 129842
rect 377213 129784 377218 129840
rect 377274 129784 377996 129840
rect 377213 129782 377996 129784
rect 377213 129779 377279 129782
rect 377990 129780 377996 129782
rect 378060 129780 378066 129844
rect 498510 129780 498516 129844
rect 498580 129842 498586 129844
rect 498745 129842 498811 129845
rect 498580 129840 498811 129842
rect 498580 129784 498750 129840
rect 498806 129784 498811 129840
rect 498580 129782 498811 129784
rect 498580 129780 498586 129782
rect 498745 129779 498811 129782
rect 499798 129780 499804 129844
rect 499868 129842 499874 129844
rect 500217 129842 500283 129845
rect 499868 129840 500283 129842
rect 499868 129784 500222 129840
rect 500278 129784 500283 129840
rect 499868 129782 500283 129784
rect 499868 129780 499874 129782
rect 500217 129779 500283 129782
rect 54385 129706 54451 129709
rect 54702 129706 54708 129708
rect 54385 129704 54708 129706
rect 54385 129648 54390 129704
rect 54446 129648 54708 129704
rect 54385 129646 54708 129648
rect 54385 129643 54451 129646
rect 54702 129644 54708 129646
rect 54772 129644 54778 129708
rect 54293 129570 54359 129573
rect 57278 129570 57284 129572
rect 54293 129568 57284 129570
rect 54293 129512 54298 129568
rect 54354 129512 57284 129568
rect 54293 129510 57284 129512
rect 54293 129507 54359 129510
rect 57278 129508 57284 129510
rect 57348 129508 57354 129572
rect 196604 124160 197186 124220
rect 197126 124130 197186 124160
rect 199193 124130 199259 124133
rect 197126 124128 199259 124130
rect 197126 124072 199198 124128
rect 199254 124072 199259 124128
rect 197126 124070 199259 124072
rect 356562 124130 356622 124190
rect 516588 124160 517162 124220
rect 359273 124130 359339 124133
rect 356562 124128 359339 124130
rect 356562 124072 359278 124128
rect 359334 124072 359339 124128
rect 356562 124070 359339 124072
rect 517102 124130 517162 124160
rect 519353 124130 519419 124133
rect 517102 124128 519419 124130
rect 517102 124072 519358 124128
rect 519414 124072 519419 124128
rect 517102 124070 519419 124072
rect 199193 124067 199259 124070
rect 359273 124067 359339 124070
rect 519353 124067 519419 124070
rect 583520 121396 584960 121636
rect -960 119370 480 119460
rect 2957 119370 3023 119373
rect -960 119368 3023 119370
rect -960 119312 2962 119368
rect 3018 119312 3023 119368
rect -960 119310 3023 119312
rect -960 119220 480 119310
rect 2957 119307 3023 119310
rect 580901 108762 580967 108765
rect 583520 108762 584960 108852
rect 580901 108760 584960 108762
rect 580901 108704 580906 108760
rect 580962 108704 584960 108760
rect 580901 108702 584960 108704
rect 580901 108699 580967 108702
rect 583520 108612 584960 108702
rect -960 106858 480 106948
rect 2773 106858 2839 106861
rect -960 106856 2839 106858
rect -960 106800 2778 106856
rect 2834 106800 2839 106856
rect -960 106798 2839 106800
rect -960 106708 480 106798
rect 2773 106795 2839 106798
rect 583520 95828 584960 96068
rect -960 94196 480 94436
rect 583520 83044 584960 83284
rect 57605 82514 57671 82517
rect 57605 82512 60062 82514
rect 57605 82456 57610 82512
rect 57666 82456 60062 82512
rect 57605 82454 60062 82456
rect 57605 82451 57671 82454
rect 60002 81894 60062 82454
rect 216765 81970 216831 81973
rect 377949 81970 378015 81973
rect 216765 81968 219450 81970
rect 216765 81912 216770 81968
rect 216826 81924 219450 81968
rect 377949 81968 379530 81970
rect 216826 81912 220064 81924
rect 216765 81910 220064 81912
rect 216765 81907 216831 81910
rect 219390 81864 220064 81910
rect 377949 81912 377954 81968
rect 378010 81924 379530 81968
rect 378010 81912 380052 81924
rect 377949 81910 380052 81912
rect 377949 81907 378015 81910
rect 379470 81864 380052 81910
rect -960 81698 480 81788
rect 3417 81698 3483 81701
rect -960 81696 3483 81698
rect -960 81640 3422 81696
rect 3478 81640 3483 81696
rect -960 81638 3483 81640
rect -960 81548 480 81638
rect 3417 81635 3483 81638
rect 56777 81426 56843 81429
rect 56777 81424 60062 81426
rect 56777 81368 56782 81424
rect 56838 81368 60062 81424
rect 56777 81366 60062 81368
rect 56777 81363 56843 81366
rect 60002 80942 60062 81366
rect 216857 81018 216923 81021
rect 377857 81018 377923 81021
rect 216857 81016 219450 81018
rect 216857 80960 216862 81016
rect 216918 80972 219450 81016
rect 377857 81016 379530 81018
rect 216918 80960 220064 80972
rect 216857 80958 220064 80960
rect 216857 80955 216923 80958
rect 219390 80912 220064 80958
rect 377857 80960 377862 81016
rect 377918 80972 379530 81016
rect 377918 80960 380052 80972
rect 377857 80958 380052 80960
rect 377857 80955 377923 80958
rect 379470 80912 380052 80958
rect 57329 79386 57395 79389
rect 57329 79384 60062 79386
rect 57329 79328 57334 79384
rect 57390 79328 60062 79384
rect 57329 79326 60062 79328
rect 57329 79323 57395 79326
rect 60002 78766 60062 79326
rect 217777 78842 217843 78845
rect 377305 78842 377371 78845
rect 217777 78840 219450 78842
rect 217777 78784 217782 78840
rect 217838 78796 219450 78840
rect 377305 78840 379530 78842
rect 217838 78784 220064 78796
rect 217777 78782 220064 78784
rect 217777 78779 217843 78782
rect 219390 78736 220064 78782
rect 377305 78784 377310 78840
rect 377366 78796 379530 78840
rect 377366 78784 380052 78796
rect 377305 78782 380052 78784
rect 377305 78779 377371 78782
rect 379470 78736 380052 78782
rect 56869 78434 56935 78437
rect 56869 78432 60062 78434
rect 56869 78376 56874 78432
rect 56930 78376 60062 78432
rect 56869 78374 60062 78376
rect 56869 78371 56935 78374
rect 60002 77814 60062 78374
rect 217961 77890 218027 77893
rect 378041 77890 378107 77893
rect 217961 77888 219450 77890
rect 217961 77832 217966 77888
rect 218022 77844 219450 77888
rect 378041 77888 379530 77890
rect 218022 77832 220064 77844
rect 217961 77830 220064 77832
rect 217961 77827 218027 77830
rect 219390 77784 220064 77830
rect 378041 77832 378046 77888
rect 378102 77844 379530 77888
rect 378102 77832 380052 77844
rect 378041 77830 380052 77832
rect 378041 77827 378107 77830
rect 379470 77784 380052 77830
rect 57145 76666 57211 76669
rect 57145 76664 60062 76666
rect 57145 76608 57150 76664
rect 57206 76608 60062 76664
rect 57145 76606 60062 76608
rect 57145 76603 57211 76606
rect 60002 76046 60062 76606
rect 217501 76122 217567 76125
rect 376937 76122 377003 76125
rect 217501 76120 219450 76122
rect 217501 76064 217506 76120
rect 217562 76076 219450 76120
rect 376937 76120 379530 76122
rect 217562 76064 220064 76076
rect 217501 76062 220064 76064
rect 217501 76059 217567 76062
rect 219390 76016 220064 76062
rect 376937 76064 376942 76120
rect 376998 76076 379530 76120
rect 376998 76064 380052 76076
rect 376937 76062 380052 76064
rect 376937 76059 377003 76062
rect 379470 76016 380052 76062
rect 57697 75578 57763 75581
rect 57697 75576 60062 75578
rect 57697 75520 57702 75576
rect 57758 75520 60062 75576
rect 57697 75518 60062 75520
rect 57697 75515 57763 75518
rect 60002 74958 60062 75518
rect 216949 75034 217015 75037
rect 377121 75034 377187 75037
rect 216949 75032 219450 75034
rect 216949 74976 216954 75032
rect 217010 74988 219450 75032
rect 377121 75032 379530 75034
rect 217010 74976 220064 74988
rect 216949 74974 220064 74976
rect 216949 74971 217015 74974
rect 219390 74928 220064 74974
rect 377121 74976 377126 75032
rect 377182 74988 379530 75032
rect 377182 74976 380052 74988
rect 377121 74974 380052 74976
rect 377121 74971 377187 74974
rect 379470 74928 380052 74974
rect 57421 73810 57487 73813
rect 57421 73808 60062 73810
rect 57421 73752 57426 73808
rect 57482 73752 60062 73808
rect 57421 73750 60062 73752
rect 57421 73747 57487 73750
rect 60002 73190 60062 73750
rect 217409 73266 217475 73269
rect 377489 73266 377555 73269
rect 217409 73264 219450 73266
rect 217409 73208 217414 73264
rect 217470 73220 219450 73264
rect 377489 73264 379530 73266
rect 217470 73208 220064 73220
rect 217409 73206 220064 73208
rect 217409 73203 217475 73206
rect 219390 73160 220064 73206
rect 377489 73208 377494 73264
rect 377550 73220 379530 73264
rect 377550 73208 380052 73220
rect 377489 73206 380052 73208
rect 377489 73203 377555 73206
rect 379470 73160 380052 73206
rect 580901 70410 580967 70413
rect 583520 70410 584960 70500
rect 580901 70408 584960 70410
rect 580901 70352 580906 70408
rect 580962 70352 584960 70408
rect 580901 70350 584960 70352
rect 580901 70347 580967 70350
rect 583520 70260 584960 70350
rect -960 69186 480 69276
rect 2773 69186 2839 69189
rect -960 69184 2839 69186
rect -960 69128 2778 69184
rect 2834 69128 2839 69184
rect -960 69126 2839 69128
rect -960 69036 480 69126
rect 2773 69123 2839 69126
rect 518893 64834 518959 64837
rect 516558 64832 518959 64834
rect 516558 64776 518898 64832
rect 518954 64776 518959 64832
rect 516558 64774 518959 64776
rect 199377 64698 199443 64701
rect 359549 64698 359615 64701
rect 196558 64696 199443 64698
rect 196558 64640 199382 64696
rect 199438 64640 199443 64696
rect 196558 64638 199443 64640
rect 196558 64350 196618 64638
rect 199377 64635 199443 64638
rect 356562 64696 359615 64698
rect 356562 64640 359554 64696
rect 359610 64640 359615 64696
rect 356562 64638 359615 64640
rect 356562 64350 356622 64638
rect 359549 64635 359615 64638
rect 516558 64350 516618 64774
rect 518893 64771 518959 64774
rect 199285 63338 199351 63341
rect 359181 63338 359247 63341
rect 519445 63338 519511 63341
rect 196558 63336 199351 63338
rect 196558 63280 199290 63336
rect 199346 63280 199351 63336
rect 196558 63278 199351 63280
rect 196558 62718 196618 63278
rect 199285 63275 199351 63278
rect 356562 63336 359247 63338
rect 356562 63280 359186 63336
rect 359242 63280 359247 63336
rect 356562 63278 359247 63280
rect 356562 62718 356622 63278
rect 359181 63275 359247 63278
rect 516558 63336 519511 63338
rect 516558 63280 519450 63336
rect 519506 63280 519511 63336
rect 516558 63278 519511 63280
rect 516558 62718 516618 63278
rect 519445 63275 519511 63278
rect 199101 61978 199167 61981
rect 358813 61978 358879 61981
rect 518985 61978 519051 61981
rect 196558 61976 199167 61978
rect 196558 61920 199106 61976
rect 199162 61920 199167 61976
rect 196558 61918 199167 61920
rect 196558 61358 196618 61918
rect 199101 61915 199167 61918
rect 356562 61976 358879 61978
rect 356562 61920 358818 61976
rect 358874 61920 358879 61976
rect 356562 61918 358879 61920
rect 356562 61358 356622 61918
rect 358813 61915 358879 61918
rect 516558 61976 519051 61978
rect 516558 61920 518990 61976
rect 519046 61920 519051 61976
rect 516558 61918 519051 61920
rect 516558 61358 516618 61918
rect 518985 61915 519051 61918
rect 198825 60482 198891 60485
rect 358905 60482 358971 60485
rect 519077 60482 519143 60485
rect 196558 60480 198891 60482
rect 196558 60424 198830 60480
rect 198886 60424 198891 60480
rect 196558 60422 198891 60424
rect 196558 59862 196618 60422
rect 198825 60419 198891 60422
rect 356562 60480 358971 60482
rect 356562 60424 358910 60480
rect 358966 60424 358971 60480
rect 356562 60422 358971 60424
rect 356562 59862 356622 60422
rect 358905 60419 358971 60422
rect 516558 60480 519143 60482
rect 516558 60424 519082 60480
rect 519138 60424 519143 60480
rect 516558 60422 519143 60424
rect 516558 59862 516618 60422
rect 519077 60419 519143 60422
rect 198733 59258 198799 59261
rect 358997 59258 359063 59261
rect 519261 59258 519327 59261
rect 196558 59256 198799 59258
rect 196558 59200 198738 59256
rect 198794 59200 198799 59256
rect 196558 59198 198799 59200
rect 196558 58638 196618 59198
rect 198733 59195 198799 59198
rect 356562 59256 359063 59258
rect 356562 59200 359002 59256
rect 359058 59200 359063 59256
rect 356562 59198 359063 59200
rect 356562 58638 356622 59198
rect 358997 59195 359063 59198
rect 516558 59256 519327 59258
rect 516558 59200 519266 59256
rect 519322 59200 519327 59256
rect 516558 59198 519327 59200
rect 516558 58638 516618 59198
rect 519261 59195 519327 59198
rect 583520 57476 584960 57716
rect -960 56388 480 56628
rect 202086 54980 202092 55044
rect 202156 55042 202162 55044
rect 376937 55042 377003 55045
rect 202156 54996 219450 55042
rect 376937 55040 379530 55042
rect 202156 54982 220064 54996
rect 202156 54980 202162 54982
rect 46606 53892 46612 53956
rect 46676 53954 46682 53956
rect 60002 53954 60062 54966
rect 219390 54936 220064 54982
rect 376937 54984 376942 55040
rect 376998 54996 379530 55040
rect 376998 54984 380052 54996
rect 376937 54982 380052 54984
rect 376937 54979 377003 54982
rect 379470 54936 380052 54982
rect 46676 53894 60062 53954
rect 46676 53892 46682 53894
rect 57881 53410 57947 53413
rect 57881 53408 60062 53410
rect 57881 53352 57886 53408
rect 57942 53352 60062 53408
rect 57881 53350 60062 53352
rect 57881 53347 57947 53350
rect 60002 53334 60062 53350
rect 219390 53304 220064 53364
rect 379470 53304 380052 53364
rect 216673 53274 216739 53277
rect 219390 53274 219450 53304
rect 216673 53272 219450 53274
rect 216673 53216 216678 53272
rect 216734 53216 219450 53272
rect 216673 53214 219450 53216
rect 376937 53274 377003 53277
rect 379470 53274 379530 53304
rect 376937 53272 379530 53274
rect 376937 53216 376942 53272
rect 376998 53216 379530 53272
rect 376937 53214 379530 53216
rect 216673 53211 216739 53214
rect 376937 53211 377003 53214
rect 206318 53076 206324 53140
rect 206388 53138 206394 53140
rect 376017 53138 376083 53141
rect 206388 53092 219450 53138
rect 376017 53136 379530 53138
rect 206388 53078 220064 53092
rect 206388 53076 206394 53078
rect 46790 52668 46796 52732
rect 46860 52730 46866 52732
rect 60002 52730 60062 53062
rect 219390 53032 220064 53078
rect 376017 53080 376022 53136
rect 376078 53092 379530 53136
rect 376078 53080 380052 53092
rect 376017 53078 380052 53080
rect 376017 53075 376083 53078
rect 379470 53032 380052 53078
rect 46860 52670 60062 52730
rect 46860 52668 46866 52670
rect 77109 44844 77175 44845
rect 83089 44844 83155 44845
rect 84193 44844 84259 44845
rect 94497 44844 94563 44845
rect 96981 44844 97047 44845
rect 98085 44844 98151 44845
rect 77109 44840 77142 44844
rect 77206 44842 77212 44844
rect 77109 44784 77114 44840
rect 77109 44780 77142 44784
rect 77206 44782 77266 44842
rect 83089 44840 83126 44844
rect 83190 44842 83196 44844
rect 83089 44784 83094 44840
rect 77206 44780 77212 44782
rect 83089 44780 83126 44784
rect 83190 44782 83246 44842
rect 84193 44840 84214 44844
rect 84278 44842 84284 44844
rect 84193 44784 84198 44840
rect 83190 44780 83196 44782
rect 84193 44780 84214 44784
rect 84278 44782 84350 44842
rect 94497 44840 94550 44844
rect 94614 44842 94620 44844
rect 94497 44784 94502 44840
rect 84278 44780 84284 44782
rect 94497 44780 94550 44784
rect 94614 44782 94654 44842
rect 96981 44840 96998 44844
rect 97062 44842 97068 44844
rect 98080 44842 98086 44844
rect 96981 44784 96986 44840
rect 94614 44780 94620 44782
rect 96981 44780 96998 44784
rect 97062 44782 97138 44842
rect 97994 44782 98086 44842
rect 97062 44780 97068 44782
rect 98080 44780 98086 44782
rect 98150 44780 98156 44844
rect 218830 44780 218836 44844
rect 218900 44842 218906 44844
rect 218973 44842 219039 44845
rect 219249 44844 219315 44845
rect 219198 44842 219204 44844
rect 218900 44840 219039 44842
rect 218900 44784 218978 44840
rect 219034 44784 219039 44840
rect 218900 44782 219039 44784
rect 219158 44782 219204 44842
rect 219268 44840 219315 44844
rect 219310 44784 219315 44840
rect 218900 44780 218906 44782
rect 77109 44779 77175 44780
rect 83089 44779 83155 44780
rect 84193 44779 84259 44780
rect 94497 44779 94563 44780
rect 96981 44779 97047 44780
rect 98085 44779 98151 44780
rect 218973 44779 219039 44782
rect 219198 44780 219204 44782
rect 219268 44780 219315 44784
rect 219249 44779 219315 44780
rect 235993 44844 236059 44845
rect 237097 44844 237163 44845
rect 243077 44844 243143 44845
rect 244273 44844 244339 44845
rect 396073 44844 396139 44845
rect 235993 44840 236054 44844
rect 235993 44784 235998 44840
rect 235993 44780 236054 44784
rect 236118 44842 236124 44844
rect 236118 44782 236150 44842
rect 237097 44840 237142 44844
rect 237206 44842 237212 44844
rect 237097 44784 237102 44840
rect 236118 44780 236124 44782
rect 237097 44780 237142 44784
rect 237206 44782 237254 44842
rect 243077 44840 243126 44844
rect 243190 44842 243196 44844
rect 244208 44842 244214 44844
rect 243077 44784 243082 44840
rect 237206 44780 237212 44782
rect 243077 44780 243126 44784
rect 243190 44782 243234 44842
rect 244182 44782 244214 44842
rect 243190 44780 243196 44782
rect 244208 44780 244214 44782
rect 244278 44840 244339 44844
rect 396048 44842 396054 44844
rect 244334 44784 244339 44840
rect 244278 44780 244339 44784
rect 395982 44782 396054 44842
rect 396118 44840 396139 44844
rect 396134 44784 396139 44840
rect 396048 44780 396054 44782
rect 396118 44780 396139 44784
rect 235993 44779 236059 44780
rect 237097 44779 237163 44780
rect 243077 44779 243143 44780
rect 244273 44779 244339 44780
rect 396073 44779 396139 44780
rect 397085 44844 397151 44845
rect 403065 44844 403131 44845
rect 414565 44844 414631 44845
rect 397085 44840 397142 44844
rect 397206 44842 397212 44844
rect 397085 44784 397090 44840
rect 397085 44780 397142 44784
rect 397206 44782 397242 44842
rect 403065 44840 403126 44844
rect 403065 44784 403070 44840
rect 397206 44780 397212 44782
rect 403065 44780 403126 44784
rect 403190 44842 403196 44844
rect 414544 44842 414550 44844
rect 403190 44782 403222 44842
rect 414474 44782 414550 44842
rect 414614 44840 414631 44844
rect 414626 44784 414631 44840
rect 403190 44780 403196 44782
rect 414544 44780 414550 44782
rect 414614 44780 414631 44784
rect 397085 44779 397151 44780
rect 403065 44779 403131 44780
rect 414565 44779 414631 44780
rect 416957 44844 417023 44845
rect 416957 44840 416998 44844
rect 417062 44842 417068 44844
rect 416957 44784 416962 44840
rect 416957 44780 416998 44784
rect 417062 44782 417114 44842
rect 417062 44780 417068 44782
rect 416957 44779 417023 44780
rect 100753 44708 100819 44709
rect 101765 44708 101831 44709
rect 57278 44644 57284 44708
rect 57348 44706 57354 44708
rect 99440 44706 99446 44708
rect 57348 44646 99446 44706
rect 57348 44644 57354 44646
rect 99440 44644 99446 44646
rect 99510 44644 99516 44708
rect 100702 44706 100708 44708
rect 100662 44646 100708 44706
rect 100772 44704 100819 44708
rect 101752 44706 101758 44708
rect 100814 44648 100819 44704
rect 100702 44644 100708 44646
rect 100772 44644 100819 44648
rect 101674 44646 101758 44706
rect 101822 44704 101831 44708
rect 101826 44648 101831 44704
rect 101752 44644 101758 44646
rect 101822 44644 101831 44648
rect 100753 44643 100819 44644
rect 101765 44643 101831 44644
rect 102777 44708 102843 44709
rect 103881 44708 103947 44709
rect 143533 44708 143599 44709
rect 102777 44704 102846 44708
rect 102777 44648 102782 44704
rect 102838 44648 102846 44704
rect 102777 44644 102846 44648
rect 102910 44706 102916 44708
rect 102910 44646 102934 44706
rect 103881 44704 103934 44708
rect 103998 44706 104004 44708
rect 143504 44706 143510 44708
rect 103881 44648 103886 44704
rect 102910 44644 102916 44646
rect 103881 44644 103934 44648
rect 103998 44646 104038 44706
rect 143442 44646 143510 44706
rect 143574 44704 143599 44708
rect 143594 44648 143599 44704
rect 103998 44644 104004 44646
rect 143504 44644 143510 44646
rect 143574 44644 143599 44648
rect 102777 44643 102843 44644
rect 103881 44643 103947 44644
rect 143533 44643 143599 44644
rect 145925 44708 145991 44709
rect 255865 44708 255931 44709
rect 256969 44708 257035 44709
rect 258073 44708 258139 44709
rect 262857 44708 262923 44709
rect 145925 44704 145958 44708
rect 146022 44706 146028 44708
rect 145925 44648 145930 44704
rect 145925 44644 145958 44648
rect 146022 44646 146082 44706
rect 146022 44644 146028 44646
rect 205030 44644 205036 44708
rect 205100 44706 205106 44708
rect 250736 44706 250742 44708
rect 205100 44646 250742 44706
rect 205100 44644 205106 44646
rect 250736 44644 250742 44646
rect 250806 44644 250812 44708
rect 255865 44704 255910 44708
rect 255974 44706 255980 44708
rect 255865 44648 255870 44704
rect 255865 44644 255910 44648
rect 255974 44646 256022 44706
rect 256969 44704 256998 44708
rect 257062 44706 257068 44708
rect 256969 44648 256974 44704
rect 255974 44644 255980 44646
rect 256969 44644 256998 44648
rect 257062 44646 257126 44706
rect 258073 44704 258086 44708
rect 258150 44706 258156 44708
rect 262840 44706 262846 44708
rect 258073 44648 258078 44704
rect 257062 44644 257068 44646
rect 258073 44644 258086 44648
rect 258150 44646 258230 44706
rect 262766 44646 262846 44706
rect 262910 44704 262923 44708
rect 262918 44648 262923 44704
rect 258150 44644 258156 44646
rect 262840 44644 262846 44646
rect 262910 44644 262923 44648
rect 145925 44643 145991 44644
rect 255865 44643 255931 44644
rect 256969 44643 257035 44644
rect 258073 44643 258139 44644
rect 262857 44643 262923 44644
rect 315849 44708 315915 44709
rect 410701 44708 410767 44709
rect 419441 44708 419507 44709
rect 423949 44708 424015 44709
rect 315849 44704 315886 44708
rect 315950 44706 315956 44708
rect 315849 44648 315854 44704
rect 315849 44644 315886 44648
rect 315950 44646 316006 44706
rect 410701 44704 410742 44708
rect 410806 44706 410812 44708
rect 410701 44648 410706 44704
rect 315950 44644 315956 44646
rect 410701 44644 410742 44648
rect 410806 44646 410858 44706
rect 410806 44644 410812 44646
rect 419440 44644 419446 44708
rect 419510 44706 419516 44708
rect 423928 44706 423934 44708
rect 419510 44646 419598 44706
rect 423858 44646 423934 44706
rect 423998 44704 424015 44708
rect 424010 44648 424015 44704
rect 583520 44692 584960 44932
rect 419510 44644 419516 44646
rect 423928 44644 423934 44646
rect 423998 44644 424015 44648
rect 315849 44643 315915 44644
rect 410701 44643 410767 44644
rect 419441 44643 419507 44644
rect 423949 44643 424015 44644
rect 113265 44572 113331 44573
rect 259453 44572 259519 44573
rect 50470 44508 50476 44572
rect 50540 44570 50546 44572
rect 108280 44570 108286 44572
rect 50540 44510 108286 44570
rect 50540 44508 50546 44510
rect 108280 44508 108286 44510
rect 108350 44508 108356 44572
rect 113265 44568 113318 44572
rect 113382 44570 113388 44572
rect 113265 44512 113270 44568
rect 113265 44508 113318 44512
rect 113382 44510 113422 44570
rect 113382 44508 113388 44510
rect 140920 44508 140926 44572
rect 140990 44508 140996 44572
rect 205214 44508 205220 44572
rect 205284 44570 205290 44572
rect 258488 44570 258494 44572
rect 205284 44510 258494 44570
rect 205284 44508 205290 44510
rect 258488 44508 258494 44510
rect 258558 44508 258564 44572
rect 259440 44570 259446 44572
rect 259362 44510 259446 44570
rect 259510 44568 259519 44572
rect 259514 44512 259519 44568
rect 259440 44508 259446 44510
rect 259510 44508 259519 44512
rect 113265 44507 113331 44508
rect 55622 44372 55628 44436
rect 55692 44434 55698 44436
rect 138422 44434 138428 44436
rect 55692 44374 138428 44434
rect 55692 44372 55698 44374
rect 138422 44372 138428 44374
rect 138492 44372 138498 44436
rect 140928 44434 140988 44508
rect 259453 44507 259519 44508
rect 260649 44572 260715 44573
rect 261753 44572 261819 44573
rect 263869 44572 263935 44573
rect 308489 44572 308555 44573
rect 404169 44572 404235 44573
rect 405457 44572 405523 44573
rect 260649 44568 260670 44572
rect 260734 44570 260740 44572
rect 260649 44512 260654 44568
rect 260649 44508 260670 44512
rect 260734 44510 260806 44570
rect 260734 44508 260740 44510
rect 261752 44508 261758 44572
rect 261822 44570 261828 44572
rect 261822 44510 261910 44570
rect 263869 44568 263934 44572
rect 263869 44512 263874 44568
rect 263930 44512 263934 44568
rect 261822 44508 261828 44510
rect 263869 44508 263934 44512
rect 263998 44570 264004 44572
rect 263998 44510 264026 44570
rect 263998 44508 264004 44510
rect 305952 44508 305958 44572
rect 306022 44508 306028 44572
rect 308489 44568 308542 44572
rect 308606 44570 308612 44572
rect 308489 44512 308494 44568
rect 308489 44508 308542 44512
rect 308606 44510 308646 44570
rect 404169 44568 404214 44572
rect 404278 44570 404284 44572
rect 405432 44570 405438 44572
rect 404169 44512 404174 44568
rect 308606 44508 308612 44510
rect 404169 44508 404214 44512
rect 404278 44510 404326 44570
rect 405366 44510 405438 44570
rect 405502 44568 405523 44572
rect 405518 44512 405523 44568
rect 404278 44508 404284 44510
rect 405432 44508 405438 44510
rect 405502 44508 405523 44512
rect 260649 44507 260715 44508
rect 261753 44507 261819 44508
rect 263869 44507 263935 44508
rect 140822 44374 140988 44434
rect 53598 44236 53604 44300
rect 53668 44298 53674 44300
rect 140822 44298 140882 44374
rect 201166 44372 201172 44436
rect 201236 44434 201242 44436
rect 305960 44434 306020 44508
rect 308489 44507 308555 44508
rect 404169 44507 404235 44508
rect 405457 44507 405523 44508
rect 406469 44572 406535 44573
rect 418153 44572 418219 44573
rect 406469 44568 406526 44572
rect 406590 44570 406596 44572
rect 418102 44570 418108 44572
rect 406469 44512 406474 44568
rect 406469 44508 406526 44512
rect 406590 44510 406626 44570
rect 418062 44510 418108 44570
rect 418172 44568 418219 44572
rect 418214 44512 418219 44568
rect 406590 44508 406596 44510
rect 418102 44508 418108 44510
rect 418172 44508 418219 44512
rect 406469 44507 406535 44508
rect 418153 44507 418219 44508
rect 420637 44572 420703 44573
rect 421741 44572 421807 44573
rect 422845 44572 422911 44573
rect 425973 44572 426039 44573
rect 439221 44572 439287 44573
rect 420637 44568 420670 44572
rect 420734 44570 420740 44572
rect 420637 44512 420642 44568
rect 420637 44508 420670 44512
rect 420734 44510 420794 44570
rect 421741 44568 421758 44572
rect 421822 44570 421828 44572
rect 422840 44570 422846 44572
rect 421741 44512 421746 44568
rect 420734 44508 420740 44510
rect 421741 44508 421758 44512
rect 421822 44510 421898 44570
rect 422754 44510 422846 44570
rect 421822 44508 421828 44510
rect 422840 44508 422846 44510
rect 422910 44508 422916 44572
rect 423520 44508 423526 44572
rect 423590 44508 423596 44572
rect 425968 44570 425974 44572
rect 425882 44510 425974 44570
rect 425968 44508 425974 44510
rect 426038 44508 426044 44572
rect 439160 44570 439166 44572
rect 439130 44510 439166 44570
rect 439230 44568 439287 44572
rect 439282 44512 439287 44568
rect 439160 44508 439166 44510
rect 439230 44508 439287 44512
rect 420637 44507 420703 44508
rect 421741 44507 421807 44508
rect 422845 44507 422911 44508
rect 201236 44374 306020 44434
rect 362217 44434 362283 44437
rect 423528 44434 423588 44508
rect 425973 44507 426039 44508
rect 439221 44507 439287 44508
rect 455873 44572 455939 44573
rect 458449 44572 458515 44573
rect 455873 44568 455894 44572
rect 455958 44570 455964 44572
rect 455873 44512 455878 44568
rect 455873 44508 455894 44512
rect 455958 44510 456030 44570
rect 458449 44568 458478 44572
rect 458542 44570 458548 44572
rect 458449 44512 458454 44568
rect 455958 44508 455964 44510
rect 458449 44508 458478 44512
rect 458542 44510 458606 44570
rect 458542 44508 458548 44510
rect 480912 44508 480918 44572
rect 480982 44508 480988 44572
rect 455873 44507 455939 44508
rect 458449 44507 458515 44508
rect 362217 44432 423588 44434
rect 362217 44376 362222 44432
rect 362278 44376 423588 44432
rect 362217 44374 423588 44376
rect 425237 44436 425303 44437
rect 425237 44432 425284 44436
rect 425348 44434 425354 44436
rect 425237 44376 425242 44432
rect 201236 44372 201242 44374
rect 362217 44371 362283 44374
rect 425237 44372 425284 44376
rect 425348 44374 425394 44434
rect 425348 44372 425354 44374
rect 425237 44371 425303 44372
rect 53668 44238 140882 44298
rect 53668 44236 53674 44238
rect 198406 44236 198412 44300
rect 198476 44298 198482 44300
rect 323342 44298 323348 44300
rect 198476 44238 323348 44298
rect 198476 44236 198482 44238
rect 323342 44236 323348 44238
rect 323412 44236 323418 44300
rect 360694 44236 360700 44300
rect 360764 44298 360770 44300
rect 480920 44298 480980 44508
rect 360764 44238 480980 44298
rect 360764 44236 360770 44238
rect 158437 44164 158503 44165
rect 160829 44164 160895 44165
rect 300853 44164 300919 44165
rect -960 44026 480 44116
rect 53230 44100 53236 44164
rect 53300 44162 53306 44164
rect 153326 44162 153332 44164
rect 53300 44102 153332 44162
rect 53300 44100 53306 44102
rect 153326 44100 153332 44102
rect 153396 44100 153402 44164
rect 158437 44160 158484 44164
rect 158548 44162 158554 44164
rect 158437 44104 158442 44160
rect 158437 44100 158484 44104
rect 158548 44102 158594 44162
rect 160829 44160 160876 44164
rect 160940 44162 160946 44164
rect 160829 44104 160834 44160
rect 158548 44100 158554 44102
rect 160829 44100 160876 44104
rect 160940 44102 160986 44162
rect 160940 44100 160946 44102
rect 206870 44100 206876 44164
rect 206940 44162 206946 44164
rect 295926 44162 295932 44164
rect 206940 44102 295932 44162
rect 206940 44100 206946 44102
rect 295926 44100 295932 44102
rect 295996 44100 296002 44164
rect 300853 44160 300900 44164
rect 300964 44162 300970 44164
rect 300853 44104 300858 44160
rect 300853 44100 300900 44104
rect 300964 44102 301010 44162
rect 300964 44100 300970 44102
rect 357934 44100 357940 44164
rect 358004 44162 358010 44164
rect 483422 44162 483428 44164
rect 358004 44102 483428 44162
rect 358004 44100 358010 44102
rect 483422 44100 483428 44102
rect 483492 44100 483498 44164
rect 158437 44099 158503 44100
rect 160829 44099 160895 44100
rect 300853 44099 300919 44100
rect 3417 44026 3483 44029
rect -960 44024 3483 44026
rect -960 43968 3422 44024
rect 3478 43968 3483 44024
rect -960 43966 3483 43968
rect -960 43876 480 43966
rect 3417 43963 3483 43966
rect 52310 43964 52316 44028
rect 52380 44026 52386 44028
rect 150934 44026 150940 44028
rect 52380 43966 150940 44026
rect 52380 43964 52386 43966
rect 150934 43964 150940 43966
rect 151004 43964 151010 44028
rect 202638 43964 202644 44028
rect 202708 44026 202714 44028
rect 290958 44026 290964 44028
rect 202708 43966 290964 44026
rect 202708 43964 202714 43966
rect 290958 43964 290964 43966
rect 291028 43964 291034 44028
rect 364926 43964 364932 44028
rect 364996 44026 365002 44028
rect 478454 44026 478460 44028
rect 364996 43966 478460 44026
rect 364996 43964 365002 43966
rect 478454 43964 478460 43966
rect 478524 43964 478530 44028
rect 279233 43892 279299 43893
rect 50838 43828 50844 43892
rect 50908 43890 50914 43892
rect 148542 43890 148548 43892
rect 50908 43830 148548 43890
rect 50908 43828 50914 43830
rect 148542 43828 148548 43830
rect 148612 43828 148618 43892
rect 198590 43828 198596 43892
rect 198660 43890 198666 43892
rect 279182 43890 279188 43892
rect 198660 43830 279066 43890
rect 279142 43830 279188 43890
rect 279252 43888 279299 43892
rect 279294 43832 279299 43888
rect 198660 43828 198666 43830
rect 115933 43756 115999 43757
rect 46422 43692 46428 43756
rect 46492 43754 46498 43756
rect 111006 43754 111012 43756
rect 46492 43694 111012 43754
rect 46492 43692 46498 43694
rect 111006 43692 111012 43694
rect 111076 43692 111082 43756
rect 115933 43752 115980 43756
rect 116044 43754 116050 43756
rect 115933 43696 115938 43752
rect 115933 43692 115980 43696
rect 116044 43694 116090 43754
rect 116044 43692 116050 43694
rect 197854 43692 197860 43756
rect 197924 43754 197930 43756
rect 278446 43754 278452 43756
rect 197924 43694 278452 43754
rect 197924 43692 197930 43694
rect 278446 43692 278452 43694
rect 278516 43692 278522 43756
rect 279006 43754 279066 43830
rect 279182 43828 279188 43830
rect 279252 43828 279299 43832
rect 367686 43828 367692 43892
rect 367756 43890 367762 43892
rect 468518 43890 468524 43892
rect 367756 43830 468524 43890
rect 367756 43828 367762 43830
rect 468518 43828 468524 43830
rect 468588 43828 468594 43892
rect 279233 43827 279299 43828
rect 285990 43754 285996 43756
rect 279006 43694 285996 43754
rect 285990 43692 285996 43694
rect 286060 43692 286066 43756
rect 374494 43692 374500 43756
rect 374564 43754 374570 43756
rect 473486 43754 473492 43756
rect 374564 43694 473492 43754
rect 374564 43692 374570 43694
rect 473486 43692 473492 43694
rect 473556 43692 473562 43756
rect 115933 43691 115999 43692
rect 59302 43556 59308 43620
rect 59372 43618 59378 43620
rect 123518 43618 123524 43620
rect 59372 43558 123524 43618
rect 59372 43556 59378 43558
rect 123518 43556 123524 43558
rect 123588 43556 123594 43620
rect 201350 43556 201356 43620
rect 201420 43618 201426 43620
rect 280838 43618 280844 43620
rect 201420 43558 280844 43618
rect 201420 43556 201426 43558
rect 280838 43556 280844 43558
rect 280908 43556 280914 43620
rect 371734 43556 371740 43620
rect 371804 43618 371810 43620
rect 371804 43558 451290 43618
rect 371804 43556 371810 43558
rect 407573 43484 407639 43485
rect 421005 43484 421071 43485
rect 428181 43484 428247 43485
rect 57094 43420 57100 43484
rect 57164 43482 57170 43484
rect 105302 43482 105308 43484
rect 57164 43422 105308 43482
rect 57164 43420 57170 43422
rect 105302 43420 105308 43422
rect 105372 43420 105378 43484
rect 204846 43420 204852 43484
rect 204916 43482 204922 43484
rect 273478 43482 273484 43484
rect 204916 43422 273484 43482
rect 204916 43420 204922 43422
rect 273478 43420 273484 43422
rect 273548 43420 273554 43484
rect 407573 43480 407620 43484
rect 407684 43482 407690 43484
rect 407573 43424 407578 43480
rect 407573 43420 407620 43424
rect 407684 43422 407730 43482
rect 421005 43480 421052 43484
rect 421116 43482 421122 43484
rect 421005 43424 421010 43480
rect 407684 43420 407690 43422
rect 421005 43420 421052 43424
rect 421116 43422 421162 43482
rect 428181 43480 428228 43484
rect 428292 43482 428298 43484
rect 451230 43482 451290 43558
rect 463550 43482 463556 43484
rect 428181 43424 428186 43480
rect 421116 43420 421122 43422
rect 428181 43420 428228 43424
rect 428292 43422 428338 43482
rect 451230 43422 463556 43482
rect 428292 43420 428298 43422
rect 463550 43420 463556 43422
rect 463620 43420 463626 43484
rect 407573 43419 407639 43420
rect 421005 43419 421071 43420
rect 428181 43419 428247 43420
rect 59118 43284 59124 43348
rect 59188 43346 59194 43348
rect 101070 43346 101076 43348
rect 59188 43286 101076 43346
rect 59188 43284 59194 43286
rect 101070 43284 101076 43286
rect 101140 43284 101146 43348
rect 200614 43284 200620 43348
rect 200684 43346 200690 43348
rect 265934 43346 265940 43348
rect 200684 43286 265940 43346
rect 200684 43284 200690 43286
rect 265934 43284 265940 43286
rect 266004 43284 266010 43348
rect 85389 43212 85455 43213
rect 92381 43212 92447 43213
rect 95877 43212 95943 43213
rect 128353 43212 128419 43213
rect 85389 43208 85436 43212
rect 85500 43210 85506 43212
rect 85389 43152 85394 43208
rect 85389 43148 85436 43152
rect 85500 43150 85546 43210
rect 92381 43208 92428 43212
rect 92492 43210 92498 43212
rect 92381 43152 92386 43208
rect 85500 43148 85506 43150
rect 92381 43148 92428 43152
rect 92492 43150 92538 43210
rect 95877 43208 95924 43212
rect 95988 43210 95994 43212
rect 128302 43210 128308 43212
rect 95877 43152 95882 43208
rect 92492 43148 92498 43150
rect 95877 43148 95924 43152
rect 95988 43150 96034 43210
rect 128262 43150 128308 43210
rect 128372 43208 128419 43212
rect 128414 43152 128419 43208
rect 95988 43148 95994 43150
rect 128302 43148 128308 43150
rect 128372 43148 128419 43152
rect 85389 43147 85455 43148
rect 92381 43147 92447 43148
rect 95877 43147 95943 43148
rect 128353 43147 128419 43148
rect 265157 43212 265223 43213
rect 272149 43212 272215 43213
rect 325877 43212 325943 43213
rect 398189 43212 398255 43213
rect 401685 43212 401751 43213
rect 265157 43208 265204 43212
rect 265268 43210 265274 43212
rect 265157 43152 265162 43208
rect 265157 43148 265204 43152
rect 265268 43150 265314 43210
rect 272149 43208 272196 43212
rect 272260 43210 272266 43212
rect 272149 43152 272154 43208
rect 265268 43148 265274 43150
rect 272149 43148 272196 43152
rect 272260 43150 272306 43210
rect 325877 43208 325924 43212
rect 325988 43210 325994 43212
rect 325877 43152 325882 43208
rect 272260 43148 272266 43150
rect 325877 43148 325924 43152
rect 325988 43150 326034 43210
rect 398189 43208 398236 43212
rect 398300 43210 398306 43212
rect 398189 43152 398194 43208
rect 325988 43148 325994 43150
rect 398189 43148 398236 43152
rect 398300 43150 398346 43210
rect 401685 43208 401732 43212
rect 401796 43210 401802 43212
rect 401685 43152 401690 43208
rect 398300 43148 398306 43150
rect 401685 43148 401732 43152
rect 401796 43150 401842 43210
rect 401796 43148 401802 43150
rect 265157 43147 265223 43148
rect 272149 43147 272215 43148
rect 325877 43147 325943 43148
rect 398189 43147 398255 43148
rect 401685 43147 401751 43148
rect 76005 42804 76071 42805
rect 78213 42804 78279 42805
rect 80421 42804 80487 42805
rect 86493 42804 86559 42805
rect 87597 42804 87663 42805
rect 88333 42804 88399 42805
rect 76005 42800 76052 42804
rect 76116 42802 76122 42804
rect 76005 42744 76010 42800
rect 76005 42740 76052 42744
rect 76116 42742 76162 42802
rect 78213 42800 78260 42804
rect 78324 42802 78330 42804
rect 78213 42744 78218 42800
rect 76116 42740 76122 42742
rect 78213 42740 78260 42744
rect 78324 42742 78370 42802
rect 80421 42800 80468 42804
rect 80532 42802 80538 42804
rect 80421 42744 80426 42800
rect 78324 42740 78330 42742
rect 80421 42740 80468 42744
rect 80532 42742 80578 42802
rect 86493 42800 86540 42804
rect 86604 42802 86610 42804
rect 86493 42744 86498 42800
rect 80532 42740 80538 42742
rect 86493 42740 86540 42744
rect 86604 42742 86650 42802
rect 87597 42800 87644 42804
rect 87708 42802 87714 42804
rect 87597 42744 87602 42800
rect 86604 42740 86610 42742
rect 87597 42740 87644 42744
rect 87708 42742 87754 42802
rect 88333 42800 88380 42804
rect 88444 42802 88450 42804
rect 88609 42802 88675 42805
rect 90725 42804 90791 42805
rect 91277 42804 91343 42805
rect 93301 42804 93367 42805
rect 93669 42804 93735 42805
rect 96245 42804 96311 42805
rect 106365 42804 106431 42805
rect 88742 42802 88748 42804
rect 88333 42744 88338 42800
rect 87708 42740 87714 42742
rect 88333 42740 88380 42744
rect 88444 42742 88490 42802
rect 88609 42800 88748 42802
rect 88609 42744 88614 42800
rect 88670 42744 88748 42800
rect 88609 42742 88748 42744
rect 88444 42740 88450 42742
rect 76005 42739 76071 42740
rect 78213 42739 78279 42740
rect 80421 42739 80487 42740
rect 86493 42739 86559 42740
rect 87597 42739 87663 42740
rect 88333 42739 88399 42740
rect 88609 42739 88675 42742
rect 88742 42740 88748 42742
rect 88812 42740 88818 42804
rect 90725 42800 90772 42804
rect 90836 42802 90842 42804
rect 90725 42744 90730 42800
rect 90725 42740 90772 42744
rect 90836 42742 90882 42802
rect 91277 42800 91324 42804
rect 91388 42802 91394 42804
rect 93301 42802 93348 42804
rect 91277 42744 91282 42800
rect 90836 42740 90842 42742
rect 91277 42740 91324 42744
rect 91388 42742 91434 42802
rect 93256 42800 93348 42802
rect 93256 42744 93306 42800
rect 93256 42742 93348 42744
rect 91388 42740 91394 42742
rect 93301 42740 93348 42742
rect 93412 42740 93418 42804
rect 93669 42800 93716 42804
rect 93780 42802 93786 42804
rect 93669 42744 93674 42800
rect 93669 42740 93716 42744
rect 93780 42742 93826 42802
rect 96245 42800 96292 42804
rect 96356 42802 96362 42804
rect 96245 42744 96250 42800
rect 93780 42740 93786 42742
rect 96245 42740 96292 42744
rect 96356 42742 96402 42802
rect 106365 42800 106412 42804
rect 106476 42802 106482 42804
rect 107009 42802 107075 42805
rect 108573 42804 108639 42805
rect 107510 42802 107516 42804
rect 106365 42744 106370 42800
rect 96356 42740 96362 42742
rect 106365 42740 106412 42744
rect 106476 42742 106522 42802
rect 107009 42800 107516 42802
rect 107009 42744 107014 42800
rect 107070 42744 107516 42800
rect 107009 42742 107516 42744
rect 106476 42740 106482 42742
rect 90725 42739 90791 42740
rect 91277 42739 91343 42740
rect 93301 42739 93367 42740
rect 93669 42739 93735 42740
rect 96245 42739 96311 42740
rect 106365 42739 106431 42740
rect 107009 42739 107075 42742
rect 107510 42740 107516 42742
rect 107580 42740 107586 42804
rect 108573 42800 108620 42804
rect 108684 42802 108690 42804
rect 111885 42802 111951 42805
rect 113173 42804 113239 42805
rect 112110 42802 112116 42804
rect 108573 42744 108578 42800
rect 108573 42740 108620 42744
rect 108684 42742 108730 42802
rect 111885 42800 112116 42802
rect 111885 42744 111890 42800
rect 111946 42744 112116 42800
rect 111885 42742 112116 42744
rect 108684 42740 108690 42742
rect 108573 42739 108639 42740
rect 111885 42739 111951 42742
rect 112110 42740 112116 42742
rect 112180 42740 112186 42804
rect 113173 42800 113220 42804
rect 113284 42802 113290 42804
rect 114185 42802 114251 42805
rect 115749 42804 115815 42805
rect 114318 42802 114324 42804
rect 113173 42744 113178 42800
rect 113173 42740 113220 42744
rect 113284 42742 113330 42802
rect 114185 42800 114324 42802
rect 114185 42744 114190 42800
rect 114246 42744 114324 42800
rect 114185 42742 114324 42744
rect 113284 42740 113290 42742
rect 113173 42739 113239 42740
rect 114185 42739 114251 42742
rect 114318 42740 114324 42742
rect 114388 42740 114394 42804
rect 115749 42800 115796 42804
rect 115860 42802 115866 42804
rect 116301 42802 116367 42805
rect 116894 42802 116900 42804
rect 115749 42744 115754 42800
rect 115749 42740 115796 42744
rect 115860 42742 115906 42802
rect 116301 42800 116900 42802
rect 116301 42744 116306 42800
rect 116362 42744 116900 42800
rect 116301 42742 116900 42744
rect 115860 42740 115866 42742
rect 115749 42739 115815 42740
rect 116301 42739 116367 42742
rect 116894 42740 116900 42742
rect 116964 42740 116970 42804
rect 118233 42802 118299 42805
rect 119061 42804 119127 42805
rect 133413 42804 133479 42805
rect 118366 42802 118372 42804
rect 118233 42800 118372 42802
rect 118233 42744 118238 42800
rect 118294 42744 118372 42800
rect 118233 42742 118372 42744
rect 118233 42739 118299 42742
rect 118366 42740 118372 42742
rect 118436 42740 118442 42804
rect 119061 42800 119108 42804
rect 119172 42802 119178 42804
rect 119061 42744 119066 42800
rect 119061 42740 119108 42744
rect 119172 42742 119218 42802
rect 133413 42800 133460 42804
rect 133524 42802 133530 42804
rect 135897 42802 135963 42805
rect 155953 42804 156019 42805
rect 136030 42802 136036 42804
rect 133413 42744 133418 42800
rect 119172 42740 119178 42742
rect 133413 42740 133460 42744
rect 133524 42742 133570 42802
rect 135897 42800 136036 42802
rect 135897 42744 135902 42800
rect 135958 42744 136036 42800
rect 135897 42742 136036 42744
rect 133524 42740 133530 42742
rect 119061 42739 119127 42740
rect 133413 42739 133479 42740
rect 135897 42739 135963 42742
rect 136030 42740 136036 42742
rect 136100 42740 136106 42804
rect 155902 42802 155908 42804
rect 155862 42742 155908 42802
rect 155972 42800 156019 42804
rect 156014 42744 156019 42800
rect 155902 42740 155908 42742
rect 155972 42740 156019 42744
rect 155953 42739 156019 42740
rect 183461 42804 183527 42805
rect 238109 42804 238175 42805
rect 183461 42800 183508 42804
rect 183572 42802 183578 42804
rect 183461 42744 183466 42800
rect 183461 42740 183508 42744
rect 183572 42742 183618 42802
rect 238109 42800 238156 42804
rect 238220 42802 238226 42804
rect 239121 42802 239187 42805
rect 240501 42804 240567 42805
rect 241605 42804 241671 42805
rect 245285 42804 245351 42805
rect 246389 42804 246455 42805
rect 250069 42804 250135 42805
rect 251173 42804 251239 42805
rect 253381 42804 253447 42805
rect 260925 42804 260991 42805
rect 239254 42802 239260 42804
rect 238109 42744 238114 42800
rect 183572 42740 183578 42742
rect 238109 42740 238156 42744
rect 238220 42742 238266 42802
rect 239121 42800 239260 42802
rect 239121 42744 239126 42800
rect 239182 42744 239260 42800
rect 239121 42742 239260 42744
rect 238220 42740 238226 42742
rect 183461 42739 183527 42740
rect 238109 42739 238175 42740
rect 239121 42739 239187 42742
rect 239254 42740 239260 42742
rect 239324 42740 239330 42804
rect 240501 42800 240548 42804
rect 240612 42802 240618 42804
rect 240501 42744 240506 42800
rect 240501 42740 240548 42744
rect 240612 42742 240658 42802
rect 241605 42800 241652 42804
rect 241716 42802 241722 42804
rect 241605 42744 241610 42800
rect 240612 42740 240618 42742
rect 241605 42740 241652 42744
rect 241716 42742 241762 42802
rect 245285 42800 245332 42804
rect 245396 42802 245402 42804
rect 245285 42744 245290 42800
rect 241716 42740 241722 42742
rect 245285 42740 245332 42744
rect 245396 42742 245442 42802
rect 246389 42800 246436 42804
rect 246500 42802 246506 42804
rect 246389 42744 246394 42800
rect 245396 42740 245402 42742
rect 246389 42740 246436 42744
rect 246500 42742 246546 42802
rect 250069 42800 250116 42804
rect 250180 42802 250186 42804
rect 250069 42744 250074 42800
rect 246500 42740 246506 42742
rect 250069 42740 250116 42744
rect 250180 42742 250226 42802
rect 251173 42800 251220 42804
rect 251284 42802 251290 42804
rect 251173 42744 251178 42800
rect 250180 42740 250186 42742
rect 251173 42740 251220 42744
rect 251284 42742 251330 42802
rect 253381 42800 253428 42804
rect 253492 42802 253498 42804
rect 253381 42744 253386 42800
rect 251284 42740 251290 42742
rect 253381 42740 253428 42744
rect 253492 42742 253538 42802
rect 260925 42800 260972 42804
rect 261036 42802 261042 42804
rect 268193 42802 268259 42805
rect 268326 42802 268332 42804
rect 260925 42744 260930 42800
rect 253492 42740 253498 42742
rect 260925 42740 260972 42744
rect 261036 42742 261082 42802
rect 268193 42800 268332 42802
rect 268193 42744 268198 42800
rect 268254 42744 268332 42800
rect 268193 42742 268332 42744
rect 261036 42740 261042 42742
rect 240501 42739 240567 42740
rect 241605 42739 241671 42740
rect 245285 42739 245351 42740
rect 246389 42739 246455 42740
rect 250069 42739 250135 42740
rect 251173 42739 251239 42740
rect 253381 42739 253447 42740
rect 260925 42739 260991 42740
rect 268193 42739 268259 42742
rect 268326 42740 268332 42742
rect 268396 42740 268402 42804
rect 268469 42802 268535 42805
rect 271229 42804 271295 42805
rect 273253 42804 273319 42805
rect 268694 42802 268700 42804
rect 268469 42800 268700 42802
rect 268469 42744 268474 42800
rect 268530 42744 268700 42800
rect 268469 42742 268700 42744
rect 268469 42739 268535 42742
rect 268694 42740 268700 42742
rect 268764 42740 268770 42804
rect 271229 42800 271276 42804
rect 271340 42802 271346 42804
rect 271229 42744 271234 42800
rect 271229 42740 271276 42744
rect 271340 42742 271386 42802
rect 273253 42800 273300 42804
rect 273364 42802 273370 42804
rect 276105 42802 276171 42805
rect 276933 42804 276999 42805
rect 276238 42802 276244 42804
rect 273253 42744 273258 42800
rect 271340 42740 271346 42742
rect 273253 42740 273300 42744
rect 273364 42742 273410 42802
rect 276105 42800 276244 42802
rect 276105 42744 276110 42800
rect 276166 42744 276244 42800
rect 276105 42742 276244 42744
rect 273364 42740 273370 42742
rect 271229 42739 271295 42740
rect 273253 42739 273319 42740
rect 276105 42739 276171 42742
rect 276238 42740 276244 42742
rect 276308 42740 276314 42804
rect 276933 42800 276980 42804
rect 277044 42802 277050 42804
rect 276933 42744 276938 42800
rect 276933 42740 276980 42744
rect 277044 42742 277090 42802
rect 277044 42740 277050 42742
rect 278078 42740 278084 42804
rect 278148 42802 278154 42804
rect 278313 42802 278379 42805
rect 278148 42800 278379 42802
rect 278148 42744 278318 42800
rect 278374 42744 278379 42800
rect 278148 42742 278379 42744
rect 278148 42740 278154 42742
rect 276933 42739 276999 42740
rect 278313 42739 278379 42742
rect 293309 42804 293375 42805
rect 298461 42804 298527 42805
rect 293309 42800 293356 42804
rect 293420 42802 293426 42804
rect 293309 42744 293314 42800
rect 293309 42740 293356 42744
rect 293420 42742 293466 42802
rect 298461 42800 298508 42804
rect 298572 42802 298578 42804
rect 302509 42802 302575 42805
rect 310973 42804 311039 42805
rect 313365 42804 313431 42805
rect 318333 42804 318399 42805
rect 320909 42804 320975 42805
rect 343173 42804 343239 42805
rect 343449 42804 343515 42805
rect 303470 42802 303476 42804
rect 298461 42744 298466 42800
rect 293420 42740 293426 42742
rect 298461 42740 298508 42744
rect 298572 42742 298618 42802
rect 302509 42800 303476 42802
rect 302509 42744 302514 42800
rect 302570 42744 303476 42800
rect 302509 42742 303476 42744
rect 298572 42740 298578 42742
rect 293309 42739 293375 42740
rect 298461 42739 298527 42740
rect 302509 42739 302575 42742
rect 303470 42740 303476 42742
rect 303540 42740 303546 42804
rect 310973 42800 311020 42804
rect 311084 42802 311090 42804
rect 310973 42744 310978 42800
rect 310973 42740 311020 42744
rect 311084 42742 311130 42802
rect 313365 42800 313412 42804
rect 313476 42802 313482 42804
rect 313365 42744 313370 42800
rect 311084 42740 311090 42742
rect 313365 42740 313412 42744
rect 313476 42742 313522 42802
rect 318333 42800 318380 42804
rect 318444 42802 318450 42804
rect 318333 42744 318338 42800
rect 313476 42740 313482 42742
rect 318333 42740 318380 42744
rect 318444 42742 318490 42802
rect 320909 42800 320956 42804
rect 321020 42802 321026 42804
rect 343173 42802 343220 42804
rect 320909 42744 320914 42800
rect 318444 42740 318450 42742
rect 320909 42740 320956 42744
rect 321020 42742 321066 42802
rect 343128 42800 343220 42802
rect 343128 42744 343178 42800
rect 343128 42742 343220 42744
rect 321020 42740 321026 42742
rect 343173 42740 343220 42742
rect 343284 42740 343290 42804
rect 343398 42802 343404 42804
rect 343358 42742 343404 42802
rect 343468 42800 343515 42804
rect 343510 42744 343515 42800
rect 343398 42740 343404 42742
rect 343468 42740 343515 42744
rect 310973 42739 311039 42740
rect 313365 42739 313431 42740
rect 318333 42739 318399 42740
rect 320909 42739 320975 42740
rect 343173 42739 343239 42740
rect 343449 42739 343515 42740
rect 399385 42802 399451 42805
rect 408309 42804 408375 42805
rect 408677 42804 408743 42805
rect 409965 42804 410031 42805
rect 411253 42804 411319 42805
rect 399518 42802 399524 42804
rect 399385 42800 399524 42802
rect 399385 42744 399390 42800
rect 399446 42744 399524 42800
rect 399385 42742 399524 42744
rect 399385 42739 399451 42742
rect 399518 42740 399524 42742
rect 399588 42740 399594 42804
rect 408309 42800 408356 42804
rect 408420 42802 408426 42804
rect 408309 42744 408314 42800
rect 408309 42740 408356 42744
rect 408420 42742 408466 42802
rect 408677 42800 408724 42804
rect 408788 42802 408794 42804
rect 408677 42744 408682 42800
rect 408420 42740 408426 42742
rect 408677 42740 408724 42744
rect 408788 42742 408834 42802
rect 409965 42800 410012 42804
rect 410076 42802 410082 42804
rect 409965 42744 409970 42800
rect 408788 42740 408794 42742
rect 409965 42740 410012 42744
rect 410076 42742 410122 42802
rect 411253 42800 411300 42804
rect 411364 42802 411370 42804
rect 411897 42802 411963 42805
rect 413277 42804 413343 42805
rect 413645 42804 413711 42805
rect 415485 42804 415551 42805
rect 426433 42804 426499 42805
rect 412398 42802 412404 42804
rect 411253 42744 411258 42800
rect 410076 42740 410082 42742
rect 411253 42740 411300 42744
rect 411364 42742 411410 42802
rect 411897 42800 412404 42802
rect 411897 42744 411902 42800
rect 411958 42744 412404 42800
rect 411897 42742 412404 42744
rect 411364 42740 411370 42742
rect 408309 42739 408375 42740
rect 408677 42739 408743 42740
rect 409965 42739 410031 42740
rect 411253 42739 411319 42740
rect 411897 42739 411963 42742
rect 412398 42740 412404 42742
rect 412468 42740 412474 42804
rect 413277 42802 413324 42804
rect 413232 42800 413324 42802
rect 413232 42744 413282 42800
rect 413232 42742 413324 42744
rect 413277 42740 413324 42742
rect 413388 42740 413394 42804
rect 413645 42800 413692 42804
rect 413756 42802 413762 42804
rect 413645 42744 413650 42800
rect 413645 42740 413692 42744
rect 413756 42742 413802 42802
rect 415485 42800 415532 42804
rect 415596 42802 415602 42804
rect 426382 42802 426388 42804
rect 415485 42744 415490 42800
rect 413756 42740 413762 42742
rect 415485 42740 415532 42744
rect 415596 42742 415642 42802
rect 426342 42742 426388 42802
rect 426452 42800 426499 42804
rect 426494 42744 426499 42800
rect 415596 42740 415602 42742
rect 426382 42740 426388 42742
rect 426452 42740 426499 42744
rect 413277 42739 413343 42740
rect 413645 42739 413711 42740
rect 415485 42739 415551 42740
rect 426433 42739 426499 42740
rect 427629 42804 427695 42805
rect 428549 42804 428615 42805
rect 429653 42804 429719 42805
rect 430941 42804 431007 42805
rect 427629 42800 427676 42804
rect 427740 42802 427746 42804
rect 427629 42744 427634 42800
rect 427629 42740 427676 42744
rect 427740 42742 427786 42802
rect 428549 42800 428596 42804
rect 428660 42802 428666 42804
rect 428549 42744 428554 42800
rect 427740 42740 427746 42742
rect 428549 42740 428596 42744
rect 428660 42742 428706 42802
rect 429653 42800 429700 42804
rect 429764 42802 429770 42804
rect 429653 42744 429658 42800
rect 428660 42740 428666 42742
rect 429653 42740 429700 42744
rect 429764 42742 429810 42802
rect 430941 42800 430988 42804
rect 431052 42802 431058 42804
rect 432137 42802 432203 42805
rect 433333 42804 433399 42805
rect 434621 42804 434687 42805
rect 435909 42804 435975 42805
rect 432270 42802 432276 42804
rect 430941 42744 430946 42800
rect 429764 42740 429770 42742
rect 430941 42740 430988 42744
rect 431052 42742 431098 42802
rect 432137 42800 432276 42802
rect 432137 42744 432142 42800
rect 432198 42744 432276 42800
rect 432137 42742 432276 42744
rect 431052 42740 431058 42742
rect 427629 42739 427695 42740
rect 428549 42739 428615 42740
rect 429653 42739 429719 42740
rect 430941 42739 431007 42740
rect 432137 42739 432203 42742
rect 432270 42740 432276 42742
rect 432340 42740 432346 42804
rect 433333 42800 433380 42804
rect 433444 42802 433450 42804
rect 433333 42744 433338 42800
rect 433333 42740 433380 42744
rect 433444 42742 433490 42802
rect 434621 42800 434668 42804
rect 434732 42802 434738 42804
rect 434621 42744 434626 42800
rect 433444 42740 433450 42742
rect 434621 42740 434668 42744
rect 434732 42742 434778 42802
rect 435909 42800 435956 42804
rect 436020 42802 436026 42804
rect 436369 42802 436435 42805
rect 438485 42804 438551 42805
rect 440877 42804 440943 42805
rect 443453 42804 443519 42805
rect 445845 42804 445911 42805
rect 448237 42804 448303 42805
rect 453389 42804 453455 42805
rect 485957 42804 486023 42805
rect 436870 42802 436876 42804
rect 435909 42744 435914 42800
rect 434732 42740 434738 42742
rect 435909 42740 435956 42744
rect 436020 42742 436066 42802
rect 436369 42800 436876 42802
rect 436369 42744 436374 42800
rect 436430 42744 436876 42800
rect 436369 42742 436876 42744
rect 436020 42740 436026 42742
rect 433333 42739 433399 42740
rect 434621 42739 434687 42740
rect 435909 42739 435975 42740
rect 436369 42739 436435 42742
rect 436870 42740 436876 42742
rect 436940 42740 436946 42804
rect 438485 42800 438532 42804
rect 438596 42802 438602 42804
rect 438485 42744 438490 42800
rect 438485 42740 438532 42744
rect 438596 42742 438642 42802
rect 440877 42800 440924 42804
rect 440988 42802 440994 42804
rect 440877 42744 440882 42800
rect 438596 42740 438602 42742
rect 440877 42740 440924 42744
rect 440988 42742 441034 42802
rect 443453 42800 443500 42804
rect 443564 42802 443570 42804
rect 443453 42744 443458 42800
rect 440988 42740 440994 42742
rect 443453 42740 443500 42744
rect 443564 42742 443610 42802
rect 445845 42800 445892 42804
rect 445956 42802 445962 42804
rect 445845 42744 445850 42800
rect 443564 42740 443570 42742
rect 445845 42740 445892 42744
rect 445956 42742 446002 42802
rect 448237 42800 448284 42804
rect 448348 42802 448354 42804
rect 448237 42744 448242 42800
rect 445956 42740 445962 42742
rect 448237 42740 448284 42744
rect 448348 42742 448394 42802
rect 453389 42800 453436 42804
rect 453500 42802 453506 42804
rect 453389 42744 453394 42800
rect 448348 42740 448354 42742
rect 453389 42740 453436 42744
rect 453500 42742 453546 42802
rect 485957 42800 486004 42804
rect 486068 42802 486074 42804
rect 485957 42744 485962 42800
rect 453500 42740 453506 42742
rect 485957 42740 486004 42744
rect 486068 42742 486114 42802
rect 486068 42740 486074 42742
rect 503110 42740 503116 42804
rect 503180 42802 503186 42804
rect 503253 42802 503319 42805
rect 503529 42804 503595 42805
rect 503180 42800 503319 42802
rect 503180 42744 503258 42800
rect 503314 42744 503319 42800
rect 503180 42742 503319 42744
rect 503180 42740 503186 42742
rect 438485 42739 438551 42740
rect 440877 42739 440943 42740
rect 443453 42739 443519 42740
rect 445845 42739 445911 42740
rect 448237 42739 448303 42740
rect 453389 42739 453455 42740
rect 485957 42739 486023 42740
rect 503253 42739 503319 42742
rect 503478 42740 503484 42804
rect 503548 42802 503595 42804
rect 503548 42800 503640 42802
rect 503590 42744 503640 42800
rect 503548 42742 503640 42744
rect 503548 42740 503595 42742
rect 503529 42739 503595 42740
rect 183185 42668 183251 42669
rect 60222 42604 60228 42668
rect 60292 42666 60298 42668
rect 125910 42666 125916 42668
rect 60292 42606 125916 42666
rect 60292 42604 60298 42606
rect 125910 42604 125916 42606
rect 125980 42604 125986 42668
rect 183134 42666 183140 42668
rect 183094 42606 183140 42666
rect 183204 42664 183251 42668
rect 183246 42608 183251 42664
rect 183134 42604 183140 42606
rect 183204 42604 183251 42608
rect 215886 42604 215892 42668
rect 215956 42666 215962 42668
rect 288198 42666 288204 42668
rect 215956 42606 288204 42666
rect 215956 42604 215962 42606
rect 288198 42604 288204 42606
rect 288268 42604 288274 42668
rect 370446 42604 370452 42668
rect 370516 42666 370522 42668
rect 465942 42666 465948 42668
rect 370516 42606 465948 42666
rect 370516 42604 370522 42606
rect 465942 42604 465948 42606
rect 466012 42604 466018 42668
rect 183185 42603 183251 42604
rect 165797 42532 165863 42533
rect 54886 42468 54892 42532
rect 54956 42530 54962 42532
rect 120758 42530 120764 42532
rect 54956 42470 120764 42530
rect 54956 42468 54962 42470
rect 120758 42468 120764 42470
rect 120828 42468 120834 42532
rect 165797 42528 165844 42532
rect 165908 42530 165914 42532
rect 165797 42472 165802 42528
rect 165797 42468 165844 42472
rect 165908 42470 165954 42530
rect 165908 42468 165914 42470
rect 210366 42468 210372 42532
rect 210436 42530 210442 42532
rect 270902 42530 270908 42532
rect 210436 42470 270908 42530
rect 210436 42468 210442 42470
rect 270902 42468 270908 42470
rect 270972 42468 270978 42532
rect 376150 42468 376156 42532
rect 376220 42530 376226 42532
rect 470910 42530 470916 42532
rect 376220 42470 470916 42530
rect 376220 42468 376226 42470
rect 470910 42468 470916 42470
rect 470980 42468 470986 42532
rect 165797 42467 165863 42468
rect 266353 42396 266419 42397
rect 57830 42332 57836 42396
rect 57900 42394 57906 42396
rect 117998 42394 118004 42396
rect 57900 42334 118004 42394
rect 57900 42332 57906 42334
rect 117998 42332 118004 42334
rect 118068 42332 118074 42396
rect 214414 42332 214420 42396
rect 214484 42394 214490 42396
rect 263542 42394 263548 42396
rect 214484 42334 263548 42394
rect 214484 42332 214490 42334
rect 263542 42332 263548 42334
rect 263612 42332 263618 42396
rect 266302 42394 266308 42396
rect 266262 42334 266308 42394
rect 266372 42392 266419 42396
rect 266414 42336 266419 42392
rect 266302 42332 266308 42334
rect 266372 42332 266419 42336
rect 266353 42331 266419 42332
rect 266629 42394 266695 42397
rect 269757 42396 269823 42397
rect 267590 42394 267596 42396
rect 266629 42392 267596 42394
rect 266629 42336 266634 42392
rect 266690 42336 267596 42392
rect 266629 42334 267596 42336
rect 266629 42331 266695 42334
rect 267590 42332 267596 42334
rect 267660 42332 267666 42396
rect 269757 42392 269804 42396
rect 269868 42394 269874 42396
rect 269757 42336 269762 42392
rect 269757 42332 269804 42336
rect 269868 42334 269914 42394
rect 269868 42332 269874 42334
rect 378726 42332 378732 42396
rect 378796 42394 378802 42396
rect 460974 42394 460980 42396
rect 378796 42334 460980 42394
rect 378796 42332 378802 42334
rect 460974 42332 460980 42334
rect 461044 42332 461050 42396
rect 269757 42331 269823 42332
rect 58934 42196 58940 42260
rect 59004 42258 59010 42260
rect 105854 42258 105860 42260
rect 59004 42198 105860 42258
rect 59004 42196 59010 42198
rect 105854 42196 105860 42198
rect 105924 42196 105930 42260
rect 109309 42258 109375 42261
rect 111149 42260 111215 42261
rect 109534 42258 109540 42260
rect 109309 42256 109540 42258
rect 109309 42200 109314 42256
rect 109370 42200 109540 42256
rect 109309 42198 109540 42200
rect 109309 42195 109375 42198
rect 109534 42196 109540 42198
rect 109604 42196 109610 42260
rect 111149 42256 111196 42260
rect 111260 42258 111266 42260
rect 111149 42200 111154 42256
rect 111149 42196 111196 42200
rect 111260 42198 111306 42258
rect 111260 42196 111266 42198
rect 206134 42196 206140 42260
rect 206204 42258 206210 42260
rect 255998 42258 256004 42260
rect 206204 42198 256004 42258
rect 206204 42196 206210 42198
rect 255998 42196 256004 42198
rect 256068 42196 256074 42260
rect 273529 42258 273595 42261
rect 274398 42258 274404 42260
rect 273529 42256 274404 42258
rect 273529 42200 273534 42256
rect 273590 42200 274404 42256
rect 273529 42198 274404 42200
rect 111149 42195 111215 42196
rect 273529 42195 273595 42198
rect 274398 42196 274404 42198
rect 274468 42196 274474 42260
rect 274725 42258 274791 42261
rect 275318 42258 275324 42260
rect 274725 42256 275324 42258
rect 274725 42200 274730 42256
rect 274786 42200 275324 42256
rect 274725 42198 275324 42200
rect 274725 42195 274791 42198
rect 275318 42196 275324 42198
rect 275388 42196 275394 42260
rect 374678 42196 374684 42260
rect 374748 42258 374754 42260
rect 451038 42258 451044 42260
rect 374748 42198 451044 42258
rect 374748 42196 374754 42198
rect 451038 42196 451044 42198
rect 451108 42196 451114 42260
rect 58750 42060 58756 42124
rect 58820 42122 58826 42124
rect 103830 42122 103836 42124
rect 58820 42062 103836 42122
rect 58820 42060 58826 42062
rect 103830 42060 103836 42062
rect 103900 42060 103906 42124
rect 207974 42060 207980 42124
rect 208044 42122 208050 42124
rect 253606 42122 253612 42124
rect 208044 42062 253612 42122
rect 208044 42060 208050 42062
rect 253606 42060 253612 42062
rect 253676 42060 253682 42124
rect 254117 42122 254183 42125
rect 254526 42122 254532 42124
rect 254117 42120 254532 42122
rect 254117 42064 254122 42120
rect 254178 42064 254532 42120
rect 254117 42062 254532 42064
rect 254117 42059 254183 42062
rect 254526 42060 254532 42062
rect 254596 42060 254602 42124
rect 363454 42060 363460 42124
rect 363524 42122 363530 42124
rect 433558 42122 433564 42124
rect 363524 42062 433564 42122
rect 363524 42060 363530 42062
rect 433558 42060 433564 42062
rect 433628 42060 433634 42124
rect 435173 42122 435239 42125
rect 435766 42122 435772 42124
rect 435173 42120 435772 42122
rect 435173 42064 435178 42120
rect 435234 42064 435772 42120
rect 435173 42062 435772 42064
rect 435173 42059 435239 42062
rect 435766 42060 435772 42062
rect 435836 42060 435842 42124
rect 248597 41988 248663 41989
rect 58566 41924 58572 41988
rect 58636 41986 58642 41988
rect 98494 41986 98500 41988
rect 58636 41926 98500 41986
rect 58636 41924 58642 41926
rect 98494 41924 98500 41926
rect 98564 41924 98570 41988
rect 208894 41924 208900 41988
rect 208964 41986 208970 41988
rect 248270 41986 248276 41988
rect 208964 41926 248276 41986
rect 208964 41924 208970 41926
rect 248270 41924 248276 41926
rect 248340 41924 248346 41988
rect 248597 41984 248644 41988
rect 248708 41986 248714 41988
rect 251725 41986 251791 41989
rect 431125 41988 431191 41989
rect 252318 41986 252324 41988
rect 248597 41928 248602 41984
rect 248597 41924 248644 41928
rect 248708 41926 248754 41986
rect 251725 41984 252324 41986
rect 251725 41928 251730 41984
rect 251786 41928 252324 41984
rect 251725 41926 252324 41928
rect 248708 41924 248714 41926
rect 248597 41923 248663 41924
rect 251725 41923 251791 41926
rect 252318 41924 252324 41926
rect 252388 41924 252394 41988
rect 375966 41924 375972 41988
rect 376036 41986 376042 41988
rect 416630 41986 416636 41988
rect 376036 41926 416636 41986
rect 376036 41924 376042 41926
rect 416630 41924 416636 41926
rect 416700 41924 416706 41988
rect 431125 41984 431172 41988
rect 431236 41986 431242 41988
rect 431125 41928 431130 41984
rect 431125 41924 431172 41928
rect 431236 41926 431282 41986
rect 431236 41924 431242 41926
rect 431125 41923 431191 41924
rect 78765 41850 78831 41853
rect 79542 41850 79548 41852
rect 78765 41848 79548 41850
rect 78765 41792 78770 41848
rect 78826 41792 79548 41848
rect 78765 41790 79548 41792
rect 78765 41787 78831 41790
rect 79542 41788 79548 41790
rect 79612 41788 79618 41852
rect 81801 41850 81867 41853
rect 89989 41852 90055 41853
rect 247677 41852 247743 41853
rect 81934 41850 81940 41852
rect 81801 41848 81940 41850
rect 81801 41792 81806 41848
rect 81862 41792 81940 41848
rect 81801 41790 81940 41792
rect 81801 41787 81867 41790
rect 81934 41788 81940 41790
rect 82004 41788 82010 41852
rect 89989 41848 90036 41852
rect 90100 41850 90106 41852
rect 89989 41792 89994 41848
rect 89989 41788 90036 41792
rect 90100 41790 90146 41850
rect 247677 41848 247724 41852
rect 247788 41850 247794 41852
rect 400305 41850 400371 41853
rect 400438 41850 400444 41852
rect 247677 41792 247682 41848
rect 90100 41788 90106 41790
rect 247677 41788 247724 41792
rect 247788 41790 247834 41850
rect 400305 41848 400444 41850
rect 400305 41792 400310 41848
rect 400366 41792 400444 41848
rect 400305 41790 400444 41792
rect 247788 41788 247794 41790
rect 89989 41787 90055 41788
rect 247677 41787 247743 41788
rect 400305 41787 400371 41790
rect 400438 41788 400444 41790
rect 400508 41788 400514 41852
rect 200798 41652 200804 41716
rect 200868 41714 200874 41716
rect 283782 41714 283788 41716
rect 200868 41654 283788 41714
rect 200868 41652 200874 41654
rect 283782 41652 283788 41654
rect 283852 41652 283858 41716
rect 55070 41516 55076 41580
rect 55140 41578 55146 41580
rect 130878 41578 130884 41580
rect 55140 41518 130884 41578
rect 55140 41516 55146 41518
rect 130878 41516 130884 41518
rect 130948 41516 130954 41580
rect 378910 41516 378916 41580
rect 378980 41578 378986 41580
rect 475878 41578 475884 41580
rect 378980 41518 475884 41578
rect 378980 41516 378986 41518
rect 475878 41516 475884 41518
rect 475948 41516 475954 41580
rect 163262 41380 163268 41444
rect 163332 41380 163338 41444
rect 418470 41380 418476 41444
rect 418540 41380 418546 41444
rect 438342 41380 438348 41444
rect 438412 41380 438418 41444
rect 50654 41244 50660 41308
rect 50724 41306 50730 41308
rect 163270 41306 163330 41380
rect 50724 41246 163330 41306
rect 50724 41244 50730 41246
rect 219934 41244 219940 41308
rect 220004 41306 220010 41308
rect 418478 41306 418538 41380
rect 220004 41246 418538 41306
rect 220004 41244 220010 41246
rect 377806 41108 377812 41172
rect 377876 41170 377882 41172
rect 438350 41170 438410 41380
rect 377876 41110 438410 41170
rect 377876 41108 377882 41110
rect 377254 40972 377260 41036
rect 377324 41034 377330 41036
rect 433333 41034 433399 41037
rect 377324 41032 433399 41034
rect 377324 40976 433338 41032
rect 433394 40976 433399 41032
rect 377324 40974 433399 40976
rect 377324 40972 377330 40974
rect 433333 40971 433399 40974
rect 379462 40836 379468 40900
rect 379532 40898 379538 40900
rect 428549 40898 428615 40901
rect 379532 40896 428615 40898
rect 379532 40840 428554 40896
rect 428610 40840 428615 40896
rect 379532 40838 428615 40840
rect 379532 40836 379538 40838
rect 428549 40835 428615 40838
rect 53414 39884 53420 39948
rect 53484 39946 53490 39948
rect 165797 39946 165863 39949
rect 53484 39944 165863 39946
rect 53484 39888 165802 39944
rect 165858 39888 165863 39944
rect 53484 39886 165863 39888
rect 53484 39884 53490 39886
rect 165797 39883 165863 39886
rect 217542 39884 217548 39948
rect 217612 39946 217618 39948
rect 250069 39946 250135 39949
rect 217612 39944 250135 39946
rect 217612 39888 250074 39944
rect 250130 39888 250135 39944
rect 217612 39886 250135 39888
rect 217612 39884 217618 39886
rect 250069 39883 250135 39886
rect 580441 32058 580507 32061
rect 580901 32058 580967 32061
rect 583520 32058 584960 32148
rect 580441 32056 584960 32058
rect 580441 32000 580446 32056
rect 580502 32000 580906 32056
rect 580962 32000 584960 32056
rect 580441 31998 584960 32000
rect 580441 31995 580507 31998
rect 580901 31995 580967 31998
rect 583520 31908 584960 31998
rect -960 31378 480 31468
rect 2773 31378 2839 31381
rect -960 31376 2839 31378
rect -960 31320 2778 31376
rect 2834 31320 2839 31376
rect -960 31318 2839 31320
rect -960 31228 480 31318
rect 2773 31315 2839 31318
rect 583520 19124 584960 19364
rect -960 18716 480 18956
rect -960 6204 480 6444
rect 583520 6340 584960 6580
<< via3 >>
rect 53052 646172 53116 646236
rect 51580 646036 51644 646100
rect 54340 645900 54404 645964
rect 430620 622100 430684 622164
rect 430804 607820 430868 607884
rect 430620 535468 430684 535532
rect 430804 535332 430868 535396
rect 59308 492492 59372 492556
rect 196572 492492 196636 492556
rect 213316 492492 213380 492556
rect 217364 492492 217428 492556
rect 219940 492492 220004 492556
rect 357940 492492 358004 492556
rect 197860 492356 197924 492420
rect 217548 492356 217612 492420
rect 360700 492356 360764 492420
rect 46796 492220 46860 492284
rect 201356 492220 201420 492284
rect 202644 492220 202708 492284
rect 364932 492220 364996 492284
rect 53604 492084 53668 492148
rect 50844 491948 50908 492012
rect 201172 492084 201236 492148
rect 206876 492084 206940 492148
rect 367692 492084 367756 492148
rect 204852 491948 204916 492012
rect 371740 491948 371804 492012
rect 46612 491812 46676 491876
rect 205036 491812 205100 491876
rect 219204 491812 219268 491876
rect 374500 491812 374564 491876
rect 59124 491676 59188 491740
rect 196756 491676 196820 491740
rect 198044 491676 198108 491740
rect 205220 491676 205284 491740
rect 55076 491540 55140 491604
rect 198412 491540 198476 491604
rect 211660 491540 211724 491604
rect 200620 491404 200684 491468
rect 50292 491268 50356 491332
rect 52316 491328 52380 491332
rect 52316 491272 52366 491328
rect 52366 491272 52380 491328
rect 52316 491268 52380 491272
rect 198596 491268 198660 491332
rect 213868 490452 213932 490516
rect 57100 489636 57164 489700
rect 206508 489092 206572 489156
rect 199148 487732 199212 487796
rect 378180 487732 378244 487796
rect 47716 486916 47780 486980
rect 210372 486508 210436 486572
rect 208900 486372 208964 486436
rect 47900 483924 47964 483988
rect 44956 483788 45020 483852
rect 44772 483652 44836 483716
rect 206140 483652 206204 483716
rect 374684 483652 374748 483716
rect 200804 479436 200868 479500
rect 378732 479436 378796 479500
rect 217180 478212 217244 478276
rect 206324 478076 206388 478140
rect 370452 478076 370516 478140
rect 208348 476716 208412 476780
rect 359780 476716 359844 476780
rect 219020 475492 219084 475556
rect 214420 475356 214484 475420
rect 375972 475356 376036 475420
rect 208532 473996 208596 474060
rect 377260 473996 377324 474060
rect 207980 472500 208044 472564
rect 376156 472500 376220 472564
rect 359964 471140 360028 471204
rect 214604 469916 214668 469980
rect 215340 469780 215404 469844
rect 212580 468420 212644 468484
rect 363460 467196 363524 467260
rect 202276 467060 202340 467124
rect 378916 467060 378980 467124
rect 48084 465700 48148 465764
rect 359412 465700 359476 465764
rect 58940 463388 59004 463452
rect 199332 463388 199396 463452
rect 46428 463252 46492 463316
rect 53420 463116 53484 463180
rect 202092 463116 202156 463180
rect 216076 462980 216140 463044
rect 376708 462980 376772 463044
rect 198780 462844 198844 462908
rect 359596 462844 359660 462908
rect 179644 462164 179708 462228
rect 510844 462164 510908 462228
rect 202460 461620 202524 461684
rect 60228 461484 60292 461548
rect 203196 461484 203260 461548
rect 178356 461408 178420 461412
rect 178356 461352 178370 461408
rect 178370 461352 178420 461408
rect 178356 461348 178420 461352
rect 198964 461348 199028 461412
rect 339724 461272 339788 461276
rect 339724 461216 339738 461272
rect 339738 461216 339788 461272
rect 339724 461212 339788 461216
rect 190868 461000 190932 461004
rect 190868 460944 190918 461000
rect 190918 460944 190932 461000
rect 190868 460940 190932 460944
rect 338252 461000 338316 461004
rect 338252 460944 338302 461000
rect 338302 460944 338316 461000
rect 338252 460940 338316 460944
rect 350948 461000 351012 461004
rect 350948 460944 350998 461000
rect 350998 460944 351012 461000
rect 350948 460940 351012 460944
rect 498516 461000 498580 461004
rect 498516 460944 498530 461000
rect 498530 460944 498580 461000
rect 498516 460940 498580 460944
rect 499804 461000 499868 461004
rect 499804 460944 499854 461000
rect 499854 460944 499868 461000
rect 499804 460940 499868 460944
rect 58756 460804 58820 460868
rect 54892 460668 54956 460732
rect 50476 460532 50540 460596
rect 55628 460396 55692 460460
rect 203012 460396 203076 460460
rect 54708 460260 54772 460324
rect 209820 460260 209884 460324
rect 52132 460124 52196 460188
rect 218652 460124 218716 460188
rect 376892 460124 376956 460188
rect 58572 459988 58636 460052
rect 48636 459580 48700 459644
rect 50660 459580 50724 459644
rect 51764 459580 51828 459644
rect 53236 459580 53300 459644
rect 55444 459640 55508 459644
rect 55444 459584 55494 459640
rect 55494 459584 55508 459640
rect 55444 459580 55508 459584
rect 216996 459580 217060 459644
rect 205404 459308 205468 459372
rect 208164 459172 208228 459236
rect 57468 459036 57532 459100
rect 57836 458900 57900 458964
rect 213132 458900 213196 458964
rect 57652 458764 57716 458828
rect 215892 458764 215956 458828
rect 199148 388452 199212 388516
rect 199516 388452 199580 388516
rect 48636 380972 48700 381036
rect 50292 375260 50356 375324
rect 198044 375260 198108 375324
rect 105492 375048 105556 375052
rect 105492 374992 105506 375048
rect 105506 374992 105556 375048
rect 105492 374988 105556 374992
rect 263732 375048 263796 375052
rect 263732 374992 263746 375048
rect 263746 374992 263796 375048
rect 263732 374988 263796 374992
rect 315252 374988 315316 375052
rect 407804 375048 407868 375052
rect 407804 374992 407818 375048
rect 407818 374992 407868 375048
rect 407804 374988 407868 374992
rect 418292 375048 418356 375052
rect 418292 374992 418306 375048
rect 418306 374992 418356 375048
rect 418292 374988 418356 374992
rect 440372 375048 440436 375052
rect 440372 374992 440386 375048
rect 440386 374992 440436 375048
rect 440372 374988 440436 374992
rect 443132 375048 443196 375052
rect 443132 374992 443146 375048
rect 443146 374992 443196 375048
rect 443132 374988 443196 374992
rect 140926 374912 140990 374916
rect 140926 374856 140962 374912
rect 140962 374856 140990 374912
rect 140926 374852 140990 374856
rect 317828 374716 317892 374780
rect 163366 374640 163430 374644
rect 163366 374584 163410 374640
rect 163410 374584 163430 374640
rect 163366 374580 163430 374584
rect 165950 374640 166014 374644
rect 165950 374584 165986 374640
rect 165986 374584 166014 374640
rect 165950 374580 166014 374584
rect 410742 374640 410806 374644
rect 410742 374584 410762 374640
rect 410762 374584 410806 374640
rect 410742 374580 410806 374584
rect 143510 374504 143574 374508
rect 143510 374448 143538 374504
rect 143538 374448 143574 374504
rect 143510 374444 143574 374448
rect 153438 374504 153502 374508
rect 153438 374448 153474 374504
rect 153474 374448 153502 374504
rect 153438 374444 153502 374448
rect 158484 374504 158548 374508
rect 158484 374448 158534 374504
rect 158534 374448 158548 374504
rect 158484 374444 158548 374448
rect 160918 374504 160982 374508
rect 160918 374448 160926 374504
rect 160926 374448 160982 374504
rect 160918 374444 160982 374448
rect 244228 374504 244292 374508
rect 244228 374448 244278 374504
rect 244278 374448 244292 374504
rect 244228 374444 244292 374448
rect 248702 374504 248766 374508
rect 248702 374448 248750 374504
rect 248750 374448 248766 374504
rect 248702 374444 248766 374448
rect 250062 374504 250126 374508
rect 250062 374448 250074 374504
rect 250074 374448 250126 374504
rect 250062 374444 250126 374448
rect 271142 374504 271206 374508
rect 271142 374448 271198 374504
rect 271198 374448 271206 374504
rect 271142 374444 271206 374448
rect 275766 374444 275830 374508
rect 320918 374504 320982 374508
rect 320918 374448 320970 374504
rect 320970 374448 320982 374504
rect 320918 374444 320982 374448
rect 433318 374504 433382 374508
rect 433318 374448 433338 374504
rect 433338 374448 433382 374504
rect 433318 374444 433382 374448
rect 433590 374504 433654 374508
rect 433590 374448 433614 374504
rect 433614 374448 433654 374504
rect 433590 374444 433654 374448
rect 445966 374504 446030 374508
rect 445966 374448 445998 374504
rect 445998 374448 446030 374504
rect 445966 374444 446030 374448
rect 448278 374504 448342 374508
rect 448278 374448 448298 374504
rect 448298 374448 448342 374504
rect 448278 374444 448342 374448
rect 148916 374368 148980 374372
rect 148916 374312 148966 374368
rect 148966 374312 148980 374368
rect 148916 374308 148980 374312
rect 146156 374232 146220 374236
rect 146156 374176 146206 374232
rect 146206 374176 146220 374232
rect 146156 374172 146220 374176
rect 217548 374172 217612 374236
rect 415716 374232 415780 374236
rect 415716 374176 415730 374232
rect 415730 374176 415780 374232
rect 415716 374172 415780 374176
rect 434852 374232 434916 374236
rect 434852 374176 434866 374232
rect 434866 374176 434916 374232
rect 434852 374172 434916 374176
rect 266308 374036 266372 374100
rect 258028 373960 258092 373964
rect 258028 373904 258078 373960
rect 258078 373904 258092 373960
rect 258028 373900 258092 373904
rect 376892 373900 376956 373964
rect 435220 373900 435284 373964
rect 98132 373764 98196 373828
rect 103284 373764 103348 373828
rect 110460 373824 110524 373828
rect 110460 373768 110474 373824
rect 110474 373768 110524 373824
rect 110460 373764 110524 373768
rect 95004 373688 95068 373692
rect 95004 373632 95054 373688
rect 95054 373632 95068 373688
rect 95004 373628 95068 373632
rect 95924 373628 95988 373692
rect 97580 373628 97644 373692
rect 113588 373688 113652 373692
rect 113588 373632 113602 373688
rect 113602 373632 113652 373688
rect 113588 373628 113652 373632
rect 116164 373688 116228 373692
rect 116164 373632 116178 373688
rect 116178 373632 116228 373688
rect 116164 373628 116228 373632
rect 118372 373688 118436 373692
rect 118372 373632 118386 373688
rect 118386 373632 118436 373688
rect 118372 373628 118436 373632
rect 121316 373688 121380 373692
rect 121316 373632 121366 373688
rect 121366 373632 121380 373688
rect 121316 373628 121380 373632
rect 124076 373688 124140 373692
rect 124076 373632 124126 373688
rect 124126 373632 124140 373688
rect 124076 373628 124140 373632
rect 125732 373688 125796 373692
rect 125732 373632 125746 373688
rect 125746 373632 125796 373688
rect 125732 373628 125796 373632
rect 128860 373688 128924 373692
rect 128860 373632 128910 373688
rect 128910 373632 128924 373688
rect 128860 373628 128924 373632
rect 131068 373688 131132 373692
rect 131068 373632 131082 373688
rect 131082 373632 131132 373688
rect 131068 373628 131132 373632
rect 133644 373688 133708 373692
rect 133644 373632 133694 373688
rect 133694 373632 133708 373688
rect 133644 373628 133708 373632
rect 136404 373688 136468 373692
rect 136404 373632 136454 373688
rect 136454 373632 136468 373688
rect 136404 373628 136468 373632
rect 139164 373688 139228 373692
rect 139164 373632 139214 373688
rect 139214 373632 139228 373688
rect 139164 373628 139228 373632
rect 151676 373688 151740 373692
rect 151676 373632 151726 373688
rect 151726 373632 151740 373688
rect 151676 373628 151740 373632
rect 212764 373764 212828 373828
rect 217364 373764 217428 373828
rect 268516 373764 268580 373828
rect 404860 373824 404924 373828
rect 404860 373768 404874 373824
rect 404874 373768 404924 373824
rect 404860 373764 404924 373768
rect 421052 373824 421116 373828
rect 421052 373768 421066 373824
rect 421066 373768 421116 373824
rect 421052 373764 421116 373768
rect 423076 373824 423140 373828
rect 423076 373768 423090 373824
rect 423090 373768 423140 373824
rect 423076 373764 423140 373768
rect 425468 373824 425532 373828
rect 425468 373768 425482 373824
rect 425482 373768 425532 373824
rect 425468 373764 425532 373768
rect 439452 373824 439516 373828
rect 439452 373768 439466 373824
rect 439466 373768 439516 373824
rect 439452 373764 439516 373768
rect 460980 373824 461044 373828
rect 460980 373768 460994 373824
rect 460994 373768 461044 373824
rect 460980 373764 461044 373768
rect 236500 373688 236564 373692
rect 236500 373632 236514 373688
rect 236514 373632 236564 373688
rect 236500 373628 236564 373632
rect 242940 373688 243004 373692
rect 242940 373632 242954 373688
rect 242954 373632 243004 373688
rect 242940 373628 243004 373632
rect 450308 373688 450372 373692
rect 450308 373632 450322 373688
rect 450322 373632 450372 373688
rect 450308 373628 450372 373632
rect 98316 373552 98380 373556
rect 98316 373496 98330 373552
rect 98330 373496 98380 373552
rect 98316 373492 98380 373496
rect 107884 373552 107948 373556
rect 107884 373496 107898 373552
rect 107898 373496 107948 373552
rect 107884 373492 107948 373496
rect 156460 373552 156524 373556
rect 156460 373496 156510 373552
rect 156510 373496 156524 373552
rect 156460 373492 156524 373496
rect 452884 373552 452948 373556
rect 452884 373496 452898 373552
rect 452898 373496 452948 373552
rect 452884 373492 452948 373496
rect 458220 373552 458284 373556
rect 458220 373496 458234 373552
rect 458234 373496 458284 373552
rect 458220 373492 458284 373496
rect 462820 373552 462884 373556
rect 462820 373496 462834 373552
rect 462834 373496 462884 373552
rect 462820 373492 462884 373496
rect 90220 373416 90284 373420
rect 90220 373360 90234 373416
rect 90234 373360 90284 373416
rect 90220 373356 90284 373360
rect 96108 373416 96172 373420
rect 96108 373360 96122 373416
rect 96122 373360 96172 373416
rect 96108 373356 96172 373360
rect 217364 373356 217428 373420
rect 269252 373416 269316 373420
rect 269252 373360 269266 373416
rect 269266 373360 269316 373416
rect 269252 373356 269316 373360
rect 455460 373416 455524 373420
rect 455460 373360 455474 373416
rect 455474 373360 455524 373416
rect 455460 373356 455524 373360
rect 88380 373280 88444 373284
rect 88380 373224 88394 373280
rect 88394 373224 88444 373280
rect 88380 373220 88444 373224
rect 100892 373280 100956 373284
rect 100892 373224 100906 373280
rect 100906 373224 100956 373280
rect 100892 373220 100956 373224
rect 235948 373220 236012 373284
rect 253980 373280 254044 373284
rect 253980 373224 253994 373280
rect 253994 373224 254044 373280
rect 253980 373220 254044 373224
rect 255452 373280 255516 373284
rect 255452 373224 255466 373280
rect 255466 373224 255516 373280
rect 255452 373220 255516 373224
rect 256740 373280 256804 373284
rect 256740 373224 256754 373280
rect 256754 373224 256804 373280
rect 256740 373220 256804 373224
rect 92428 373144 92492 373148
rect 92428 373088 92442 373144
rect 92442 373088 92492 373144
rect 92428 373084 92492 373088
rect 93716 373144 93780 373148
rect 93716 373088 93730 373144
rect 93730 373088 93780 373144
rect 93716 373084 93780 373088
rect 247172 373144 247236 373148
rect 247172 373088 247186 373144
rect 247186 373088 247236 373144
rect 247172 373084 247236 373088
rect 261340 373144 261404 373148
rect 261340 373088 261354 373144
rect 261354 373088 261404 373144
rect 261340 373084 261404 373088
rect 265020 373144 265084 373148
rect 265020 373088 265034 373144
rect 265034 373088 265084 373144
rect 265020 373084 265084 373088
rect 300900 373144 300964 373148
rect 300900 373088 300914 373144
rect 300914 373088 300964 373144
rect 300900 373084 300964 373088
rect 438164 373144 438228 373148
rect 438164 373088 438214 373144
rect 438214 373088 438228 373144
rect 438164 373084 438228 373088
rect 216628 372812 216692 372876
rect 52132 372676 52196 372740
rect 55444 372676 55508 372740
rect 216812 372676 216876 372740
rect 376708 372676 376772 372740
rect 377996 372736 378060 372740
rect 377996 372680 378046 372736
rect 378046 372680 378060 372736
rect 377996 372676 378060 372680
rect 84700 372600 84764 372604
rect 84700 372544 84750 372600
rect 84750 372544 84764 372600
rect 84700 372540 84764 372544
rect 86724 372600 86788 372604
rect 86724 372544 86774 372600
rect 86774 372544 86788 372600
rect 86724 372540 86788 372544
rect 88012 372600 88076 372604
rect 88012 372544 88062 372600
rect 88062 372544 88076 372600
rect 88012 372540 88076 372544
rect 89300 372600 89364 372604
rect 89300 372544 89350 372600
rect 89350 372544 89364 372600
rect 89300 372540 89364 372544
rect 90036 372540 90100 372604
rect 91508 372600 91572 372604
rect 91508 372544 91558 372600
rect 91558 372544 91572 372600
rect 91508 372540 91572 372544
rect 93348 372600 93412 372604
rect 93348 372544 93398 372600
rect 93398 372544 93412 372600
rect 93348 372540 93412 372544
rect 99972 372600 100036 372604
rect 99972 372544 100022 372600
rect 100022 372544 100036 372600
rect 99972 372540 100036 372544
rect 104572 372600 104636 372604
rect 104572 372544 104622 372600
rect 104622 372544 104636 372600
rect 104572 372540 104636 372544
rect 112852 372540 112916 372604
rect 114508 372600 114572 372604
rect 114508 372544 114522 372600
rect 114522 372544 114572 372600
rect 114508 372540 114572 372544
rect 208348 372540 208412 372604
rect 238156 372600 238220 372604
rect 238156 372544 238170 372600
rect 238170 372544 238220 372600
rect 238156 372540 238220 372544
rect 239076 372600 239140 372604
rect 239076 372544 239126 372600
rect 239126 372544 239140 372600
rect 239076 372540 239140 372544
rect 244780 372540 244844 372604
rect 251956 372540 252020 372604
rect 252876 372540 252940 372604
rect 259500 372600 259564 372604
rect 259500 372544 259514 372600
rect 259514 372544 259564 372600
rect 259500 372540 259564 372544
rect 260052 372540 260116 372604
rect 262260 372600 262324 372604
rect 262260 372544 262274 372600
rect 262274 372544 262324 372600
rect 262260 372540 262324 372544
rect 267044 372540 267108 372604
rect 272564 372540 272628 372604
rect 273852 372540 273916 372604
rect 326660 372540 326724 372604
rect 425284 372540 425348 372604
rect 426388 372600 426452 372604
rect 426388 372544 426438 372600
rect 426438 372544 426452 372600
rect 426388 372540 426452 372544
rect 428596 372540 428660 372604
rect 79916 372404 79980 372468
rect 84516 372464 84580 372468
rect 84516 372408 84566 372464
rect 84566 372408 84580 372464
rect 84516 372404 84580 372408
rect 183140 372404 183204 372468
rect 279004 372404 279068 372468
rect 376708 372404 376772 372468
rect 433564 372404 433628 372468
rect 78260 372328 78324 372332
rect 78260 372272 78310 372328
rect 78310 372272 78324 372328
rect 78260 372268 78324 372272
rect 109540 372268 109604 372332
rect 118188 372268 118252 372332
rect 277532 372268 277596 372332
rect 470732 372268 470796 372332
rect 113220 372132 113284 372196
rect 273300 372132 273364 372196
rect 292804 372132 292868 372196
rect 343220 372192 343284 372196
rect 343220 372136 343234 372192
rect 343234 372136 343284 372192
rect 343220 372132 343284 372136
rect 343404 372192 343468 372196
rect 343404 372136 343454 372192
rect 343454 372136 343468 372192
rect 343404 372132 343468 372136
rect 81940 371996 82004 372060
rect 183324 371920 183388 371924
rect 240548 371996 240612 372060
rect 400260 372132 400324 372196
rect 406148 372132 406212 372196
rect 503116 372192 503180 372196
rect 503116 372136 503166 372192
rect 503166 372136 503180 372192
rect 503116 372132 503180 372136
rect 396212 371996 396276 372060
rect 398972 371996 399036 372060
rect 183324 371864 183338 371920
rect 183338 371864 183388 371920
rect 183324 371860 183388 371864
rect 241652 371860 241716 371924
rect 245884 371860 245948 371924
rect 397500 371920 397564 371924
rect 397500 371864 397514 371920
rect 397514 371864 397564 371920
rect 76604 371724 76668 371788
rect 77156 371784 77220 371788
rect 77156 371728 77206 371784
rect 77206 371728 77220 371784
rect 77156 371724 77220 371728
rect 119844 371724 119908 371788
rect 101996 371648 102060 371652
rect 101996 371592 102046 371648
rect 102046 371592 102060 371648
rect 101996 371588 102060 371592
rect 106964 371648 107028 371652
rect 106964 371592 107014 371648
rect 107014 371592 107028 371648
rect 106964 371588 107028 371592
rect 108804 371648 108868 371652
rect 108804 371592 108854 371648
rect 108854 371592 108868 371648
rect 108804 371588 108868 371592
rect 111564 371648 111628 371652
rect 111564 371592 111614 371648
rect 111614 371592 111628 371648
rect 111564 371588 111628 371592
rect 117084 371588 117148 371652
rect 216996 371588 217060 371652
rect 276428 371724 276492 371788
rect 302924 371724 302988 371788
rect 397500 371860 397564 371864
rect 413692 371860 413756 371924
rect 483244 371860 483308 371924
rect 402284 371724 402348 371788
rect 410012 371724 410076 371788
rect 411852 371724 411916 371788
rect 430620 371784 430684 371788
rect 430620 371728 430634 371784
rect 430634 371728 430684 371784
rect 430620 371724 430684 371728
rect 241652 371588 241716 371652
rect 251220 371648 251284 371652
rect 251220 371592 251234 371648
rect 251234 371592 251284 371648
rect 251220 371588 251284 371592
rect 258396 371588 258460 371652
rect 407252 371588 407316 371652
rect 412772 371588 412836 371652
rect 465396 371588 465460 371652
rect 83780 371512 83844 371516
rect 83780 371456 83830 371512
rect 83830 371456 83844 371512
rect 83780 371452 83844 371456
rect 81020 371316 81084 371380
rect 247908 371452 247972 371516
rect 250300 371452 250364 371516
rect 253612 371452 253676 371516
rect 256188 371452 256252 371516
rect 260972 371452 261036 371516
rect 263548 371512 263612 371516
rect 263548 371456 263598 371512
rect 263598 371456 263612 371512
rect 263548 371452 263612 371456
rect 265756 371452 265820 371516
rect 267780 371512 267844 371516
rect 267780 371456 267794 371512
rect 267794 371456 267844 371512
rect 267780 371452 267844 371456
rect 277532 371452 277596 371516
rect 411300 371512 411364 371516
rect 411300 371456 411314 371512
rect 411314 371456 411364 371512
rect 411300 371452 411364 371456
rect 418844 371452 418908 371516
rect 422340 371512 422404 371516
rect 422340 371456 422354 371512
rect 422354 371456 422404 371512
rect 422340 371452 422404 371456
rect 427676 371452 427740 371516
rect 100708 371316 100772 371380
rect 102732 371376 102796 371380
rect 102732 371320 102782 371376
rect 102782 371320 102796 371376
rect 102732 371316 102796 371320
rect 105308 371316 105372 371380
rect 107516 371316 107580 371380
rect 115796 371316 115860 371380
rect 270908 371316 270972 371380
rect 273668 371316 273732 371380
rect 276244 371316 276308 371380
rect 278268 371316 278332 371380
rect 280292 371316 280356 371380
rect 283788 371316 283852 371380
rect 285812 371316 285876 371380
rect 287652 371316 287716 371380
rect 290596 371316 290660 371380
rect 295380 371376 295444 371380
rect 295380 371320 295394 371376
rect 295394 371320 295444 371376
rect 295380 371316 295444 371320
rect 298140 371376 298204 371380
rect 298140 371320 298154 371376
rect 298154 371320 298204 371376
rect 298140 371316 298204 371320
rect 305316 371316 305380 371380
rect 308628 371316 308692 371380
rect 310652 371316 310716 371380
rect 313412 371316 313476 371380
rect 322980 371376 323044 371380
rect 322980 371320 322994 371376
rect 322994 371320 323044 371376
rect 322980 371316 323044 371320
rect 396580 371316 396644 371380
rect 403020 371376 403084 371380
rect 403020 371320 403034 371376
rect 403034 371320 403084 371376
rect 403020 371316 403084 371320
rect 403572 371316 403636 371380
rect 408540 371376 408604 371380
rect 408540 371320 408554 371376
rect 408554 371320 408604 371376
rect 408540 371316 408604 371320
rect 414060 371376 414124 371380
rect 414060 371320 414074 371376
rect 414074 371320 414124 371376
rect 414060 371316 414124 371320
rect 415532 371316 415596 371380
rect 416820 371376 416884 371380
rect 416820 371320 416834 371376
rect 416834 371320 416884 371376
rect 416820 371316 416884 371320
rect 418108 371376 418172 371380
rect 418108 371320 418158 371376
rect 418158 371320 418172 371376
rect 418108 371316 418172 371320
rect 420316 371316 420380 371380
rect 421236 371316 421300 371380
rect 423996 371316 424060 371380
rect 427860 371376 427924 371380
rect 427860 371320 427874 371376
rect 427874 371320 427924 371376
rect 427860 371316 427924 371320
rect 429332 371316 429396 371380
rect 431172 371316 431236 371380
rect 432092 371316 432156 371380
rect 436324 371316 436388 371380
rect 438348 371316 438412 371380
rect 467972 371316 468036 371380
rect 473308 371376 473372 371380
rect 473308 371320 473358 371376
rect 473358 371320 473372 371376
rect 473308 371316 473372 371320
rect 480300 371376 480364 371380
rect 480300 371320 480314 371376
rect 480314 371320 480364 371376
rect 480300 371316 480364 371320
rect 485820 371376 485884 371380
rect 485820 371320 485834 371376
rect 485834 371320 485884 371376
rect 485820 371316 485884 371320
rect 503484 371316 503548 371380
rect 208532 371180 208596 371244
rect 359964 371180 360028 371244
rect 475332 371180 475396 371244
rect 216812 371044 216876 371108
rect 377260 371044 377324 371108
rect 478092 371044 478156 371108
rect 216628 370500 216692 370564
rect 377812 370364 377876 370428
rect 215340 369820 215404 369884
rect 379468 369820 379532 369884
rect 209820 369140 209884 369204
rect 211660 369140 211724 369204
rect 213316 369140 213380 369204
rect 213868 369140 213932 369204
rect 359780 369004 359844 369068
rect 199516 366284 199580 366348
rect 178540 351868 178604 351932
rect 179644 350568 179708 350572
rect 179644 350512 179694 350568
rect 179694 350512 179708 350568
rect 179644 350508 179708 350512
rect 190868 350508 190932 350572
rect 198964 350508 199028 350572
rect 338436 350568 338500 350572
rect 338436 350512 338486 350568
rect 338486 350512 338500 350568
rect 338436 350508 338500 350512
rect 339724 350508 339788 350572
rect 350948 350508 351012 350572
rect 498516 350508 498580 350572
rect 499804 350508 499868 350572
rect 510844 350568 510908 350572
rect 510844 350512 510894 350568
rect 510894 350512 510908 350568
rect 510844 350508 510908 350512
rect 218836 350372 218900 350436
rect 377260 349692 377324 349756
rect 54340 320180 54404 320244
rect 57100 319908 57164 319972
rect 53052 269180 53116 269244
rect 250484 265024 250548 265028
rect 250484 264968 250498 265024
rect 250498 264968 250548 265024
rect 250484 264964 250548 264968
rect 274220 265024 274284 265028
rect 274220 264968 274234 265024
rect 274234 264968 274284 265024
rect 274220 264964 274284 264968
rect 93462 264828 93526 264892
rect 111006 264888 111070 264892
rect 111006 264832 111026 264888
rect 111026 264832 111070 264888
rect 111006 264828 111070 264832
rect 125966 264888 126030 264892
rect 125966 264832 126022 264888
rect 126022 264832 126030 264888
rect 125966 264828 126030 264832
rect 128308 264888 128372 264892
rect 128308 264832 128358 264888
rect 128358 264832 128372 264888
rect 128308 264828 128372 264832
rect 130998 264828 131062 264892
rect 133446 264888 133510 264892
rect 133446 264832 133474 264888
rect 133474 264832 133510 264888
rect 133446 264828 133510 264832
rect 135894 264888 135958 264892
rect 135894 264832 135902 264888
rect 135902 264832 135958 264888
rect 135894 264828 135958 264832
rect 138478 264888 138542 264892
rect 138478 264832 138534 264888
rect 138534 264832 138542 264888
rect 138478 264828 138542 264832
rect 196756 264828 196820 264892
rect 318470 264828 318534 264892
rect 359412 264828 359476 264892
rect 473438 264888 473502 264892
rect 473438 264832 473450 264888
rect 473450 264832 473502 264888
rect 140926 264692 140990 264756
rect 143510 264752 143574 264756
rect 143510 264696 143538 264752
rect 143538 264696 143574 264752
rect 143510 264692 143574 264696
rect 145958 264752 146022 264756
rect 145958 264696 145986 264752
rect 145986 264696 146022 264752
rect 145958 264692 146022 264696
rect 148542 264752 148606 264756
rect 148542 264696 148562 264752
rect 148562 264696 148606 264752
rect 148542 264692 148606 264696
rect 196572 264692 196636 264756
rect 310990 264692 311054 264756
rect 359596 264692 359660 264756
rect 445966 264692 446030 264756
rect 468542 264692 468606 264756
rect 470990 264752 471054 264756
rect 473438 264828 473502 264832
rect 480918 264888 480982 264892
rect 480918 264832 480958 264888
rect 480958 264832 480982 264888
rect 480918 264828 480982 264832
rect 470990 264696 471022 264752
rect 471022 264696 471054 264752
rect 470990 264692 471054 264696
rect 478470 264692 478534 264756
rect 483366 264752 483430 264756
rect 483366 264696 483386 264752
rect 483386 264696 483430 264752
rect 483366 264692 483430 264696
rect 485950 264752 486014 264756
rect 485950 264696 485962 264752
rect 485962 264696 486014 264752
rect 485950 264692 486014 264696
rect 293446 264616 293510 264620
rect 293446 264560 293462 264616
rect 293462 264560 293510 264616
rect 293446 264556 293510 264560
rect 418494 264556 418558 264620
rect 421078 264616 421142 264620
rect 421078 264560 421102 264616
rect 421102 264560 421142 264616
rect 421078 264556 421142 264560
rect 423526 264616 423590 264620
rect 423526 264560 423550 264616
rect 423550 264560 423590 264616
rect 423526 264556 423590 264560
rect 425974 264616 426038 264620
rect 425974 264560 425978 264616
rect 425978 264560 426034 264616
rect 426034 264560 426038 264616
rect 425974 264556 426038 264560
rect 429782 264616 429846 264620
rect 429782 264560 429806 264616
rect 429806 264560 429846 264616
rect 429782 264556 429846 264560
rect 475886 264616 475950 264620
rect 475886 264560 475898 264616
rect 475898 264560 475950 264616
rect 475886 264556 475950 264560
rect 300900 264420 300964 264484
rect 118004 264148 118068 264212
rect 280844 264344 280908 264348
rect 280844 264288 280858 264344
rect 280858 264288 280908 264344
rect 280844 264284 280908 264288
rect 283420 264344 283484 264348
rect 283420 264288 283434 264344
rect 283434 264288 283484 264344
rect 283420 264284 283484 264288
rect 285996 264344 286060 264348
rect 285996 264288 286010 264344
rect 286010 264288 286060 264344
rect 285996 264284 286060 264288
rect 288204 264344 288268 264348
rect 288204 264288 288218 264344
rect 288218 264288 288268 264344
rect 288204 264284 288268 264288
rect 290964 264344 291028 264348
rect 290964 264288 290978 264344
rect 290978 264288 291028 264344
rect 290964 264284 291028 264288
rect 298508 264284 298572 264348
rect 295932 264148 295996 264212
rect 51764 263604 51828 263668
rect 219020 263604 219084 263668
rect 415900 263664 415964 263668
rect 415900 263608 415914 263664
rect 415914 263608 415964 263664
rect 415900 263604 415964 263608
rect 80468 263468 80532 263532
rect 88380 263528 88444 263532
rect 88380 263472 88394 263528
rect 88394 263472 88444 263528
rect 88380 263468 88444 263472
rect 90036 263528 90100 263532
rect 90036 263472 90050 263528
rect 90050 263472 90100 263528
rect 90036 263468 90100 263472
rect 90772 263528 90836 263532
rect 90772 263472 90786 263528
rect 90786 263472 90836 263528
rect 90772 263468 90836 263472
rect 91324 263528 91388 263532
rect 91324 263472 91338 263528
rect 91338 263472 91388 263528
rect 91324 263468 91388 263472
rect 92428 263528 92492 263532
rect 92428 263472 92442 263528
rect 92442 263472 92492 263528
rect 92428 263468 92492 263472
rect 93716 263468 93780 263532
rect 96108 263528 96172 263532
rect 96108 263472 96122 263528
rect 96122 263472 96172 263528
rect 96108 263468 96172 263472
rect 98500 263468 98564 263532
rect 101076 263528 101140 263532
rect 101076 263472 101090 263528
rect 101090 263472 101140 263528
rect 101076 263468 101140 263472
rect 103284 263468 103348 263532
rect 105860 263468 105924 263532
rect 108252 263528 108316 263532
rect 108252 263472 108266 263528
rect 108266 263472 108316 263528
rect 108252 263468 108316 263472
rect 109724 263468 109788 263532
rect 113588 263468 113652 263532
rect 115980 263528 116044 263532
rect 115980 263472 115994 263528
rect 115994 263472 116044 263528
rect 115980 263468 116044 263472
rect 116900 263468 116964 263532
rect 118372 263468 118436 263532
rect 120948 263528 121012 263532
rect 120948 263472 120962 263528
rect 120962 263472 121012 263528
rect 120948 263468 121012 263472
rect 123524 263528 123588 263532
rect 123524 263472 123538 263528
rect 123538 263472 123588 263528
rect 123524 263468 123588 263472
rect 150940 263528 151004 263532
rect 150940 263472 150990 263528
rect 150990 263472 151004 263528
rect 150940 263468 151004 263472
rect 155908 263528 155972 263532
rect 155908 263472 155958 263528
rect 155958 263472 155972 263528
rect 155908 263468 155972 263472
rect 158484 263528 158548 263532
rect 158484 263472 158534 263528
rect 158534 263472 158548 263528
rect 158484 263468 158548 263472
rect 160876 263468 160940 263532
rect 163452 263528 163516 263532
rect 163452 263472 163502 263528
rect 163502 263472 163516 263528
rect 163452 263468 163516 263472
rect 166028 263528 166092 263532
rect 166028 263472 166078 263528
rect 166078 263472 166092 263528
rect 166028 263468 166092 263472
rect 235948 263528 236012 263532
rect 235948 263472 235998 263528
rect 235998 263472 236012 263528
rect 235948 263468 236012 263472
rect 239628 263468 239692 263532
rect 243124 263528 243188 263532
rect 243124 263472 243138 263528
rect 243138 263472 243188 263528
rect 243124 263468 243188 263472
rect 247540 263468 247604 263532
rect 248276 263468 248340 263532
rect 253612 263528 253676 263532
rect 253612 263472 253626 263528
rect 253626 263472 253676 263528
rect 253612 263468 253676 263472
rect 256188 263528 256252 263532
rect 256188 263472 256202 263528
rect 256202 263472 256252 263528
rect 256188 263468 256252 263472
rect 258212 263528 258276 263532
rect 258212 263472 258226 263528
rect 258226 263472 258276 263528
rect 258212 263468 258276 263472
rect 261708 263468 261772 263532
rect 262812 263468 262876 263532
rect 263548 263528 263612 263532
rect 263548 263472 263598 263528
rect 263598 263472 263612 263528
rect 263548 263468 263612 263472
rect 265204 263468 265268 263532
rect 265940 263528 266004 263532
rect 265940 263472 265954 263528
rect 265954 263472 266004 263528
rect 265940 263468 266004 263472
rect 268332 263528 268396 263532
rect 268332 263472 268346 263528
rect 268346 263472 268396 263528
rect 268332 263468 268396 263472
rect 269804 263528 269868 263532
rect 269804 263472 269818 263528
rect 269818 263472 269868 263528
rect 269804 263468 269868 263472
rect 270908 263528 270972 263532
rect 270908 263472 270922 263528
rect 270922 263472 270972 263528
rect 270908 263468 270972 263472
rect 271276 263528 271340 263532
rect 271276 263472 271290 263528
rect 271290 263472 271340 263528
rect 271276 263468 271340 263472
rect 272196 263468 272260 263532
rect 273300 263528 273364 263532
rect 273300 263472 273314 263528
rect 273314 263472 273364 263528
rect 273300 263468 273364 263472
rect 275876 263528 275940 263532
rect 275876 263472 275926 263528
rect 275926 263472 275940 263528
rect 275876 263468 275940 263472
rect 276060 263528 276124 263532
rect 276060 263472 276110 263528
rect 276110 263472 276124 263528
rect 276060 263468 276124 263472
rect 279188 263528 279252 263532
rect 279188 263472 279238 263528
rect 279238 263472 279252 263528
rect 279188 263468 279252 263472
rect 305868 263528 305932 263532
rect 305868 263472 305882 263528
rect 305882 263472 305932 263528
rect 305868 263468 305932 263472
rect 308444 263528 308508 263532
rect 308444 263472 308458 263528
rect 308458 263472 308508 263528
rect 308444 263468 308508 263472
rect 323348 263468 323412 263532
rect 325924 263468 325988 263532
rect 343220 263468 343284 263532
rect 398236 263468 398300 263532
rect 401732 263468 401796 263532
rect 405412 263468 405476 263532
rect 408356 263528 408420 263532
rect 408356 263472 408370 263528
rect 408370 263472 408420 263528
rect 408356 263468 408420 263472
rect 410748 263528 410812 263532
rect 410748 263472 410762 263528
rect 410762 263472 410812 263528
rect 410748 263468 410812 263472
rect 413692 263528 413756 263532
rect 413692 263472 413706 263528
rect 413706 263472 413756 263528
rect 413692 263468 413756 263472
rect 416084 263468 416148 263532
rect 419396 263528 419460 263532
rect 419396 263472 419410 263528
rect 419410 263472 419460 263528
rect 419396 263468 419460 263472
rect 425284 263528 425348 263532
rect 425284 263472 425298 263528
rect 425298 263472 425348 263528
rect 425284 263468 425348 263472
rect 426388 263528 426452 263532
rect 426388 263472 426438 263528
rect 426438 263472 426452 263528
rect 426388 263468 426452 263472
rect 427492 263528 427556 263532
rect 427492 263472 427506 263528
rect 427506 263472 427556 263528
rect 427492 263468 427556 263472
rect 428228 263528 428292 263532
rect 428228 263472 428242 263528
rect 428242 263472 428292 263528
rect 428228 263468 428292 263472
rect 430988 263528 431052 263532
rect 430988 263472 431002 263528
rect 431002 263472 431052 263528
rect 430988 263468 431052 263472
rect 432276 263528 432340 263532
rect 432276 263472 432290 263528
rect 432290 263472 432340 263528
rect 432276 263468 432340 263472
rect 433380 263528 433444 263532
rect 433380 263472 433394 263528
rect 433394 263472 433444 263528
rect 433380 263468 433444 263472
rect 434484 263468 434548 263532
rect 435956 263528 436020 263532
rect 435956 263472 435970 263528
rect 435970 263472 436020 263528
rect 435956 263468 436020 263472
rect 438164 263468 438228 263532
rect 440924 263528 440988 263532
rect 440924 263472 440938 263528
rect 440938 263472 440988 263528
rect 440924 263468 440988 263472
rect 443500 263528 443564 263532
rect 443500 263472 443514 263528
rect 443514 263472 443564 263528
rect 443500 263468 443564 263472
rect 448284 263528 448348 263532
rect 448284 263472 448298 263528
rect 448298 263472 448348 263528
rect 448284 263468 448348 263472
rect 451044 263528 451108 263532
rect 451044 263472 451058 263528
rect 451058 263472 451108 263528
rect 451044 263468 451108 263472
rect 453436 263528 453500 263532
rect 453436 263472 453450 263528
rect 453450 263472 453500 263528
rect 453436 263468 453500 263472
rect 455828 263528 455892 263532
rect 455828 263472 455842 263528
rect 455842 263472 455892 263528
rect 455828 263468 455892 263472
rect 503484 263528 503548 263532
rect 503484 263472 503534 263528
rect 503534 263472 503548 263528
rect 503484 263468 503548 263472
rect 83044 263332 83108 263396
rect 113404 263332 113468 263396
rect 153516 263332 153580 263396
rect 198780 263332 198844 263396
rect 320956 263332 321020 263396
rect 463556 263332 463620 263396
rect 77156 263196 77220 263260
rect 81756 263196 81820 263260
rect 85436 263196 85500 263260
rect 95924 263196 95988 263260
rect 99420 263256 99484 263260
rect 99420 263200 99470 263256
rect 99470 263200 99484 263256
rect 99420 263196 99484 263200
rect 313412 263196 313476 263260
rect 315804 263196 315868 263260
rect 76052 263060 76116 263124
rect 103836 263060 103900 263124
rect 217180 263060 217244 263124
rect 278452 263060 278516 263124
rect 465948 263196 466012 263260
rect 83964 262924 84028 262988
rect 87644 262984 87708 262988
rect 87644 262928 87658 262984
rect 87658 262928 87708 262984
rect 87644 262924 87708 262928
rect 88748 262924 88812 262988
rect 100708 262984 100772 262988
rect 100708 262928 100758 262984
rect 100758 262928 100772 262984
rect 100708 262924 100772 262928
rect 119108 262924 119172 262988
rect 237052 262924 237116 262988
rect 244228 262924 244292 262988
rect 258396 262984 258460 262988
rect 258396 262928 258410 262984
rect 258410 262928 258460 262984
rect 258396 262924 258460 262928
rect 260972 262984 261036 262988
rect 260972 262928 260986 262984
rect 260986 262928 261036 262984
rect 260972 262924 261036 262928
rect 273484 262924 273548 262988
rect 79548 262788 79612 262852
rect 112116 262788 112180 262852
rect 94452 262652 94516 262716
rect 101812 262712 101876 262716
rect 101812 262656 101826 262712
rect 101826 262656 101876 262712
rect 101812 262652 101876 262656
rect 102732 262652 102796 262716
rect 105308 262652 105372 262716
rect 108620 262652 108684 262716
rect 343404 263060 343468 263124
rect 460980 263060 461044 263124
rect 378180 262924 378244 262988
rect 420684 262924 420748 262988
rect 421788 262984 421852 262988
rect 421788 262928 421802 262984
rect 421802 262928 421852 262984
rect 421788 262924 421852 262928
rect 433564 262984 433628 262988
rect 433564 262928 433578 262984
rect 433578 262928 433628 262984
rect 433564 262924 433628 262928
rect 435772 262924 435836 262988
rect 438532 262924 438596 262988
rect 397132 262788 397196 262852
rect 413324 262788 413388 262852
rect 418108 262848 418172 262852
rect 418108 262792 418158 262848
rect 418158 262792 418172 262848
rect 418108 262788 418172 262792
rect 458404 262652 458468 262716
rect 86540 262516 86604 262580
rect 115796 262516 115860 262580
rect 423996 262576 424060 262580
rect 423996 262520 424010 262576
rect 424010 262520 424060 262576
rect 423996 262516 424060 262520
rect 106412 262380 106476 262444
rect 183140 262380 183204 262444
rect 252324 262380 252388 262444
rect 260604 262380 260668 262444
rect 267596 262380 267660 262444
rect 404124 262380 404188 262444
rect 412404 262380 412468 262444
rect 78260 262244 78324 262308
rect 97028 262244 97092 262308
rect 98132 262244 98196 262308
rect 107516 262304 107580 262308
rect 107516 262248 107566 262304
rect 107566 262248 107580 262304
rect 107516 262244 107580 262248
rect 111196 262244 111260 262308
rect 114324 262244 114388 262308
rect 183508 262244 183572 262308
rect 238156 262244 238220 262308
rect 240548 262244 240612 262308
rect 241652 262244 241716 262308
rect 245332 262244 245396 262308
rect 246436 262244 246500 262308
rect 248644 262244 248708 262308
rect 250116 262244 250180 262308
rect 251220 262304 251284 262308
rect 251220 262248 251270 262304
rect 251270 262248 251284 262304
rect 251220 262244 251284 262248
rect 253428 262244 253492 262308
rect 254532 262244 254596 262308
rect 255820 262244 255884 262308
rect 256924 262244 256988 262308
rect 259500 262304 259564 262308
rect 259500 262248 259514 262304
rect 259514 262248 259564 262304
rect 259500 262244 259564 262248
rect 263916 262244 263980 262308
rect 266308 262244 266372 262308
rect 268700 262244 268764 262308
rect 276980 262244 277044 262308
rect 278084 262244 278148 262308
rect 303476 262244 303540 262308
rect 396028 262244 396092 262308
rect 199332 262108 199396 262172
rect 399524 262244 399588 262308
rect 400444 262244 400508 262308
rect 403020 262304 403084 262308
rect 403020 262248 403034 262304
rect 403034 262248 403084 262304
rect 403020 262244 403084 262248
rect 406516 262244 406580 262308
rect 407620 262244 407684 262308
rect 408724 262244 408788 262308
rect 410012 262244 410076 262308
rect 411300 262304 411364 262308
rect 411300 262248 411350 262304
rect 411350 262248 411364 262304
rect 411300 262244 411364 262248
rect 414612 262244 414676 262308
rect 417004 262244 417068 262308
rect 422892 262244 422956 262308
rect 428596 262244 428660 262308
rect 431172 262244 431236 262308
rect 436876 262244 436940 262308
rect 439268 262244 439332 262308
rect 503116 262244 503180 262308
rect 377996 260884 378060 260948
rect 47716 260748 47780 260812
rect 44956 260340 45020 260404
rect 44772 260068 44836 260132
rect 377812 260068 377876 260132
rect 510844 241436 510908 241500
rect 178540 240212 178604 240276
rect 179644 240212 179708 240276
rect 190868 240272 190932 240276
rect 190868 240216 190918 240272
rect 190918 240216 190932 240272
rect 190868 240212 190932 240216
rect 217548 240212 217612 240276
rect 338436 240212 338500 240276
rect 339724 240212 339788 240276
rect 350948 240212 351012 240276
rect 379652 240212 379716 240276
rect 498516 240212 498580 240276
rect 499804 240212 499868 240276
rect 377260 239804 377324 239868
rect 379652 239592 379716 239596
rect 379652 239536 379702 239592
rect 379702 239536 379716 239592
rect 379652 239532 379716 239536
rect 377996 239396 378060 239460
rect 47900 238580 47964 238644
rect 57100 237416 57164 237420
rect 57100 237360 57150 237416
rect 57150 237360 57164 237416
rect 57100 237356 57164 237360
rect 51580 219404 51644 219468
rect 57468 162964 57532 163028
rect 96046 154728 96110 154732
rect 96046 154672 96066 154728
rect 96066 154672 96110 154728
rect 96046 154668 96110 154672
rect 113318 154728 113382 154732
rect 113318 154672 113362 154728
rect 113362 154672 113382 154728
rect 113318 154668 113382 154672
rect 163366 154728 163430 154732
rect 163366 154672 163374 154728
rect 163374 154672 163430 154728
rect 163366 154668 163430 154672
rect 165950 154668 166014 154732
rect 261078 154532 261142 154596
rect 273590 154532 273654 154596
rect 57652 154396 57716 154460
rect 148548 154396 148612 154460
rect 202460 154396 202524 154460
rect 315804 154396 315868 154460
rect 418476 154456 418540 154460
rect 418476 154400 418490 154456
rect 418490 154400 418540 154456
rect 418476 154396 418540 154400
rect 421052 154456 421116 154460
rect 421052 154400 421066 154456
rect 421066 154400 421116 154456
rect 421052 154396 421116 154400
rect 426020 154456 426084 154460
rect 426020 154400 426034 154456
rect 426034 154400 426084 154456
rect 426020 154396 426084 154400
rect 443500 154456 443564 154460
rect 443500 154400 443514 154456
rect 443514 154400 443564 154456
rect 443500 154396 443564 154400
rect 57836 154260 57900 154324
rect 138428 154320 138492 154324
rect 138428 154264 138442 154320
rect 138442 154264 138492 154320
rect 98500 154184 98564 154188
rect 98500 154128 98514 154184
rect 98514 154128 98564 154184
rect 98500 154124 98564 154128
rect 101076 154184 101140 154188
rect 101076 154128 101090 154184
rect 101090 154128 101140 154184
rect 101076 154124 101140 154128
rect 105860 154184 105924 154188
rect 105860 154128 105874 154184
rect 105874 154128 105924 154184
rect 105860 154124 105924 154128
rect 108252 154184 108316 154188
rect 108252 154128 108266 154184
rect 108266 154128 108316 154184
rect 108252 154124 108316 154128
rect 138428 154260 138492 154264
rect 208164 154260 208228 154324
rect 313412 154260 313476 154324
rect 475884 154320 475948 154324
rect 475884 154264 475898 154320
rect 475898 154264 475948 154320
rect 475884 154260 475948 154264
rect 478460 154320 478524 154324
rect 478460 154264 478474 154320
rect 478474 154264 478524 154320
rect 478460 154260 478524 154264
rect 140820 154124 140884 154188
rect 143580 154184 143644 154188
rect 143580 154128 143594 154184
rect 143594 154128 143644 154184
rect 143580 154124 143644 154128
rect 203012 154124 203076 154188
rect 288204 154184 288268 154188
rect 288204 154128 288218 154184
rect 288218 154128 288268 154184
rect 288204 154124 288268 154128
rect 293356 154184 293420 154188
rect 293356 154128 293370 154184
rect 293370 154128 293420 154184
rect 293356 154124 293420 154128
rect 145972 154048 146036 154052
rect 145972 153992 145986 154048
rect 145986 153992 146036 154048
rect 145972 153988 146036 153992
rect 150940 154048 151004 154052
rect 150940 153992 150954 154048
rect 150954 153992 151004 154048
rect 150940 153988 151004 153992
rect 216076 153988 216140 154052
rect 305868 154124 305932 154188
rect 473492 154184 473556 154188
rect 473492 154128 473506 154184
rect 473506 154128 473556 154184
rect 473492 154124 473556 154128
rect 480852 154184 480916 154188
rect 480852 154128 480866 154184
rect 480866 154128 480916 154184
rect 480852 154124 480916 154128
rect 298508 154048 298572 154052
rect 298508 153992 298522 154048
rect 298522 153992 298572 154048
rect 298508 153988 298572 153992
rect 303476 154048 303540 154052
rect 303476 153992 303490 154048
rect 303490 153992 303540 154048
rect 303476 153988 303540 153992
rect 470916 154048 470980 154052
rect 470916 153992 470930 154048
rect 470930 153992 470980 154048
rect 470916 153988 470980 153992
rect 483244 154048 483308 154052
rect 483244 153992 483258 154048
rect 483258 153992 483308 154048
rect 483244 153988 483308 153992
rect 153332 153912 153396 153916
rect 153332 153856 153346 153912
rect 153346 153856 153396 153912
rect 153332 153852 153396 153856
rect 213132 153852 213196 153916
rect 270908 153852 270972 153916
rect 295932 153852 295996 153916
rect 308444 153912 308508 153916
rect 308444 153856 308458 153912
rect 308458 153856 308508 153912
rect 308444 153852 308508 153856
rect 423444 153912 423508 153916
rect 423444 153856 423458 153912
rect 423458 153856 423508 153912
rect 423444 153852 423508 153856
rect 486004 153912 486068 153916
rect 486004 153856 486018 153912
rect 486018 153856 486068 153912
rect 486004 153852 486068 153856
rect 85436 153172 85500 153236
rect 95924 153172 95988 153236
rect 99420 153172 99484 153236
rect 236132 153172 236196 153236
rect 261708 153172 261772 153236
rect 265204 153172 265268 153236
rect 272196 153172 272260 153236
rect 300900 153172 300964 153236
rect 398236 153172 398300 153236
rect 401732 153172 401796 153236
rect 416084 153172 416148 153236
rect 455828 153172 455892 153236
rect 463556 153172 463620 153236
rect 76052 153036 76116 153100
rect 78260 153036 78324 153100
rect 79548 153036 79612 153100
rect 81940 153036 82004 153100
rect 83044 153036 83108 153100
rect 86540 153036 86604 153100
rect 87644 153036 87708 153100
rect 88748 153036 88812 153100
rect 90036 153036 90100 153100
rect 91324 153036 91388 153100
rect 93348 153036 93412 153100
rect 94452 153036 94516 153100
rect 97028 153036 97092 153100
rect 98132 153036 98196 153100
rect 100708 153036 100772 153100
rect 102732 153036 102796 153100
rect 103836 153036 103900 153100
rect 106412 153096 106476 153100
rect 106412 153040 106426 153096
rect 106426 153040 106476 153096
rect 106412 153036 106476 153040
rect 108804 153036 108868 153100
rect 111012 153036 111076 153100
rect 111196 153096 111260 153100
rect 111196 153040 111210 153096
rect 111210 153040 111260 153096
rect 111196 153036 111260 153040
rect 112116 153036 112180 153100
rect 114508 153096 114572 153100
rect 114508 153040 114558 153096
rect 114558 153040 114572 153096
rect 114508 153036 114572 153040
rect 115796 153036 115860 153100
rect 117084 153036 117148 153100
rect 118372 153036 118436 153100
rect 119108 153036 119172 153100
rect 125916 153036 125980 153100
rect 128492 153036 128556 153100
rect 130884 153036 130948 153100
rect 133460 153036 133524 153100
rect 136036 153036 136100 153100
rect 155908 153096 155972 153100
rect 155908 153040 155958 153096
rect 155958 153040 155972 153096
rect 155908 153036 155972 153040
rect 218652 153036 218716 153100
rect 238156 153036 238220 153100
rect 240548 153036 240612 153100
rect 241652 153036 241716 153100
rect 242940 153096 243004 153100
rect 242940 153040 242954 153096
rect 242954 153040 243004 153096
rect 242940 153036 243004 153040
rect 244228 153096 244292 153100
rect 244228 153040 244278 153096
rect 244278 153040 244292 153096
rect 244228 153036 244292 153040
rect 246436 153036 246500 153100
rect 247724 153036 247788 153100
rect 248644 153036 248708 153100
rect 250116 153036 250180 153100
rect 250668 153036 250732 153100
rect 251220 153096 251284 153100
rect 251220 153040 251234 153096
rect 251234 153040 251284 153096
rect 251220 153036 251284 153040
rect 253428 153036 253492 153100
rect 253612 153096 253676 153100
rect 253612 153040 253626 153096
rect 253626 153040 253676 153096
rect 253612 153036 253676 153040
rect 254532 153036 254596 153100
rect 255820 153036 255884 153100
rect 256188 153036 256252 153100
rect 256924 153036 256988 153100
rect 258212 153036 258276 153100
rect 259500 153096 259564 153100
rect 259500 153040 259550 153096
rect 259550 153040 259564 153096
rect 259500 153036 259564 153040
rect 262812 153036 262876 153100
rect 263916 153036 263980 153100
rect 266308 153096 266372 153100
rect 266308 153040 266358 153096
rect 266358 153040 266372 153096
rect 266308 153036 266372 153040
rect 268700 153036 268764 153100
rect 269804 153036 269868 153100
rect 271092 153036 271156 153100
rect 274404 153036 274468 153100
rect 275324 153036 275388 153100
rect 278452 153036 278516 153100
rect 279004 153036 279068 153100
rect 280844 153036 280908 153100
rect 283788 153036 283852 153100
rect 285996 153036 286060 153100
rect 290964 153036 291028 153100
rect 320956 153036 321020 153100
rect 396028 153096 396092 153100
rect 396028 153040 396078 153096
rect 396078 153040 396092 153096
rect 396028 153036 396092 153040
rect 399524 153036 399588 153100
rect 400444 153036 400508 153100
rect 403020 153096 403084 153100
rect 403020 153040 403070 153096
rect 403070 153040 403084 153096
rect 403020 153036 403084 153040
rect 405044 153036 405108 153100
rect 406516 153036 406580 153100
rect 407620 153036 407684 153100
rect 408724 153036 408788 153100
rect 410012 153096 410076 153100
rect 410012 153040 410026 153096
rect 410026 153040 410076 153096
rect 410012 153036 410076 153040
rect 411300 153096 411364 153100
rect 411300 153040 411350 153096
rect 411350 153040 411364 153096
rect 411300 153036 411364 153040
rect 413508 153036 413572 153100
rect 414428 153036 414492 153100
rect 415532 153096 415596 153100
rect 415532 153040 415546 153096
rect 415546 153040 415596 153096
rect 415532 153036 415596 153040
rect 417004 153036 417068 153100
rect 418108 153036 418172 153100
rect 420684 153036 420748 153100
rect 421788 153036 421852 153100
rect 422892 153036 422956 153100
rect 423996 153036 424060 153100
rect 425284 153036 425348 153100
rect 426388 153036 426452 153100
rect 428596 153036 428660 153100
rect 429700 153036 429764 153100
rect 431172 153036 431236 153100
rect 431724 153036 431788 153100
rect 433564 153036 433628 153100
rect 434668 153036 434732 153100
rect 435956 153036 436020 153100
rect 436876 153036 436940 153100
rect 438348 153036 438412 153100
rect 439268 153036 439332 153100
rect 440924 153036 440988 153100
rect 445892 153036 445956 153100
rect 448284 153036 448348 153100
rect 451044 153036 451108 153100
rect 453436 153036 453500 153100
rect 458404 153036 458468 153100
rect 158484 152900 158548 152964
rect 206508 152900 206572 152964
rect 318380 152900 318444 152964
rect 48084 152764 48148 152828
rect 91508 152764 91572 152828
rect 101812 152764 101876 152828
rect 103836 152764 103900 152828
rect 107516 152764 107580 152828
rect 109540 152764 109604 152828
rect 113220 152824 113284 152828
rect 113220 152768 113234 152824
rect 113234 152768 113284 152824
rect 113220 152764 113284 152768
rect 118004 152764 118068 152828
rect 120764 152764 120828 152828
rect 122604 152764 122668 152828
rect 183140 152764 183204 152828
rect 311020 152764 311084 152828
rect 343220 152764 343284 152828
rect 468524 152764 468588 152828
rect 160876 152628 160940 152692
rect 214604 152628 214668 152692
rect 77156 152492 77220 152556
rect 93716 152492 93780 152556
rect 115980 152552 116044 152556
rect 115980 152496 115994 152552
rect 115994 152496 116044 152552
rect 115980 152492 116044 152496
rect 183508 152552 183572 152556
rect 183508 152496 183522 152552
rect 183522 152496 183572 152552
rect 183508 152492 183572 152496
rect 203196 152492 203260 152556
rect 88380 152416 88444 152420
rect 88380 152360 88394 152416
rect 88394 152360 88444 152416
rect 88380 152356 88444 152360
rect 90772 152356 90836 152420
rect 237052 152356 237116 152420
rect 245332 152356 245396 152420
rect 248276 152356 248340 152420
rect 252324 152356 252388 152420
rect 258396 152492 258460 152556
rect 260604 152628 260668 152692
rect 265940 152628 266004 152692
rect 267596 152628 267660 152692
rect 268332 152628 268396 152692
rect 273300 152628 273364 152692
rect 460980 152628 461044 152692
rect 503484 152628 503548 152692
rect 276244 152492 276308 152556
rect 343404 152492 343468 152556
rect 397132 152492 397196 152556
rect 404124 152492 404188 152556
rect 410748 152492 410812 152556
rect 412404 152492 412468 152556
rect 413692 152492 413756 152556
rect 419212 152492 419276 152556
rect 427676 152492 427740 152556
rect 433380 152492 433444 152556
rect 435772 152492 435836 152556
rect 438532 152492 438596 152556
rect 503116 152492 503180 152556
rect 263548 152356 263612 152420
rect 408172 152356 408236 152420
rect 465948 152220 466012 152284
rect 105308 152084 105372 152148
rect 202276 152084 202340 152148
rect 325556 152084 325620 152148
rect 80468 151948 80532 152012
rect 84148 151948 84212 152012
rect 238708 152008 238772 152012
rect 238708 151952 238758 152008
rect 238758 151952 238772 152008
rect 238708 151948 238772 151952
rect 276980 151948 277044 152012
rect 277348 151812 277412 151876
rect 205404 151676 205468 151740
rect 322980 151676 323044 151740
rect 430620 151676 430684 151740
rect 427860 151540 427924 151604
rect 379468 151268 379532 151332
rect 57836 150512 57900 150516
rect 57836 150456 57850 150512
rect 57850 150456 57900 150512
rect 57836 150452 57900 150456
rect 57100 133724 57164 133788
rect 377260 133724 377324 133788
rect 377812 133044 377876 133108
rect 57100 132364 57164 132428
rect 217548 130868 217612 130932
rect 377996 130868 378060 130932
rect 57284 130324 57348 130388
rect 190868 130324 190932 130388
rect 510844 130324 510908 130388
rect 178540 129780 178604 129844
rect 179644 129780 179708 129844
rect 338436 129840 338500 129844
rect 338436 129784 338486 129840
rect 338486 129784 338500 129840
rect 338436 129780 338500 129784
rect 339724 129780 339788 129844
rect 350948 129780 351012 129844
rect 377996 129780 378060 129844
rect 498516 129780 498580 129844
rect 499804 129780 499868 129844
rect 54708 129644 54772 129708
rect 57284 129508 57348 129572
rect 202092 54980 202156 55044
rect 46612 53892 46676 53956
rect 206324 53076 206388 53140
rect 46796 52668 46860 52732
rect 77142 44840 77206 44844
rect 77142 44784 77170 44840
rect 77170 44784 77206 44840
rect 77142 44780 77206 44784
rect 83126 44840 83190 44844
rect 83126 44784 83150 44840
rect 83150 44784 83190 44840
rect 83126 44780 83190 44784
rect 84214 44840 84278 44844
rect 84214 44784 84254 44840
rect 84254 44784 84278 44840
rect 84214 44780 84278 44784
rect 94550 44840 94614 44844
rect 94550 44784 94558 44840
rect 94558 44784 94614 44840
rect 94550 44780 94614 44784
rect 96998 44840 97062 44844
rect 96998 44784 97042 44840
rect 97042 44784 97062 44840
rect 96998 44780 97062 44784
rect 98086 44840 98150 44844
rect 98086 44784 98090 44840
rect 98090 44784 98146 44840
rect 98146 44784 98150 44840
rect 98086 44780 98150 44784
rect 218836 44780 218900 44844
rect 219204 44840 219268 44844
rect 219204 44784 219254 44840
rect 219254 44784 219268 44840
rect 219204 44780 219268 44784
rect 236054 44780 236118 44844
rect 237142 44840 237206 44844
rect 237142 44784 237158 44840
rect 237158 44784 237206 44840
rect 237142 44780 237206 44784
rect 243126 44840 243190 44844
rect 243126 44784 243138 44840
rect 243138 44784 243190 44840
rect 243126 44780 243190 44784
rect 244214 44780 244278 44844
rect 396054 44840 396118 44844
rect 396054 44784 396078 44840
rect 396078 44784 396118 44840
rect 396054 44780 396118 44784
rect 397142 44840 397206 44844
rect 397142 44784 397146 44840
rect 397146 44784 397206 44840
rect 397142 44780 397206 44784
rect 403126 44780 403190 44844
rect 414550 44840 414614 44844
rect 414550 44784 414570 44840
rect 414570 44784 414614 44840
rect 414550 44780 414614 44784
rect 416998 44840 417062 44844
rect 416998 44784 417018 44840
rect 417018 44784 417062 44840
rect 416998 44780 417062 44784
rect 57284 44644 57348 44708
rect 99446 44644 99510 44708
rect 100708 44704 100772 44708
rect 100708 44648 100758 44704
rect 100758 44648 100772 44704
rect 100708 44644 100772 44648
rect 101758 44704 101822 44708
rect 101758 44648 101770 44704
rect 101770 44648 101822 44704
rect 101758 44644 101822 44648
rect 102846 44644 102910 44708
rect 103934 44704 103998 44708
rect 103934 44648 103942 44704
rect 103942 44648 103998 44704
rect 103934 44644 103998 44648
rect 143510 44704 143574 44708
rect 143510 44648 143538 44704
rect 143538 44648 143574 44704
rect 143510 44644 143574 44648
rect 145958 44704 146022 44708
rect 145958 44648 145986 44704
rect 145986 44648 146022 44704
rect 145958 44644 146022 44648
rect 205036 44644 205100 44708
rect 250742 44644 250806 44708
rect 255910 44704 255974 44708
rect 255910 44648 255926 44704
rect 255926 44648 255974 44704
rect 255910 44644 255974 44648
rect 256998 44704 257062 44708
rect 256998 44648 257030 44704
rect 257030 44648 257062 44704
rect 256998 44644 257062 44648
rect 258086 44704 258150 44708
rect 258086 44648 258134 44704
rect 258134 44648 258150 44704
rect 258086 44644 258150 44648
rect 262846 44704 262910 44708
rect 262846 44648 262862 44704
rect 262862 44648 262910 44704
rect 262846 44644 262910 44648
rect 315886 44704 315950 44708
rect 315886 44648 315910 44704
rect 315910 44648 315950 44704
rect 315886 44644 315950 44648
rect 410742 44704 410806 44708
rect 410742 44648 410762 44704
rect 410762 44648 410806 44704
rect 410742 44644 410806 44648
rect 419446 44704 419510 44708
rect 419446 44648 419502 44704
rect 419502 44648 419510 44704
rect 419446 44644 419510 44648
rect 423934 44704 423998 44708
rect 423934 44648 423954 44704
rect 423954 44648 423998 44704
rect 423934 44644 423998 44648
rect 50476 44508 50540 44572
rect 108286 44508 108350 44572
rect 113318 44568 113382 44572
rect 113318 44512 113326 44568
rect 113326 44512 113382 44568
rect 113318 44508 113382 44512
rect 140926 44508 140990 44572
rect 205220 44508 205284 44572
rect 258494 44508 258558 44572
rect 259446 44568 259510 44572
rect 259446 44512 259458 44568
rect 259458 44512 259510 44568
rect 259446 44508 259510 44512
rect 55628 44372 55692 44436
rect 138428 44372 138492 44436
rect 260670 44568 260734 44572
rect 260670 44512 260710 44568
rect 260710 44512 260734 44568
rect 260670 44508 260734 44512
rect 261758 44568 261822 44572
rect 261758 44512 261814 44568
rect 261814 44512 261822 44568
rect 261758 44508 261822 44512
rect 263934 44508 263998 44572
rect 305958 44508 306022 44572
rect 308542 44568 308606 44572
rect 308542 44512 308550 44568
rect 308550 44512 308606 44568
rect 308542 44508 308606 44512
rect 404214 44568 404278 44572
rect 404214 44512 404230 44568
rect 404230 44512 404278 44568
rect 404214 44508 404278 44512
rect 405438 44568 405502 44572
rect 405438 44512 405462 44568
rect 405462 44512 405502 44568
rect 405438 44508 405502 44512
rect 53604 44236 53668 44300
rect 201172 44372 201236 44436
rect 406526 44568 406590 44572
rect 406526 44512 406530 44568
rect 406530 44512 406590 44568
rect 406526 44508 406590 44512
rect 418108 44568 418172 44572
rect 418108 44512 418158 44568
rect 418158 44512 418172 44568
rect 418108 44508 418172 44512
rect 420670 44568 420734 44572
rect 420670 44512 420698 44568
rect 420698 44512 420734 44568
rect 420670 44508 420734 44512
rect 421758 44568 421822 44572
rect 421758 44512 421802 44568
rect 421802 44512 421822 44568
rect 421758 44508 421822 44512
rect 422846 44568 422910 44572
rect 422846 44512 422850 44568
rect 422850 44512 422906 44568
rect 422906 44512 422910 44568
rect 422846 44508 422910 44512
rect 423526 44508 423590 44572
rect 425974 44568 426038 44572
rect 425974 44512 425978 44568
rect 425978 44512 426034 44568
rect 426034 44512 426038 44568
rect 425974 44508 426038 44512
rect 439166 44568 439230 44572
rect 439166 44512 439226 44568
rect 439226 44512 439230 44568
rect 439166 44508 439230 44512
rect 455894 44568 455958 44572
rect 455894 44512 455934 44568
rect 455934 44512 455958 44568
rect 455894 44508 455958 44512
rect 458478 44568 458542 44572
rect 458478 44512 458510 44568
rect 458510 44512 458542 44568
rect 458478 44508 458542 44512
rect 480918 44508 480982 44572
rect 425284 44432 425348 44436
rect 425284 44376 425298 44432
rect 425298 44376 425348 44432
rect 425284 44372 425348 44376
rect 198412 44236 198476 44300
rect 323348 44236 323412 44300
rect 360700 44236 360764 44300
rect 53236 44100 53300 44164
rect 153332 44100 153396 44164
rect 158484 44160 158548 44164
rect 158484 44104 158498 44160
rect 158498 44104 158548 44160
rect 158484 44100 158548 44104
rect 160876 44160 160940 44164
rect 160876 44104 160890 44160
rect 160890 44104 160940 44160
rect 160876 44100 160940 44104
rect 206876 44100 206940 44164
rect 295932 44100 295996 44164
rect 300900 44160 300964 44164
rect 300900 44104 300914 44160
rect 300914 44104 300964 44160
rect 300900 44100 300964 44104
rect 357940 44100 358004 44164
rect 483428 44100 483492 44164
rect 52316 43964 52380 44028
rect 150940 43964 151004 44028
rect 202644 43964 202708 44028
rect 290964 43964 291028 44028
rect 364932 43964 364996 44028
rect 478460 43964 478524 44028
rect 50844 43828 50908 43892
rect 148548 43828 148612 43892
rect 198596 43828 198660 43892
rect 279188 43888 279252 43892
rect 279188 43832 279238 43888
rect 279238 43832 279252 43888
rect 46428 43692 46492 43756
rect 111012 43692 111076 43756
rect 115980 43752 116044 43756
rect 115980 43696 115994 43752
rect 115994 43696 116044 43752
rect 115980 43692 116044 43696
rect 197860 43692 197924 43756
rect 278452 43692 278516 43756
rect 279188 43828 279252 43832
rect 367692 43828 367756 43892
rect 468524 43828 468588 43892
rect 285996 43692 286060 43756
rect 374500 43692 374564 43756
rect 473492 43692 473556 43756
rect 59308 43556 59372 43620
rect 123524 43556 123588 43620
rect 201356 43556 201420 43620
rect 280844 43556 280908 43620
rect 371740 43556 371804 43620
rect 57100 43420 57164 43484
rect 105308 43420 105372 43484
rect 204852 43420 204916 43484
rect 273484 43420 273548 43484
rect 407620 43480 407684 43484
rect 407620 43424 407634 43480
rect 407634 43424 407684 43480
rect 407620 43420 407684 43424
rect 421052 43480 421116 43484
rect 421052 43424 421066 43480
rect 421066 43424 421116 43480
rect 421052 43420 421116 43424
rect 428228 43480 428292 43484
rect 428228 43424 428242 43480
rect 428242 43424 428292 43480
rect 428228 43420 428292 43424
rect 463556 43420 463620 43484
rect 59124 43284 59188 43348
rect 101076 43284 101140 43348
rect 200620 43284 200684 43348
rect 265940 43284 266004 43348
rect 85436 43208 85500 43212
rect 85436 43152 85450 43208
rect 85450 43152 85500 43208
rect 85436 43148 85500 43152
rect 92428 43208 92492 43212
rect 92428 43152 92442 43208
rect 92442 43152 92492 43208
rect 92428 43148 92492 43152
rect 95924 43208 95988 43212
rect 95924 43152 95938 43208
rect 95938 43152 95988 43208
rect 95924 43148 95988 43152
rect 128308 43208 128372 43212
rect 128308 43152 128358 43208
rect 128358 43152 128372 43208
rect 128308 43148 128372 43152
rect 265204 43208 265268 43212
rect 265204 43152 265218 43208
rect 265218 43152 265268 43208
rect 265204 43148 265268 43152
rect 272196 43208 272260 43212
rect 272196 43152 272210 43208
rect 272210 43152 272260 43208
rect 272196 43148 272260 43152
rect 325924 43208 325988 43212
rect 325924 43152 325938 43208
rect 325938 43152 325988 43208
rect 325924 43148 325988 43152
rect 398236 43208 398300 43212
rect 398236 43152 398250 43208
rect 398250 43152 398300 43208
rect 398236 43148 398300 43152
rect 401732 43208 401796 43212
rect 401732 43152 401746 43208
rect 401746 43152 401796 43208
rect 401732 43148 401796 43152
rect 76052 42800 76116 42804
rect 76052 42744 76066 42800
rect 76066 42744 76116 42800
rect 76052 42740 76116 42744
rect 78260 42800 78324 42804
rect 78260 42744 78274 42800
rect 78274 42744 78324 42800
rect 78260 42740 78324 42744
rect 80468 42800 80532 42804
rect 80468 42744 80482 42800
rect 80482 42744 80532 42800
rect 80468 42740 80532 42744
rect 86540 42800 86604 42804
rect 86540 42744 86554 42800
rect 86554 42744 86604 42800
rect 86540 42740 86604 42744
rect 87644 42800 87708 42804
rect 87644 42744 87658 42800
rect 87658 42744 87708 42800
rect 87644 42740 87708 42744
rect 88380 42800 88444 42804
rect 88380 42744 88394 42800
rect 88394 42744 88444 42800
rect 88380 42740 88444 42744
rect 88748 42740 88812 42804
rect 90772 42800 90836 42804
rect 90772 42744 90786 42800
rect 90786 42744 90836 42800
rect 90772 42740 90836 42744
rect 91324 42800 91388 42804
rect 91324 42744 91338 42800
rect 91338 42744 91388 42800
rect 91324 42740 91388 42744
rect 93348 42800 93412 42804
rect 93348 42744 93362 42800
rect 93362 42744 93412 42800
rect 93348 42740 93412 42744
rect 93716 42800 93780 42804
rect 93716 42744 93730 42800
rect 93730 42744 93780 42800
rect 93716 42740 93780 42744
rect 96292 42800 96356 42804
rect 96292 42744 96306 42800
rect 96306 42744 96356 42800
rect 96292 42740 96356 42744
rect 106412 42800 106476 42804
rect 106412 42744 106426 42800
rect 106426 42744 106476 42800
rect 106412 42740 106476 42744
rect 107516 42740 107580 42804
rect 108620 42800 108684 42804
rect 108620 42744 108634 42800
rect 108634 42744 108684 42800
rect 108620 42740 108684 42744
rect 112116 42740 112180 42804
rect 113220 42800 113284 42804
rect 113220 42744 113234 42800
rect 113234 42744 113284 42800
rect 113220 42740 113284 42744
rect 114324 42740 114388 42804
rect 115796 42800 115860 42804
rect 115796 42744 115810 42800
rect 115810 42744 115860 42800
rect 115796 42740 115860 42744
rect 116900 42740 116964 42804
rect 118372 42740 118436 42804
rect 119108 42800 119172 42804
rect 119108 42744 119122 42800
rect 119122 42744 119172 42800
rect 119108 42740 119172 42744
rect 133460 42800 133524 42804
rect 133460 42744 133474 42800
rect 133474 42744 133524 42800
rect 133460 42740 133524 42744
rect 136036 42740 136100 42804
rect 155908 42800 155972 42804
rect 155908 42744 155958 42800
rect 155958 42744 155972 42800
rect 155908 42740 155972 42744
rect 183508 42800 183572 42804
rect 183508 42744 183522 42800
rect 183522 42744 183572 42800
rect 183508 42740 183572 42744
rect 238156 42800 238220 42804
rect 238156 42744 238170 42800
rect 238170 42744 238220 42800
rect 238156 42740 238220 42744
rect 239260 42740 239324 42804
rect 240548 42800 240612 42804
rect 240548 42744 240562 42800
rect 240562 42744 240612 42800
rect 240548 42740 240612 42744
rect 241652 42800 241716 42804
rect 241652 42744 241666 42800
rect 241666 42744 241716 42800
rect 241652 42740 241716 42744
rect 245332 42800 245396 42804
rect 245332 42744 245346 42800
rect 245346 42744 245396 42800
rect 245332 42740 245396 42744
rect 246436 42800 246500 42804
rect 246436 42744 246450 42800
rect 246450 42744 246500 42800
rect 246436 42740 246500 42744
rect 250116 42800 250180 42804
rect 250116 42744 250130 42800
rect 250130 42744 250180 42800
rect 250116 42740 250180 42744
rect 251220 42800 251284 42804
rect 251220 42744 251234 42800
rect 251234 42744 251284 42800
rect 251220 42740 251284 42744
rect 253428 42800 253492 42804
rect 253428 42744 253442 42800
rect 253442 42744 253492 42800
rect 253428 42740 253492 42744
rect 260972 42800 261036 42804
rect 260972 42744 260986 42800
rect 260986 42744 261036 42800
rect 260972 42740 261036 42744
rect 268332 42740 268396 42804
rect 268700 42740 268764 42804
rect 271276 42800 271340 42804
rect 271276 42744 271290 42800
rect 271290 42744 271340 42800
rect 271276 42740 271340 42744
rect 273300 42800 273364 42804
rect 273300 42744 273314 42800
rect 273314 42744 273364 42800
rect 273300 42740 273364 42744
rect 276244 42740 276308 42804
rect 276980 42800 277044 42804
rect 276980 42744 276994 42800
rect 276994 42744 277044 42800
rect 276980 42740 277044 42744
rect 278084 42740 278148 42804
rect 293356 42800 293420 42804
rect 293356 42744 293370 42800
rect 293370 42744 293420 42800
rect 293356 42740 293420 42744
rect 298508 42800 298572 42804
rect 298508 42744 298522 42800
rect 298522 42744 298572 42800
rect 298508 42740 298572 42744
rect 303476 42740 303540 42804
rect 311020 42800 311084 42804
rect 311020 42744 311034 42800
rect 311034 42744 311084 42800
rect 311020 42740 311084 42744
rect 313412 42800 313476 42804
rect 313412 42744 313426 42800
rect 313426 42744 313476 42800
rect 313412 42740 313476 42744
rect 318380 42800 318444 42804
rect 318380 42744 318394 42800
rect 318394 42744 318444 42800
rect 318380 42740 318444 42744
rect 320956 42800 321020 42804
rect 320956 42744 320970 42800
rect 320970 42744 321020 42800
rect 320956 42740 321020 42744
rect 343220 42800 343284 42804
rect 343220 42744 343234 42800
rect 343234 42744 343284 42800
rect 343220 42740 343284 42744
rect 343404 42800 343468 42804
rect 343404 42744 343454 42800
rect 343454 42744 343468 42800
rect 343404 42740 343468 42744
rect 399524 42740 399588 42804
rect 408356 42800 408420 42804
rect 408356 42744 408370 42800
rect 408370 42744 408420 42800
rect 408356 42740 408420 42744
rect 408724 42800 408788 42804
rect 408724 42744 408738 42800
rect 408738 42744 408788 42800
rect 408724 42740 408788 42744
rect 410012 42800 410076 42804
rect 410012 42744 410026 42800
rect 410026 42744 410076 42800
rect 410012 42740 410076 42744
rect 411300 42800 411364 42804
rect 411300 42744 411314 42800
rect 411314 42744 411364 42800
rect 411300 42740 411364 42744
rect 412404 42740 412468 42804
rect 413324 42800 413388 42804
rect 413324 42744 413338 42800
rect 413338 42744 413388 42800
rect 413324 42740 413388 42744
rect 413692 42800 413756 42804
rect 413692 42744 413706 42800
rect 413706 42744 413756 42800
rect 413692 42740 413756 42744
rect 415532 42800 415596 42804
rect 415532 42744 415546 42800
rect 415546 42744 415596 42800
rect 415532 42740 415596 42744
rect 426388 42800 426452 42804
rect 426388 42744 426438 42800
rect 426438 42744 426452 42800
rect 426388 42740 426452 42744
rect 427676 42800 427740 42804
rect 427676 42744 427690 42800
rect 427690 42744 427740 42800
rect 427676 42740 427740 42744
rect 428596 42800 428660 42804
rect 428596 42744 428610 42800
rect 428610 42744 428660 42800
rect 428596 42740 428660 42744
rect 429700 42800 429764 42804
rect 429700 42744 429714 42800
rect 429714 42744 429764 42800
rect 429700 42740 429764 42744
rect 430988 42800 431052 42804
rect 430988 42744 431002 42800
rect 431002 42744 431052 42800
rect 430988 42740 431052 42744
rect 432276 42740 432340 42804
rect 433380 42800 433444 42804
rect 433380 42744 433394 42800
rect 433394 42744 433444 42800
rect 433380 42740 433444 42744
rect 434668 42800 434732 42804
rect 434668 42744 434682 42800
rect 434682 42744 434732 42800
rect 434668 42740 434732 42744
rect 435956 42800 436020 42804
rect 435956 42744 435970 42800
rect 435970 42744 436020 42800
rect 435956 42740 436020 42744
rect 436876 42740 436940 42804
rect 438532 42800 438596 42804
rect 438532 42744 438546 42800
rect 438546 42744 438596 42800
rect 438532 42740 438596 42744
rect 440924 42800 440988 42804
rect 440924 42744 440938 42800
rect 440938 42744 440988 42800
rect 440924 42740 440988 42744
rect 443500 42800 443564 42804
rect 443500 42744 443514 42800
rect 443514 42744 443564 42800
rect 443500 42740 443564 42744
rect 445892 42800 445956 42804
rect 445892 42744 445906 42800
rect 445906 42744 445956 42800
rect 445892 42740 445956 42744
rect 448284 42800 448348 42804
rect 448284 42744 448298 42800
rect 448298 42744 448348 42800
rect 448284 42740 448348 42744
rect 453436 42800 453500 42804
rect 453436 42744 453450 42800
rect 453450 42744 453500 42800
rect 453436 42740 453500 42744
rect 486004 42800 486068 42804
rect 486004 42744 486018 42800
rect 486018 42744 486068 42800
rect 486004 42740 486068 42744
rect 503116 42740 503180 42804
rect 503484 42800 503548 42804
rect 503484 42744 503534 42800
rect 503534 42744 503548 42800
rect 503484 42740 503548 42744
rect 60228 42604 60292 42668
rect 125916 42604 125980 42668
rect 183140 42664 183204 42668
rect 183140 42608 183190 42664
rect 183190 42608 183204 42664
rect 183140 42604 183204 42608
rect 215892 42604 215956 42668
rect 288204 42604 288268 42668
rect 370452 42604 370516 42668
rect 465948 42604 466012 42668
rect 54892 42468 54956 42532
rect 120764 42468 120828 42532
rect 165844 42528 165908 42532
rect 165844 42472 165858 42528
rect 165858 42472 165908 42528
rect 165844 42468 165908 42472
rect 210372 42468 210436 42532
rect 270908 42468 270972 42532
rect 376156 42468 376220 42532
rect 470916 42468 470980 42532
rect 57836 42332 57900 42396
rect 118004 42332 118068 42396
rect 214420 42332 214484 42396
rect 263548 42332 263612 42396
rect 266308 42392 266372 42396
rect 266308 42336 266358 42392
rect 266358 42336 266372 42392
rect 266308 42332 266372 42336
rect 267596 42332 267660 42396
rect 269804 42392 269868 42396
rect 269804 42336 269818 42392
rect 269818 42336 269868 42392
rect 269804 42332 269868 42336
rect 378732 42332 378796 42396
rect 460980 42332 461044 42396
rect 58940 42196 59004 42260
rect 105860 42196 105924 42260
rect 109540 42196 109604 42260
rect 111196 42256 111260 42260
rect 111196 42200 111210 42256
rect 111210 42200 111260 42256
rect 111196 42196 111260 42200
rect 206140 42196 206204 42260
rect 256004 42196 256068 42260
rect 274404 42196 274468 42260
rect 275324 42196 275388 42260
rect 374684 42196 374748 42260
rect 451044 42196 451108 42260
rect 58756 42060 58820 42124
rect 103836 42060 103900 42124
rect 207980 42060 208044 42124
rect 253612 42060 253676 42124
rect 254532 42060 254596 42124
rect 363460 42060 363524 42124
rect 433564 42060 433628 42124
rect 435772 42060 435836 42124
rect 58572 41924 58636 41988
rect 98500 41924 98564 41988
rect 208900 41924 208964 41988
rect 248276 41924 248340 41988
rect 248644 41984 248708 41988
rect 248644 41928 248658 41984
rect 248658 41928 248708 41984
rect 248644 41924 248708 41928
rect 252324 41924 252388 41988
rect 375972 41924 376036 41988
rect 416636 41924 416700 41988
rect 431172 41984 431236 41988
rect 431172 41928 431186 41984
rect 431186 41928 431236 41984
rect 431172 41924 431236 41928
rect 79548 41788 79612 41852
rect 81940 41788 82004 41852
rect 90036 41848 90100 41852
rect 90036 41792 90050 41848
rect 90050 41792 90100 41848
rect 90036 41788 90100 41792
rect 247724 41848 247788 41852
rect 247724 41792 247738 41848
rect 247738 41792 247788 41848
rect 247724 41788 247788 41792
rect 400444 41788 400508 41852
rect 200804 41652 200868 41716
rect 283788 41652 283852 41716
rect 55076 41516 55140 41580
rect 130884 41516 130948 41580
rect 378916 41516 378980 41580
rect 475884 41516 475948 41580
rect 163268 41380 163332 41444
rect 418476 41380 418540 41444
rect 438348 41380 438412 41444
rect 50660 41244 50724 41308
rect 219940 41244 220004 41308
rect 377812 41108 377876 41172
rect 377260 40972 377324 41036
rect 379468 40836 379532 40900
rect 53420 39884 53484 39948
rect 217548 39884 217612 39948
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 44955 483852 45021 483853
rect 44955 483788 44956 483852
rect 45020 483788 45021 483852
rect 44955 483787 45021 483788
rect 44771 483716 44837 483717
rect 44771 483652 44772 483716
rect 44836 483652 44837 483716
rect 44771 483651 44837 483652
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 44774 260133 44834 483651
rect 44958 260405 45018 483787
rect 45234 478894 45854 514338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 53051 646236 53117 646237
rect 53051 646172 53052 646236
rect 53116 646172 53117 646236
rect 53051 646171 53117 646172
rect 51579 646100 51645 646101
rect 51579 646036 51580 646100
rect 51644 646036 51645 646100
rect 51579 646035 51645 646036
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 46795 492284 46861 492285
rect 46795 492220 46796 492284
rect 46860 492220 46861 492284
rect 46795 492219 46861 492220
rect 46611 491876 46677 491877
rect 46611 491812 46612 491876
rect 46676 491812 46677 491876
rect 46611 491811 46677 491812
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 46427 463316 46493 463317
rect 46427 463252 46428 463316
rect 46492 463252 46493 463316
rect 46427 463251 46493 463252
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 44955 260404 45021 260405
rect 44955 260340 44956 260404
rect 45020 260340 45021 260404
rect 44955 260339 45021 260340
rect 44771 260132 44837 260133
rect 44771 260068 44772 260132
rect 44836 260068 44837 260132
rect 44771 260067 44837 260068
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 46430 43757 46490 463251
rect 46614 53957 46674 491811
rect 46611 53956 46677 53957
rect 46611 53892 46612 53956
rect 46676 53892 46677 53956
rect 46611 53891 46677 53892
rect 46798 52733 46858 492219
rect 47715 486980 47781 486981
rect 47715 486916 47716 486980
rect 47780 486916 47781 486980
rect 47715 486915 47781 486916
rect 47718 260813 47778 486915
rect 47899 483988 47965 483989
rect 47899 483924 47900 483988
rect 47964 483924 47965 483988
rect 47899 483923 47965 483924
rect 47715 260812 47781 260813
rect 47715 260748 47716 260812
rect 47780 260748 47781 260812
rect 47715 260747 47781 260748
rect 47902 238645 47962 483923
rect 48954 482614 49574 518058
rect 50843 492012 50909 492013
rect 50843 491948 50844 492012
rect 50908 491948 50909 492012
rect 50843 491947 50909 491948
rect 50291 491332 50357 491333
rect 50291 491268 50292 491332
rect 50356 491268 50357 491332
rect 50291 491267 50357 491268
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48083 465764 48149 465765
rect 48083 465700 48084 465764
rect 48148 465700 48149 465764
rect 48083 465699 48149 465700
rect 47899 238644 47965 238645
rect 47899 238580 47900 238644
rect 47964 238580 47965 238644
rect 47899 238579 47965 238580
rect 48086 152829 48146 465699
rect 48635 459644 48701 459645
rect 48635 459580 48636 459644
rect 48700 459580 48701 459644
rect 48635 459579 48701 459580
rect 48638 381037 48698 459579
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48635 381036 48701 381037
rect 48635 380972 48636 381036
rect 48700 380972 48701 381036
rect 48635 380971 48701 380972
rect 48954 374614 49574 410058
rect 50294 375325 50354 491267
rect 50475 460596 50541 460597
rect 50475 460532 50476 460596
rect 50540 460532 50541 460596
rect 50475 460531 50541 460532
rect 50291 375324 50357 375325
rect 50291 375260 50292 375324
rect 50356 375260 50357 375324
rect 50291 375259 50357 375260
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48083 152828 48149 152829
rect 48083 152764 48084 152828
rect 48148 152764 48149 152828
rect 48083 152763 48149 152764
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 46795 52732 46861 52733
rect 46795 52668 46796 52732
rect 46860 52668 46861 52732
rect 46795 52667 46861 52668
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 46427 43756 46493 43757
rect 46427 43692 46428 43756
rect 46492 43692 46493 43756
rect 46427 43691 46493 43692
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 50058
rect 50478 44573 50538 460531
rect 50659 459644 50725 459645
rect 50659 459580 50660 459644
rect 50724 459580 50725 459644
rect 50659 459579 50725 459580
rect 50475 44572 50541 44573
rect 50475 44508 50476 44572
rect 50540 44508 50541 44572
rect 50475 44507 50541 44508
rect 50662 41309 50722 459579
rect 50846 43893 50906 491947
rect 51582 219469 51642 646035
rect 52315 491332 52381 491333
rect 52315 491268 52316 491332
rect 52380 491268 52381 491332
rect 52315 491267 52381 491268
rect 52131 460188 52197 460189
rect 52131 460124 52132 460188
rect 52196 460124 52197 460188
rect 52131 460123 52197 460124
rect 51763 459644 51829 459645
rect 51763 459580 51764 459644
rect 51828 459580 51829 459644
rect 51763 459579 51829 459580
rect 51766 263669 51826 459579
rect 52134 372741 52194 460123
rect 52131 372740 52197 372741
rect 52131 372676 52132 372740
rect 52196 372676 52197 372740
rect 52131 372675 52197 372676
rect 51763 263668 51829 263669
rect 51763 263604 51764 263668
rect 51828 263604 51829 263668
rect 51763 263603 51829 263604
rect 51579 219468 51645 219469
rect 51579 219404 51580 219468
rect 51644 219404 51645 219468
rect 51579 219403 51645 219404
rect 52318 44029 52378 491267
rect 53054 269245 53114 646171
rect 54339 645964 54405 645965
rect 54339 645900 54340 645964
rect 54404 645900 54405 645964
rect 54339 645899 54405 645900
rect 53603 492148 53669 492149
rect 53603 492084 53604 492148
rect 53668 492084 53669 492148
rect 53603 492083 53669 492084
rect 53419 463180 53485 463181
rect 53419 463116 53420 463180
rect 53484 463116 53485 463180
rect 53419 463115 53485 463116
rect 53235 459644 53301 459645
rect 53235 459580 53236 459644
rect 53300 459580 53301 459644
rect 53235 459579 53301 459580
rect 53051 269244 53117 269245
rect 53051 269180 53052 269244
rect 53116 269180 53117 269244
rect 53051 269179 53117 269180
rect 53238 44165 53298 459579
rect 53235 44164 53301 44165
rect 53235 44100 53236 44164
rect 53300 44100 53301 44164
rect 53235 44099 53301 44100
rect 52315 44028 52381 44029
rect 52315 43964 52316 44028
rect 52380 43964 52381 44028
rect 52315 43963 52381 43964
rect 50843 43892 50909 43893
rect 50843 43828 50844 43892
rect 50908 43828 50909 43892
rect 50843 43827 50909 43828
rect 50659 41308 50725 41309
rect 50659 41244 50660 41308
rect 50724 41244 50725 41308
rect 50659 41243 50725 41244
rect 53422 39949 53482 463115
rect 53606 44301 53666 492083
rect 54342 320245 54402 645899
rect 55794 633454 56414 668898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 640099 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 640099 63854 640338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 640099 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 640099 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 640099 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 640099 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 640099 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 640099 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 640099 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 640099 99854 640338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 640099 103574 644058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 640099 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 640099 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 640099 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 640099 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 79568 633454 79888 633486
rect 79568 633218 79610 633454
rect 79846 633218 79888 633454
rect 79568 633134 79888 633218
rect 79568 632898 79610 633134
rect 79846 632898 79888 633134
rect 79568 632866 79888 632898
rect 110288 633454 110608 633486
rect 110288 633218 110330 633454
rect 110566 633218 110608 633454
rect 110288 633134 110608 633218
rect 110288 632898 110330 633134
rect 110566 632898 110608 633134
rect 110288 632866 110608 632898
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 79568 597454 79888 597486
rect 79568 597218 79610 597454
rect 79846 597218 79888 597454
rect 79568 597134 79888 597218
rect 79568 596898 79610 597134
rect 79846 596898 79888 597134
rect 79568 596866 79888 596898
rect 110288 597454 110608 597486
rect 110288 597218 110330 597454
rect 110566 597218 110608 597454
rect 110288 597134 110608 597218
rect 110288 596898 110330 597134
rect 110566 596898 110608 597134
rect 110288 596866 110608 596898
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 64208 579454 64528 579486
rect 64208 579218 64250 579454
rect 64486 579218 64528 579454
rect 64208 579134 64528 579218
rect 64208 578898 64250 579134
rect 64486 578898 64528 579134
rect 64208 578866 64528 578898
rect 94928 579454 95248 579486
rect 94928 579218 94970 579454
rect 95206 579218 95248 579454
rect 94928 579134 95248 579218
rect 94928 578898 94970 579134
rect 95206 578898 95248 579134
rect 94928 578866 95248 578898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 59514 565174 60134 573000
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 557000 60134 564618
rect 63234 568894 63854 573000
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 557000 63854 568338
rect 66954 572614 67574 573000
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 557000 67574 572058
rect 73794 562394 74414 573000
rect 73794 562158 73826 562394
rect 74062 562158 74146 562394
rect 74382 562158 74414 562394
rect 73794 562074 74414 562158
rect 73794 561838 73826 562074
rect 74062 561838 74146 562074
rect 74382 561838 74414 562074
rect 73794 557000 74414 561838
rect 77514 566114 78134 573000
rect 77514 565878 77546 566114
rect 77782 565878 77866 566114
rect 78102 565878 78134 566114
rect 77514 565794 78134 565878
rect 77514 565558 77546 565794
rect 77782 565558 77866 565794
rect 78102 565558 78134 565794
rect 77514 557000 78134 565558
rect 81234 567954 81854 573000
rect 81234 567718 81266 567954
rect 81502 567718 81586 567954
rect 81822 567718 81854 567954
rect 81234 567634 81854 567718
rect 81234 567398 81266 567634
rect 81502 567398 81586 567634
rect 81822 567398 81854 567634
rect 81234 557000 81854 567398
rect 84954 571674 85574 573000
rect 84954 571438 84986 571674
rect 85222 571438 85306 571674
rect 85542 571438 85574 571674
rect 84954 571354 85574 571438
rect 84954 571118 84986 571354
rect 85222 571118 85306 571354
rect 85542 571118 85574 571354
rect 84954 557000 85574 571118
rect 91794 561454 92414 573000
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 557000 92414 560898
rect 95514 565174 96134 573000
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 557000 96134 564618
rect 99234 568894 99854 573000
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 557000 99854 568338
rect 102954 572614 103574 573000
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 557000 103574 572058
rect 109794 562394 110414 573000
rect 109794 562158 109826 562394
rect 110062 562158 110146 562394
rect 110382 562158 110414 562394
rect 109794 562074 110414 562158
rect 109794 561838 109826 562074
rect 110062 561838 110146 562074
rect 110382 561838 110414 562074
rect 109794 557000 110414 561838
rect 113514 566114 114134 573000
rect 113514 565878 113546 566114
rect 113782 565878 113866 566114
rect 114102 565878 114134 566114
rect 113514 565794 114134 565878
rect 113514 565558 113546 565794
rect 113782 565558 113866 565794
rect 114102 565558 114134 565794
rect 113514 557000 114134 565558
rect 117234 567954 117854 573000
rect 117234 567718 117266 567954
rect 117502 567718 117586 567954
rect 117822 567718 117854 567954
rect 117234 567634 117854 567718
rect 117234 567398 117266 567634
rect 117502 567398 117586 567634
rect 117822 567398 117854 567634
rect 117234 557000 117854 567398
rect 120954 571674 121574 573000
rect 120954 571438 120986 571674
rect 121222 571438 121306 571674
rect 121542 571438 121574 571674
rect 120954 571354 121574 571438
rect 120954 571118 120986 571354
rect 121222 571118 121306 571354
rect 121542 571118 121574 571354
rect 120954 557000 121574 571118
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 557000 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 557000 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 640099 139574 644058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 640099 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 640099 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 640099 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 640099 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 640099 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 640099 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 640099 171854 640338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 640099 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 640099 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 640099 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 640099 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 640099 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 640099 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 159568 633454 159888 633486
rect 159568 633218 159610 633454
rect 159846 633218 159888 633454
rect 159568 633134 159888 633218
rect 159568 632898 159610 633134
rect 159846 632898 159888 633134
rect 159568 632866 159888 632898
rect 190288 633454 190608 633486
rect 190288 633218 190330 633454
rect 190566 633218 190608 633454
rect 190288 633134 190608 633218
rect 190288 632898 190330 633134
rect 190566 632898 190608 633134
rect 190288 632866 190608 632898
rect 144208 615454 144528 615486
rect 144208 615218 144250 615454
rect 144486 615218 144528 615454
rect 144208 615134 144528 615218
rect 144208 614898 144250 615134
rect 144486 614898 144528 615134
rect 144208 614866 144528 614898
rect 174928 615454 175248 615486
rect 174928 615218 174970 615454
rect 175206 615218 175248 615454
rect 174928 615134 175248 615218
rect 174928 614898 174970 615134
rect 175206 614898 175248 615134
rect 174928 614866 175248 614898
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 159568 597454 159888 597486
rect 159568 597218 159610 597454
rect 159846 597218 159888 597454
rect 159568 597134 159888 597218
rect 159568 596898 159610 597134
rect 159846 596898 159888 597134
rect 159568 596866 159888 596898
rect 190288 597454 190608 597486
rect 190288 597218 190330 597454
rect 190566 597218 190608 597454
rect 190288 597134 190608 597218
rect 190288 596898 190330 597134
rect 190566 596898 190608 597134
rect 190288 596866 190608 596898
rect 144208 579454 144528 579486
rect 144208 579218 144250 579454
rect 144486 579218 144528 579454
rect 144208 579134 144528 579218
rect 144208 578898 144250 579134
rect 144486 578898 144528 579134
rect 144208 578866 144528 578898
rect 174928 579454 175248 579486
rect 174928 579218 174970 579454
rect 175206 579218 175248 579454
rect 174928 579134 175248 579218
rect 174928 578898 174970 579134
rect 175206 578898 175248 579134
rect 174928 578866 175248 578898
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 557000 135854 568338
rect 138954 572614 139574 573000
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 557000 139574 572058
rect 145794 562394 146414 573000
rect 145794 562158 145826 562394
rect 146062 562158 146146 562394
rect 146382 562158 146414 562394
rect 145794 562074 146414 562158
rect 145794 561838 145826 562074
rect 146062 561838 146146 562074
rect 146382 561838 146414 562074
rect 145794 557000 146414 561838
rect 149514 566114 150134 573000
rect 149514 565878 149546 566114
rect 149782 565878 149866 566114
rect 150102 565878 150134 566114
rect 149514 565794 150134 565878
rect 149514 565558 149546 565794
rect 149782 565558 149866 565794
rect 150102 565558 150134 565794
rect 149514 557000 150134 565558
rect 153234 567954 153854 573000
rect 153234 567718 153266 567954
rect 153502 567718 153586 567954
rect 153822 567718 153854 567954
rect 153234 567634 153854 567718
rect 153234 567398 153266 567634
rect 153502 567398 153586 567634
rect 153822 567398 153854 567634
rect 153234 557000 153854 567398
rect 156954 571674 157574 573000
rect 156954 571438 156986 571674
rect 157222 571438 157306 571674
rect 157542 571438 157574 571674
rect 156954 571354 157574 571438
rect 156954 571118 156986 571354
rect 157222 571118 157306 571354
rect 157542 571118 157574 571354
rect 156954 557000 157574 571118
rect 163794 561454 164414 573000
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 557000 164414 560898
rect 167514 565174 168134 573000
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 557000 168134 564618
rect 171234 568894 171854 573000
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 557000 171854 568338
rect 174954 572614 175574 573000
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 557000 175574 572058
rect 181794 562394 182414 573000
rect 181794 562158 181826 562394
rect 182062 562158 182146 562394
rect 182382 562158 182414 562394
rect 181794 562074 182414 562158
rect 181794 561838 181826 562074
rect 182062 561838 182146 562074
rect 182382 561838 182414 562074
rect 181794 557000 182414 561838
rect 185514 566114 186134 573000
rect 185514 565878 185546 566114
rect 185782 565878 185866 566114
rect 186102 565878 186134 566114
rect 185514 565794 186134 565878
rect 185514 565558 185546 565794
rect 185782 565558 185866 565794
rect 186102 565558 186134 565794
rect 185514 557000 186134 565558
rect 189234 567954 189854 573000
rect 189234 567718 189266 567954
rect 189502 567718 189586 567954
rect 189822 567718 189854 567954
rect 189234 567634 189854 567718
rect 189234 567398 189266 567634
rect 189502 567398 189586 567634
rect 189822 567398 189854 567634
rect 189234 557000 189854 567398
rect 192954 571674 193574 573000
rect 192954 571438 192986 571674
rect 193222 571438 193306 571674
rect 193542 571438 193574 571674
rect 192954 571354 193574 571438
rect 192954 571118 192986 571354
rect 193222 571118 193306 571354
rect 193542 571118 193574 571354
rect 192954 557000 193574 571118
rect 199794 561454 200414 573000
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 557000 200414 560898
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 557000 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 557000 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 640099 218414 650898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 640099 222134 654618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 640099 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 640099 229574 662058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 640099 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 640099 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 640099 243854 640338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 640099 247574 644058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 640099 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 640099 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 640099 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 640099 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 640099 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 640099 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 640099 279854 640338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 640099 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 239568 633454 239888 633486
rect 239568 633218 239610 633454
rect 239846 633218 239888 633454
rect 239568 633134 239888 633218
rect 239568 632898 239610 633134
rect 239846 632898 239888 633134
rect 239568 632866 239888 632898
rect 270288 633454 270608 633486
rect 270288 633218 270330 633454
rect 270566 633218 270608 633454
rect 270288 633134 270608 633218
rect 270288 632898 270330 633134
rect 270566 632898 270608 633134
rect 270288 632866 270608 632898
rect 224208 615454 224528 615486
rect 224208 615218 224250 615454
rect 224486 615218 224528 615454
rect 224208 615134 224528 615218
rect 224208 614898 224250 615134
rect 224486 614898 224528 615134
rect 224208 614866 224528 614898
rect 254928 615454 255248 615486
rect 254928 615218 254970 615454
rect 255206 615218 255248 615454
rect 254928 615134 255248 615218
rect 254928 614898 254970 615134
rect 255206 614898 255248 615134
rect 254928 614866 255248 614898
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 239568 597454 239888 597486
rect 239568 597218 239610 597454
rect 239846 597218 239888 597454
rect 239568 597134 239888 597218
rect 239568 596898 239610 597134
rect 239846 596898 239888 597134
rect 239568 596866 239888 596898
rect 270288 597454 270608 597486
rect 270288 597218 270330 597454
rect 270566 597218 270608 597454
rect 270288 597134 270608 597218
rect 270288 596898 270330 597134
rect 270566 596898 270608 597134
rect 270288 596866 270608 596898
rect 224208 579454 224528 579486
rect 224208 579218 224250 579454
rect 224486 579218 224528 579454
rect 224208 579134 224528 579218
rect 224208 578898 224250 579134
rect 224486 578898 224528 579134
rect 224208 578866 224528 578898
rect 254928 579454 255248 579486
rect 254928 579218 254970 579454
rect 255206 579218 255248 579454
rect 254928 579134 255248 579218
rect 254928 578898 254970 579134
rect 255206 578898 255248 579134
rect 254928 578866 255248 578898
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 557000 211574 572058
rect 217794 562394 218414 573000
rect 217794 562158 217826 562394
rect 218062 562158 218146 562394
rect 218382 562158 218414 562394
rect 217794 562074 218414 562158
rect 217794 561838 217826 562074
rect 218062 561838 218146 562074
rect 218382 561838 218414 562074
rect 217794 557000 218414 561838
rect 221514 566114 222134 573000
rect 221514 565878 221546 566114
rect 221782 565878 221866 566114
rect 222102 565878 222134 566114
rect 221514 565794 222134 565878
rect 221514 565558 221546 565794
rect 221782 565558 221866 565794
rect 222102 565558 222134 565794
rect 221514 557000 222134 565558
rect 225234 567954 225854 573000
rect 225234 567718 225266 567954
rect 225502 567718 225586 567954
rect 225822 567718 225854 567954
rect 225234 567634 225854 567718
rect 225234 567398 225266 567634
rect 225502 567398 225586 567634
rect 225822 567398 225854 567634
rect 225234 557000 225854 567398
rect 228954 571674 229574 573000
rect 228954 571438 228986 571674
rect 229222 571438 229306 571674
rect 229542 571438 229574 571674
rect 228954 571354 229574 571438
rect 228954 571118 228986 571354
rect 229222 571118 229306 571354
rect 229542 571118 229574 571354
rect 228954 557000 229574 571118
rect 235794 561454 236414 573000
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 557000 236414 560898
rect 239514 565174 240134 573000
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 557000 240134 564618
rect 243234 568894 243854 573000
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 557000 243854 568338
rect 246954 572614 247574 573000
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 557000 247574 572058
rect 253794 562394 254414 573000
rect 253794 562158 253826 562394
rect 254062 562158 254146 562394
rect 254382 562158 254414 562394
rect 253794 562074 254414 562158
rect 253794 561838 253826 562074
rect 254062 561838 254146 562074
rect 254382 561838 254414 562074
rect 253794 557000 254414 561838
rect 257514 566114 258134 573000
rect 257514 565878 257546 566114
rect 257782 565878 257866 566114
rect 258102 565878 258134 566114
rect 257514 565794 258134 565878
rect 257514 565558 257546 565794
rect 257782 565558 257866 565794
rect 258102 565558 258134 565794
rect 257514 557000 258134 565558
rect 261234 567954 261854 573000
rect 261234 567718 261266 567954
rect 261502 567718 261586 567954
rect 261822 567718 261854 567954
rect 261234 567634 261854 567718
rect 261234 567398 261266 567634
rect 261502 567398 261586 567634
rect 261822 567398 261854 567634
rect 261234 557000 261854 567398
rect 264954 571674 265574 573000
rect 264954 571438 264986 571674
rect 265222 571438 265306 571674
rect 265542 571438 265574 571674
rect 264954 571354 265574 571438
rect 264954 571118 264986 571354
rect 265222 571118 265306 571354
rect 265542 571118 265574 571354
rect 264954 557000 265574 571118
rect 271794 561454 272414 573000
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 557000 272414 560898
rect 275514 565174 276134 573000
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 557000 276134 564618
rect 279234 568894 279854 573000
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 557000 279854 568338
rect 282954 572614 283574 573000
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 557000 283574 572058
rect 289794 557000 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 557000 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 557000 297854 586338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 557000 301574 590058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 64208 543454 64528 543486
rect 64208 543218 64250 543454
rect 64486 543218 64528 543454
rect 64208 543134 64528 543218
rect 64208 542898 64250 543134
rect 64486 542898 64528 543134
rect 64208 542866 64528 542898
rect 94928 543454 95248 543486
rect 94928 543218 94970 543454
rect 95206 543218 95248 543454
rect 94928 543134 95248 543218
rect 94928 542898 94970 543134
rect 95206 542898 95248 543134
rect 94928 542866 95248 542898
rect 125648 543454 125968 543486
rect 125648 543218 125690 543454
rect 125926 543218 125968 543454
rect 125648 543134 125968 543218
rect 125648 542898 125690 543134
rect 125926 542898 125968 543134
rect 125648 542866 125968 542898
rect 156368 543454 156688 543486
rect 156368 543218 156410 543454
rect 156646 543218 156688 543454
rect 156368 543134 156688 543218
rect 156368 542898 156410 543134
rect 156646 542898 156688 543134
rect 156368 542866 156688 542898
rect 187088 543454 187408 543486
rect 187088 543218 187130 543454
rect 187366 543218 187408 543454
rect 187088 543134 187408 543218
rect 187088 542898 187130 543134
rect 187366 542898 187408 543134
rect 187088 542866 187408 542898
rect 217808 543454 218128 543486
rect 217808 543218 217850 543454
rect 218086 543218 218128 543454
rect 217808 543134 218128 543218
rect 217808 542898 217850 543134
rect 218086 542898 218128 543134
rect 217808 542866 218128 542898
rect 248528 543454 248848 543486
rect 248528 543218 248570 543454
rect 248806 543218 248848 543454
rect 248528 543134 248848 543218
rect 248528 542898 248570 543134
rect 248806 542898 248848 543134
rect 248528 542866 248848 542898
rect 279248 543454 279568 543486
rect 279248 543218 279290 543454
rect 279526 543218 279568 543454
rect 279248 543134 279568 543218
rect 279248 542898 279290 543134
rect 279526 542898 279568 543134
rect 279248 542866 279568 542898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55075 491604 55141 491605
rect 55075 491540 55076 491604
rect 55140 491540 55141 491604
rect 55075 491539 55141 491540
rect 54891 460732 54957 460733
rect 54891 460668 54892 460732
rect 54956 460668 54957 460732
rect 54891 460667 54957 460668
rect 54707 460324 54773 460325
rect 54707 460260 54708 460324
rect 54772 460260 54773 460324
rect 54707 460259 54773 460260
rect 54339 320244 54405 320245
rect 54339 320180 54340 320244
rect 54404 320180 54405 320244
rect 54339 320179 54405 320180
rect 54710 129709 54770 460259
rect 54707 129708 54773 129709
rect 54707 129644 54708 129708
rect 54772 129644 54773 129708
rect 54707 129643 54773 129644
rect 53603 44300 53669 44301
rect 53603 44236 53604 44300
rect 53668 44236 53669 44300
rect 53603 44235 53669 44236
rect 54894 42533 54954 460667
rect 54891 42532 54957 42533
rect 54891 42468 54892 42532
rect 54956 42468 54957 42532
rect 54891 42467 54957 42468
rect 55078 41581 55138 491539
rect 55794 489454 56414 524898
rect 79568 525454 79888 525486
rect 79568 525218 79610 525454
rect 79846 525218 79888 525454
rect 79568 525134 79888 525218
rect 79568 524898 79610 525134
rect 79846 524898 79888 525134
rect 79568 524866 79888 524898
rect 110288 525454 110608 525486
rect 110288 525218 110330 525454
rect 110566 525218 110608 525454
rect 110288 525134 110608 525218
rect 110288 524898 110330 525134
rect 110566 524898 110608 525134
rect 110288 524866 110608 524898
rect 141008 525454 141328 525486
rect 141008 525218 141050 525454
rect 141286 525218 141328 525454
rect 141008 525134 141328 525218
rect 141008 524898 141050 525134
rect 141286 524898 141328 525134
rect 141008 524866 141328 524898
rect 171728 525454 172048 525486
rect 171728 525218 171770 525454
rect 172006 525218 172048 525454
rect 171728 525134 172048 525218
rect 171728 524898 171770 525134
rect 172006 524898 172048 525134
rect 171728 524866 172048 524898
rect 202448 525454 202768 525486
rect 202448 525218 202490 525454
rect 202726 525218 202768 525454
rect 202448 525134 202768 525218
rect 202448 524898 202490 525134
rect 202726 524898 202768 525134
rect 202448 524866 202768 524898
rect 233168 525454 233488 525486
rect 233168 525218 233210 525454
rect 233446 525218 233488 525454
rect 233168 525134 233488 525218
rect 233168 524898 233210 525134
rect 233446 524898 233488 525134
rect 233168 524866 233488 524898
rect 263888 525454 264208 525486
rect 263888 525218 263930 525454
rect 264166 525218 264208 525454
rect 263888 525134 264208 525218
rect 263888 524898 263930 525134
rect 264166 524898 264208 525134
rect 263888 524866 264208 524898
rect 294608 525454 294928 525486
rect 294608 525218 294650 525454
rect 294886 525218 294928 525454
rect 294608 525134 294928 525218
rect 294608 524898 294650 525134
rect 294886 524898 294928 525134
rect 294608 524866 294928 524898
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 59307 492556 59373 492557
rect 59307 492492 59308 492556
rect 59372 492492 59373 492556
rect 59307 492491 59373 492492
rect 59123 491740 59189 491741
rect 59123 491676 59124 491740
rect 59188 491676 59189 491740
rect 59123 491675 59189 491676
rect 57099 489700 57165 489701
rect 57099 489636 57100 489700
rect 57164 489636 57165 489700
rect 57099 489635 57165 489636
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55627 460460 55693 460461
rect 55627 460396 55628 460460
rect 55692 460396 55693 460460
rect 55627 460395 55693 460396
rect 55443 459644 55509 459645
rect 55443 459580 55444 459644
rect 55508 459580 55509 459644
rect 55443 459579 55509 459580
rect 55446 372741 55506 459579
rect 55443 372740 55509 372741
rect 55443 372676 55444 372740
rect 55508 372676 55509 372740
rect 55443 372675 55509 372676
rect 55630 44437 55690 460395
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 57102 319973 57162 489635
rect 58939 463452 59005 463453
rect 58939 463388 58940 463452
rect 59004 463388 59005 463452
rect 58939 463387 59005 463388
rect 58755 460868 58821 460869
rect 58755 460804 58756 460868
rect 58820 460804 58821 460868
rect 58755 460803 58821 460804
rect 58571 460052 58637 460053
rect 58571 459988 58572 460052
rect 58636 459988 58637 460052
rect 58571 459987 58637 459988
rect 57467 459100 57533 459101
rect 57467 459036 57468 459100
rect 57532 459036 57533 459100
rect 57467 459035 57533 459036
rect 57099 319972 57165 319973
rect 57099 319908 57100 319972
rect 57164 319908 57165 319972
rect 57099 319907 57165 319908
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 57099 237420 57165 237421
rect 57099 237356 57100 237420
rect 57164 237356 57165 237420
rect 57099 237355 57165 237356
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57102 133789 57162 237355
rect 57470 163029 57530 459035
rect 57835 458964 57901 458965
rect 57835 458900 57836 458964
rect 57900 458900 57901 458964
rect 57835 458899 57901 458900
rect 57651 458828 57717 458829
rect 57651 458764 57652 458828
rect 57716 458764 57717 458828
rect 57651 458763 57717 458764
rect 57467 163028 57533 163029
rect 57467 162964 57468 163028
rect 57532 162964 57533 163028
rect 57467 162963 57533 162964
rect 57654 154461 57714 458763
rect 57651 154460 57717 154461
rect 57651 154396 57652 154460
rect 57716 154396 57717 154460
rect 57651 154395 57717 154396
rect 57838 154325 57898 458899
rect 57835 154324 57901 154325
rect 57835 154260 57836 154324
rect 57900 154260 57901 154324
rect 57835 154259 57901 154260
rect 57835 150516 57901 150517
rect 57835 150452 57836 150516
rect 57900 150452 57901 150516
rect 57835 150451 57901 150452
rect 57099 133788 57165 133789
rect 57099 133724 57100 133788
rect 57164 133724 57165 133788
rect 57099 133723 57165 133724
rect 57099 132428 57165 132429
rect 57099 132364 57100 132428
rect 57164 132364 57165 132428
rect 57099 132363 57165 132364
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55627 44436 55693 44437
rect 55627 44372 55628 44436
rect 55692 44372 55693 44436
rect 55627 44371 55693 44372
rect 55075 41580 55141 41581
rect 55075 41516 55076 41580
rect 55140 41516 55141 41580
rect 55075 41515 55141 41516
rect 53419 39948 53485 39949
rect 53419 39884 53420 39948
rect 53484 39884 53485 39948
rect 53419 39883 53485 39884
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 56898
rect 57102 43485 57162 132363
rect 57283 130388 57349 130389
rect 57283 130324 57284 130388
rect 57348 130324 57349 130388
rect 57283 130323 57349 130324
rect 57286 129573 57346 130323
rect 57283 129572 57349 129573
rect 57283 129508 57284 129572
rect 57348 129508 57349 129572
rect 57283 129507 57349 129508
rect 57286 44709 57346 129507
rect 57283 44708 57349 44709
rect 57283 44644 57284 44708
rect 57348 44644 57349 44708
rect 57283 44643 57349 44644
rect 57099 43484 57165 43485
rect 57099 43420 57100 43484
rect 57164 43420 57165 43484
rect 57099 43419 57165 43420
rect 57838 42397 57898 150451
rect 57835 42396 57901 42397
rect 57835 42332 57836 42396
rect 57900 42332 57901 42396
rect 57835 42331 57901 42332
rect 58574 41989 58634 459987
rect 58758 42125 58818 460803
rect 58942 42261 59002 463387
rect 59126 43349 59186 491675
rect 59310 43621 59370 492491
rect 59514 476114 60134 493000
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 60134 476114
rect 59514 475794 60134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 60134 475794
rect 59514 460308 60134 475558
rect 63234 477954 63854 493000
rect 63234 477718 63266 477954
rect 63502 477718 63586 477954
rect 63822 477718 63854 477954
rect 63234 477634 63854 477718
rect 63234 477398 63266 477634
rect 63502 477398 63586 477634
rect 63822 477398 63854 477634
rect 60227 461548 60293 461549
rect 60227 461484 60228 461548
rect 60292 461484 60293 461548
rect 60227 461483 60293 461484
rect 60230 458690 60290 461483
rect 63234 460308 63854 477398
rect 66954 464614 67574 493000
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 460308 67574 464058
rect 73794 471454 74414 493000
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 460308 74414 470898
rect 77514 475174 78134 493000
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 460308 78134 474618
rect 81234 478894 81854 493000
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 460308 81854 478338
rect 84954 482614 85574 493000
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 460308 85574 482058
rect 91794 489454 92414 493000
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 460308 92414 488898
rect 95514 476114 96134 493000
rect 95514 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 96134 476114
rect 95514 475794 96134 475878
rect 95514 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 96134 475794
rect 95514 460308 96134 475558
rect 99234 477954 99854 493000
rect 99234 477718 99266 477954
rect 99502 477718 99586 477954
rect 99822 477718 99854 477954
rect 99234 477634 99854 477718
rect 99234 477398 99266 477634
rect 99502 477398 99586 477634
rect 99822 477398 99854 477634
rect 99234 460308 99854 477398
rect 102954 464614 103574 493000
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 460308 103574 464058
rect 109794 471454 110414 493000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 460308 110414 470898
rect 113514 475174 114134 493000
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 460308 114134 474618
rect 117234 478894 117854 493000
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 460308 117854 478338
rect 120954 482614 121574 493000
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 460308 121574 482058
rect 127794 489454 128414 493000
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 460308 128414 488898
rect 131514 476114 132134 493000
rect 131514 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 132134 476114
rect 131514 475794 132134 475878
rect 131514 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 132134 475794
rect 131514 460308 132134 475558
rect 135234 477954 135854 493000
rect 135234 477718 135266 477954
rect 135502 477718 135586 477954
rect 135822 477718 135854 477954
rect 135234 477634 135854 477718
rect 135234 477398 135266 477634
rect 135502 477398 135586 477634
rect 135822 477398 135854 477634
rect 135234 460308 135854 477398
rect 138954 464614 139574 493000
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 460308 139574 464058
rect 145794 471454 146414 493000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 460308 146414 470898
rect 149514 475174 150134 493000
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 460308 150134 474618
rect 153234 478894 153854 493000
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 460308 153854 478338
rect 156954 482614 157574 493000
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 460308 157574 482058
rect 163794 489454 164414 493000
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 460308 164414 488898
rect 167514 476114 168134 493000
rect 167514 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 168134 476114
rect 167514 475794 168134 475878
rect 167514 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 168134 475794
rect 167514 460308 168134 475558
rect 171234 477954 171854 493000
rect 171234 477718 171266 477954
rect 171502 477718 171586 477954
rect 171822 477718 171854 477954
rect 171234 477634 171854 477718
rect 171234 477398 171266 477634
rect 171502 477398 171586 477634
rect 171822 477398 171854 477634
rect 171234 460308 171854 477398
rect 174954 464614 175574 493000
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 460308 175574 464058
rect 181794 471454 182414 493000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 179643 462228 179709 462229
rect 179643 462164 179644 462228
rect 179708 462164 179709 462228
rect 179643 462163 179709 462164
rect 178355 461412 178421 461413
rect 178355 461348 178356 461412
rect 178420 461348 178421 461412
rect 178355 461347 178421 461348
rect 59862 458630 60290 458690
rect 178358 458690 178418 461347
rect 179646 458690 179706 462163
rect 181794 460308 182414 470898
rect 185514 475174 186134 493000
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 460308 186134 474618
rect 189234 478894 189854 493000
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 460308 189854 478338
rect 192954 482614 193574 493000
rect 196571 492556 196637 492557
rect 196571 492492 196572 492556
rect 196636 492492 196637 492556
rect 196571 492491 196637 492492
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 190867 461004 190933 461005
rect 190867 460940 190868 461004
rect 190932 460940 190933 461004
rect 190867 460939 190933 460940
rect 190870 458690 190930 460939
rect 192954 460308 193574 482058
rect 178358 458630 178524 458690
rect 179646 458630 179748 458690
rect 59862 374010 59922 458630
rect 178464 458202 178524 458630
rect 179688 458202 179748 458630
rect 190840 458630 190930 458690
rect 190840 458202 190900 458630
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 60952 399454 61300 399486
rect 60952 399218 61008 399454
rect 61244 399218 61300 399454
rect 60952 399134 61300 399218
rect 60952 398898 61008 399134
rect 61244 398898 61300 399134
rect 60952 398866 61300 398898
rect 195320 399454 195668 399486
rect 195320 399218 195376 399454
rect 195612 399218 195668 399454
rect 195320 399134 195668 399218
rect 195320 398898 195376 399134
rect 195612 398898 195668 399134
rect 195320 398866 195668 398898
rect 60272 381454 60620 381486
rect 60272 381218 60328 381454
rect 60564 381218 60620 381454
rect 60272 381134 60620 381218
rect 60272 380898 60328 381134
rect 60564 380898 60620 381134
rect 60272 380866 60620 380898
rect 196000 381454 196348 381486
rect 196000 381218 196056 381454
rect 196292 381218 196348 381454
rect 196000 381134 196348 381218
rect 196000 380898 196056 381134
rect 196292 380898 196348 381134
rect 196000 380866 196348 380898
rect 105491 375052 105557 375053
rect 76086 374990 76666 375050
rect 59862 373950 60290 374010
rect 59514 366234 60134 373000
rect 59514 365998 59546 366234
rect 59782 365998 59866 366234
rect 60102 365998 60134 366234
rect 59514 365914 60134 365998
rect 59514 365678 59546 365914
rect 59782 365678 59866 365914
rect 60102 365678 60134 365914
rect 59514 350308 60134 365678
rect 60230 349890 60290 373950
rect 63234 352894 63854 373000
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 350308 63854 352338
rect 66954 356614 67574 373000
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 350308 67574 356058
rect 73794 363454 74414 373000
rect 76606 371789 76666 374990
rect 77158 371789 77218 375050
rect 76603 371788 76669 371789
rect 76603 371724 76604 371788
rect 76668 371724 76669 371788
rect 76603 371723 76669 371724
rect 77155 371788 77221 371789
rect 77155 371724 77156 371788
rect 77220 371724 77221 371788
rect 77155 371723 77221 371724
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 350308 74414 362898
rect 77514 367174 78134 373000
rect 78262 372333 78322 375050
rect 79622 374990 79978 375050
rect 80574 374990 81082 375050
rect 81798 374990 82002 375050
rect 83158 374990 83842 375050
rect 84246 374990 84578 375050
rect 79918 372469 79978 374990
rect 79915 372468 79981 372469
rect 79915 372404 79916 372468
rect 79980 372404 79981 372468
rect 79915 372403 79981 372404
rect 78259 372332 78325 372333
rect 78259 372268 78260 372332
rect 78324 372268 78325 372332
rect 78259 372267 78325 372268
rect 81022 371381 81082 374990
rect 81019 371380 81085 371381
rect 81019 371316 81020 371380
rect 81084 371316 81085 371380
rect 81019 371315 81085 371316
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 350308 78134 366618
rect 81234 370894 81854 373000
rect 81942 372061 82002 374990
rect 81939 372060 82005 372061
rect 81939 371996 81940 372060
rect 82004 371996 82005 372060
rect 81939 371995 82005 371996
rect 83782 371517 83842 374990
rect 84518 372469 84578 374990
rect 84702 374990 85470 375050
rect 86558 374990 86786 375050
rect 87646 374990 88074 375050
rect 88326 374990 88442 375050
rect 88734 374990 89362 375050
rect 84702 372605 84762 374990
rect 84699 372604 84765 372605
rect 84699 372540 84700 372604
rect 84764 372540 84765 372604
rect 84699 372539 84765 372540
rect 84515 372468 84581 372469
rect 84515 372404 84516 372468
rect 84580 372404 84581 372468
rect 84515 372403 84581 372404
rect 83779 371516 83845 371517
rect 83779 371452 83780 371516
rect 83844 371452 83845 371516
rect 83779 371451 83845 371452
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 350308 81854 370338
rect 84954 357554 85574 373000
rect 86726 372605 86786 374990
rect 88014 372605 88074 374990
rect 88382 373285 88442 374990
rect 88379 373284 88445 373285
rect 88379 373220 88380 373284
rect 88444 373220 88445 373284
rect 88379 373219 88445 373220
rect 89302 372605 89362 374990
rect 90038 372605 90098 375050
rect 90222 374990 90774 375050
rect 91318 374990 91570 375050
rect 92406 374990 92490 375050
rect 90222 373421 90282 374990
rect 90219 373420 90285 373421
rect 90219 373356 90220 373420
rect 90284 373356 90285 373420
rect 90219 373355 90285 373356
rect 91510 372605 91570 374990
rect 92430 373149 92490 374990
rect 93350 374990 93494 375050
rect 93630 374990 93778 375050
rect 94582 374990 95066 375050
rect 92427 373148 92493 373149
rect 92427 373084 92428 373148
rect 92492 373084 92493 373148
rect 92427 373083 92493 373084
rect 86723 372604 86789 372605
rect 86723 372540 86724 372604
rect 86788 372540 86789 372604
rect 86723 372539 86789 372540
rect 88011 372604 88077 372605
rect 88011 372540 88012 372604
rect 88076 372540 88077 372604
rect 88011 372539 88077 372540
rect 89299 372604 89365 372605
rect 89299 372540 89300 372604
rect 89364 372540 89365 372604
rect 89299 372539 89365 372540
rect 90035 372604 90101 372605
rect 90035 372540 90036 372604
rect 90100 372540 90101 372604
rect 90035 372539 90101 372540
rect 91507 372604 91573 372605
rect 91507 372540 91508 372604
rect 91572 372540 91573 372604
rect 91507 372539 91573 372540
rect 84954 357318 84986 357554
rect 85222 357318 85306 357554
rect 85542 357318 85574 357554
rect 84954 357234 85574 357318
rect 84954 356998 84986 357234
rect 85222 356998 85306 357234
rect 85542 356998 85574 357234
rect 84954 350308 85574 356998
rect 91794 362514 92414 373000
rect 93350 372605 93410 374990
rect 93718 373149 93778 374990
rect 95006 373693 95066 374990
rect 95912 374370 95972 375020
rect 96078 374990 96170 375050
rect 97030 374990 97642 375050
rect 98118 374990 98194 375050
rect 95912 374310 95986 374370
rect 95926 373693 95986 374310
rect 95003 373692 95069 373693
rect 95003 373628 95004 373692
rect 95068 373628 95069 373692
rect 95003 373627 95069 373628
rect 95923 373692 95989 373693
rect 95923 373628 95924 373692
rect 95988 373628 95989 373692
rect 95923 373627 95989 373628
rect 96110 373421 96170 374990
rect 97582 373693 97642 374990
rect 98134 373829 98194 374990
rect 98318 374990 98526 375050
rect 99478 374990 100034 375050
rect 100702 374990 100770 375050
rect 98131 373828 98197 373829
rect 98131 373764 98132 373828
rect 98196 373764 98197 373828
rect 98131 373763 98197 373764
rect 97579 373692 97645 373693
rect 97579 373628 97580 373692
rect 97644 373628 97645 373692
rect 97579 373627 97645 373628
rect 98318 373557 98378 374990
rect 98315 373556 98381 373557
rect 98315 373492 98316 373556
rect 98380 373492 98381 373556
rect 98315 373491 98381 373492
rect 96107 373420 96173 373421
rect 96107 373356 96108 373420
rect 96172 373356 96173 373420
rect 96107 373355 96173 373356
rect 93715 373148 93781 373149
rect 93715 373084 93716 373148
rect 93780 373084 93781 373148
rect 93715 373083 93781 373084
rect 93347 372604 93413 372605
rect 93347 372540 93348 372604
rect 93412 372540 93413 372604
rect 93347 372539 93413 372540
rect 91794 362278 91826 362514
rect 92062 362278 92146 362514
rect 92382 362278 92414 362514
rect 91794 362194 92414 362278
rect 91794 361958 91826 362194
rect 92062 361958 92146 362194
rect 92382 361958 92414 362194
rect 91794 350308 92414 361958
rect 95514 366234 96134 373000
rect 95514 365998 95546 366234
rect 95782 365998 95866 366234
rect 96102 365998 96134 366234
rect 95514 365914 96134 365998
rect 95514 365678 95546 365914
rect 95782 365678 95866 365914
rect 96102 365678 96134 365914
rect 95514 350308 96134 365678
rect 99234 352894 99854 373000
rect 99974 372605 100034 374990
rect 99971 372604 100037 372605
rect 99971 372540 99972 372604
rect 100036 372540 100037 372604
rect 99971 372539 100037 372540
rect 100710 371381 100770 374990
rect 100894 374990 101110 375050
rect 101790 374990 102058 375050
rect 100894 373285 100954 374990
rect 100891 373284 100957 373285
rect 100891 373220 100892 373284
rect 100956 373220 100957 373284
rect 100891 373219 100957 373220
rect 101998 371653 102058 374990
rect 102734 374990 102878 375050
rect 103286 374990 103558 375050
rect 103966 374990 104634 375050
rect 101995 371652 102061 371653
rect 101995 371588 101996 371652
rect 102060 371588 102061 371652
rect 101995 371587 102061 371588
rect 102734 371381 102794 374990
rect 103286 373829 103346 374990
rect 103283 373828 103349 373829
rect 103283 373764 103284 373828
rect 103348 373764 103349 373828
rect 103283 373763 103349 373764
rect 100707 371380 100773 371381
rect 100707 371316 100708 371380
rect 100772 371316 100773 371380
rect 100707 371315 100773 371316
rect 102731 371380 102797 371381
rect 102731 371316 102732 371380
rect 102796 371316 102797 371380
rect 102731 371315 102797 371316
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 350308 99854 352338
rect 102954 356614 103574 373000
rect 104574 372605 104634 374990
rect 104571 372604 104637 372605
rect 104571 372540 104572 372604
rect 104636 372540 104637 372604
rect 104571 372539 104637 372540
rect 105310 371381 105370 375050
rect 105491 374988 105492 375052
rect 105556 375050 105557 375052
rect 105556 374990 106006 375050
rect 106414 374990 107026 375050
rect 105556 374988 105557 374990
rect 105491 374987 105557 374988
rect 106966 371653 107026 374990
rect 107518 374990 107638 375050
rect 107886 374990 108318 375050
rect 108726 374990 108866 375050
rect 106963 371652 107029 371653
rect 106963 371588 106964 371652
rect 107028 371588 107029 371652
rect 106963 371587 107029 371588
rect 107518 371381 107578 374990
rect 107886 373557 107946 374990
rect 107883 373556 107949 373557
rect 107883 373492 107884 373556
rect 107948 373492 107949 373556
rect 107883 373491 107949 373492
rect 108806 371653 108866 374990
rect 109542 374990 109814 375050
rect 110462 374990 111038 375050
rect 111174 374990 111626 375050
rect 112262 374990 112914 375050
rect 109542 372333 109602 374990
rect 110462 373829 110522 374990
rect 110459 373828 110525 373829
rect 110459 373764 110460 373828
rect 110524 373764 110525 373828
rect 110459 373763 110525 373764
rect 109539 372332 109605 372333
rect 109539 372268 109540 372332
rect 109604 372268 109605 372332
rect 109539 372267 109605 372268
rect 108803 371652 108869 371653
rect 108803 371588 108804 371652
rect 108868 371588 108869 371652
rect 108803 371587 108869 371588
rect 105307 371380 105373 371381
rect 105307 371316 105308 371380
rect 105372 371316 105373 371380
rect 105307 371315 105373 371316
rect 107515 371380 107581 371381
rect 107515 371316 107516 371380
rect 107580 371316 107581 371380
rect 107515 371315 107581 371316
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 350308 103574 356058
rect 109794 363454 110414 373000
rect 111566 371653 111626 374990
rect 112854 372605 112914 374990
rect 113222 374990 113350 375050
rect 112851 372604 112917 372605
rect 112851 372540 112852 372604
rect 112916 372540 112917 372604
rect 112851 372539 112917 372540
rect 113222 372197 113282 374990
rect 113592 374370 113652 375020
rect 114438 374990 114570 375050
rect 113590 374310 113652 374370
rect 113590 373693 113650 374310
rect 113587 373692 113653 373693
rect 113587 373628 113588 373692
rect 113652 373628 113653 373692
rect 113587 373627 113653 373628
rect 113219 372196 113285 372197
rect 113219 372132 113220 372196
rect 113284 372132 113285 372196
rect 113219 372131 113285 372132
rect 111563 371652 111629 371653
rect 111563 371588 111564 371652
rect 111628 371588 111629 371652
rect 111563 371587 111629 371588
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 350308 110414 362898
rect 113514 367174 114134 373000
rect 114510 372605 114570 374990
rect 115768 374370 115828 375020
rect 116070 374990 116226 375050
rect 117022 374990 117146 375050
rect 118110 374990 118250 375050
rect 115768 374310 115858 374370
rect 114507 372604 114573 372605
rect 114507 372540 114508 372604
rect 114572 372540 114573 372604
rect 114507 372539 114573 372540
rect 115798 371381 115858 374310
rect 116166 373693 116226 374990
rect 116163 373692 116229 373693
rect 116163 373628 116164 373692
rect 116228 373628 116229 373692
rect 116163 373627 116229 373628
rect 117086 371653 117146 374990
rect 117083 371652 117149 371653
rect 117083 371588 117084 371652
rect 117148 371588 117149 371652
rect 117083 371587 117149 371588
rect 115795 371380 115861 371381
rect 115795 371316 115796 371380
rect 115860 371316 115861 371380
rect 115795 371315 115861 371316
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 350308 114134 366618
rect 117234 370894 117854 373000
rect 118190 372333 118250 374990
rect 118374 374990 118518 375050
rect 119198 374990 119906 375050
rect 120966 374990 121378 375050
rect 123550 374990 124138 375050
rect 118374 373693 118434 374990
rect 118371 373692 118437 373693
rect 118371 373628 118372 373692
rect 118436 373628 118437 373692
rect 118371 373627 118437 373628
rect 118187 372332 118253 372333
rect 118187 372268 118188 372332
rect 118252 372268 118253 372332
rect 118187 372267 118253 372268
rect 119846 371789 119906 374990
rect 121318 373693 121378 374990
rect 124078 373693 124138 374990
rect 125734 374990 125998 375050
rect 128310 374990 128922 375050
rect 131030 374990 131130 375050
rect 133478 374990 133706 375050
rect 135926 374990 136466 375050
rect 138510 374990 139226 375050
rect 125734 373693 125794 374990
rect 128862 373693 128922 374990
rect 131070 373693 131130 374990
rect 133646 373693 133706 374990
rect 136406 373693 136466 374990
rect 139166 373693 139226 374990
rect 140928 374917 140988 375020
rect 140925 374916 140991 374917
rect 140925 374852 140926 374916
rect 140990 374852 140991 374916
rect 140925 374851 140991 374852
rect 143512 374509 143572 375020
rect 145990 374990 146218 375050
rect 148574 374990 148978 375050
rect 151022 374990 151738 375050
rect 143509 374508 143575 374509
rect 143509 374444 143510 374508
rect 143574 374444 143575 374508
rect 143509 374443 143575 374444
rect 146158 374237 146218 374990
rect 148918 374373 148978 374990
rect 148915 374372 148981 374373
rect 148915 374308 148916 374372
rect 148980 374308 148981 374372
rect 148915 374307 148981 374308
rect 146155 374236 146221 374237
rect 146155 374172 146156 374236
rect 146220 374172 146221 374236
rect 146155 374171 146221 374172
rect 151678 373693 151738 374990
rect 153440 374509 153500 375020
rect 155918 374990 156522 375050
rect 153437 374508 153503 374509
rect 153437 374444 153438 374508
rect 153502 374444 153503 374508
rect 153437 374443 153503 374444
rect 121315 373692 121381 373693
rect 121315 373628 121316 373692
rect 121380 373628 121381 373692
rect 121315 373627 121381 373628
rect 124075 373692 124141 373693
rect 124075 373628 124076 373692
rect 124140 373628 124141 373692
rect 124075 373627 124141 373628
rect 125731 373692 125797 373693
rect 125731 373628 125732 373692
rect 125796 373628 125797 373692
rect 125731 373627 125797 373628
rect 128859 373692 128925 373693
rect 128859 373628 128860 373692
rect 128924 373628 128925 373692
rect 128859 373627 128925 373628
rect 131067 373692 131133 373693
rect 131067 373628 131068 373692
rect 131132 373628 131133 373692
rect 131067 373627 131133 373628
rect 133643 373692 133709 373693
rect 133643 373628 133644 373692
rect 133708 373628 133709 373692
rect 133643 373627 133709 373628
rect 136403 373692 136469 373693
rect 136403 373628 136404 373692
rect 136468 373628 136469 373692
rect 136403 373627 136469 373628
rect 139163 373692 139229 373693
rect 139163 373628 139164 373692
rect 139228 373628 139229 373692
rect 139163 373627 139229 373628
rect 151675 373692 151741 373693
rect 151675 373628 151676 373692
rect 151740 373628 151741 373692
rect 151675 373627 151741 373628
rect 156462 373557 156522 374990
rect 158486 374509 158546 375050
rect 160920 374509 160980 375020
rect 163368 374645 163428 375020
rect 165952 374645 166012 375020
rect 183142 374990 183254 375050
rect 163365 374644 163431 374645
rect 163365 374580 163366 374644
rect 163430 374580 163431 374644
rect 163365 374579 163431 374580
rect 165949 374644 166015 374645
rect 165949 374580 165950 374644
rect 166014 374580 166015 374644
rect 165949 374579 166015 374580
rect 158483 374508 158549 374509
rect 158483 374444 158484 374508
rect 158548 374444 158549 374508
rect 158483 374443 158549 374444
rect 160917 374508 160983 374509
rect 160917 374444 160918 374508
rect 160982 374444 160983 374508
rect 160917 374443 160983 374444
rect 156459 373556 156525 373557
rect 156459 373492 156460 373556
rect 156524 373492 156525 373556
rect 156459 373491 156525 373492
rect 119843 371788 119909 371789
rect 119843 371724 119844 371788
rect 119908 371724 119909 371788
rect 119843 371723 119909 371724
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 350308 117854 370338
rect 120954 357554 121574 373000
rect 120954 357318 120986 357554
rect 121222 357318 121306 357554
rect 121542 357318 121574 357554
rect 120954 357234 121574 357318
rect 120954 356998 120986 357234
rect 121222 356998 121306 357234
rect 121542 356998 121574 357234
rect 120954 350308 121574 356998
rect 127794 362514 128414 373000
rect 127794 362278 127826 362514
rect 128062 362278 128146 362514
rect 128382 362278 128414 362514
rect 127794 362194 128414 362278
rect 127794 361958 127826 362194
rect 128062 361958 128146 362194
rect 128382 361958 128414 362194
rect 127794 350308 128414 361958
rect 131514 366234 132134 373000
rect 131514 365998 131546 366234
rect 131782 365998 131866 366234
rect 132102 365998 132134 366234
rect 131514 365914 132134 365998
rect 131514 365678 131546 365914
rect 131782 365678 131866 365914
rect 132102 365678 132134 365914
rect 131514 350308 132134 365678
rect 135234 352894 135854 373000
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 350308 135854 352338
rect 138954 356614 139574 373000
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 350308 139574 356058
rect 145794 363454 146414 373000
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 350308 146414 362898
rect 149514 367174 150134 373000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 350308 150134 366618
rect 153234 370894 153854 373000
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 350308 153854 370338
rect 156954 357554 157574 373000
rect 156954 357318 156986 357554
rect 157222 357318 157306 357554
rect 157542 357318 157574 357554
rect 156954 357234 157574 357318
rect 156954 356998 156986 357234
rect 157222 356998 157306 357234
rect 157542 356998 157574 357234
rect 156954 350308 157574 356998
rect 163794 362514 164414 373000
rect 163794 362278 163826 362514
rect 164062 362278 164146 362514
rect 164382 362278 164414 362514
rect 163794 362194 164414 362278
rect 163794 361958 163826 362194
rect 164062 361958 164146 362194
rect 164382 361958 164414 362194
rect 163794 350308 164414 361958
rect 167514 366234 168134 373000
rect 167514 365998 167546 366234
rect 167782 365998 167866 366234
rect 168102 365998 168134 366234
rect 167514 365914 168134 365998
rect 167514 365678 167546 365914
rect 167782 365678 167866 365914
rect 168102 365678 168134 365914
rect 167514 350308 168134 365678
rect 171234 352894 171854 373000
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 350308 171854 352338
rect 174954 356614 175574 373000
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 350308 175574 356058
rect 181794 363454 182414 373000
rect 183142 372469 183202 374990
rect 183360 374370 183420 375020
rect 183326 374310 183420 374370
rect 183139 372468 183205 372469
rect 183139 372404 183140 372468
rect 183204 372404 183205 372468
rect 183139 372403 183205 372404
rect 183326 371925 183386 374310
rect 183323 371924 183389 371925
rect 183323 371860 183324 371924
rect 183388 371860 183389 371924
rect 183323 371859 183389 371860
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 178539 351932 178605 351933
rect 178539 351868 178540 351932
rect 178604 351868 178605 351932
rect 178539 351867 178605 351868
rect 59862 349830 60290 349890
rect 59862 263530 59922 349830
rect 178542 348530 178602 351867
rect 179643 350572 179709 350573
rect 179643 350508 179644 350572
rect 179708 350508 179709 350572
rect 179643 350507 179709 350508
rect 178464 348470 178602 348530
rect 179646 348530 179706 350507
rect 181794 350308 182414 362898
rect 185514 367174 186134 373000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 350308 186134 366618
rect 189234 370894 189854 373000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 350308 189854 370338
rect 192954 357554 193574 373000
rect 192954 357318 192986 357554
rect 193222 357318 193306 357554
rect 193542 357318 193574 357554
rect 192954 357234 193574 357318
rect 192954 356998 192986 357234
rect 193222 356998 193306 357234
rect 193542 356998 193574 357234
rect 190867 350572 190933 350573
rect 190867 350508 190868 350572
rect 190932 350508 190933 350572
rect 190867 350507 190933 350508
rect 190870 348530 190930 350507
rect 192954 350308 193574 356998
rect 179646 348470 179748 348530
rect 178464 348202 178524 348470
rect 179688 348202 179748 348470
rect 190840 348470 190930 348530
rect 190840 348202 190900 348470
rect 60272 345454 60620 345486
rect 60272 345218 60328 345454
rect 60564 345218 60620 345454
rect 60272 345134 60620 345218
rect 60272 344898 60328 345134
rect 60564 344898 60620 345134
rect 60272 344866 60620 344898
rect 196000 345454 196348 345486
rect 196000 345218 196056 345454
rect 196292 345218 196348 345454
rect 196000 345134 196348 345218
rect 196000 344898 196056 345134
rect 196292 344898 196348 345134
rect 196000 344866 196348 344898
rect 60952 327454 61300 327486
rect 60952 327218 61008 327454
rect 61244 327218 61300 327454
rect 60952 327134 61300 327218
rect 60952 326898 61008 327134
rect 61244 326898 61300 327134
rect 60952 326866 61300 326898
rect 195320 327454 195668 327486
rect 195320 327218 195376 327454
rect 195612 327218 195668 327454
rect 195320 327134 195668 327218
rect 195320 326898 195376 327134
rect 195612 326898 195668 327134
rect 195320 326866 195668 326898
rect 60272 309454 60620 309486
rect 60272 309218 60328 309454
rect 60564 309218 60620 309454
rect 60272 309134 60620 309218
rect 60272 308898 60328 309134
rect 60564 308898 60620 309134
rect 60272 308866 60620 308898
rect 196000 309454 196348 309486
rect 196000 309218 196056 309454
rect 196292 309218 196348 309454
rect 196000 309134 196348 309218
rect 196000 308898 196056 309134
rect 196292 308898 196348 309134
rect 196000 308866 196348 308898
rect 60952 291454 61300 291486
rect 60952 291218 61008 291454
rect 61244 291218 61300 291454
rect 60952 291134 61300 291218
rect 60952 290898 61008 291134
rect 61244 290898 61300 291134
rect 60952 290866 61300 290898
rect 195320 291454 195668 291486
rect 195320 291218 195376 291454
rect 195612 291218 195668 291454
rect 195320 291134 195668 291218
rect 195320 290898 195376 291134
rect 195612 290898 195668 291134
rect 195320 290866 195668 290898
rect 60272 273454 60620 273486
rect 60272 273218 60328 273454
rect 60564 273218 60620 273454
rect 60272 273134 60620 273218
rect 60272 272898 60328 273134
rect 60564 272898 60620 273134
rect 60272 272866 60620 272898
rect 196000 273454 196348 273486
rect 196000 273218 196056 273454
rect 196292 273218 196348 273454
rect 196000 273134 196348 273218
rect 196000 272898 196056 273134
rect 196292 272898 196348 273134
rect 196000 272866 196348 272898
rect 76056 264890 76116 265106
rect 76054 264830 76116 264890
rect 77144 264890 77204 265106
rect 78232 264890 78292 265106
rect 79592 264890 79652 265106
rect 80544 264890 80604 265106
rect 81768 264890 81828 265106
rect 83128 264890 83188 265106
rect 84216 264890 84276 265106
rect 85440 264890 85500 265106
rect 77144 264830 77218 264890
rect 78232 264830 78322 264890
rect 59862 263470 60290 263530
rect 59514 241174 60134 263000
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 240308 60134 240618
rect 60230 238770 60290 263470
rect 76054 263125 76114 264830
rect 77158 263261 77218 264830
rect 77155 263260 77221 263261
rect 77155 263196 77156 263260
rect 77220 263196 77221 263260
rect 77155 263195 77221 263196
rect 76051 263124 76117 263125
rect 76051 263060 76052 263124
rect 76116 263060 76117 263124
rect 76051 263059 76117 263060
rect 63234 244894 63854 263000
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 240308 63854 244338
rect 66954 248614 67574 263000
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 240308 67574 248058
rect 73794 255454 74414 263000
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 240308 74414 254898
rect 77514 259174 78134 263000
rect 78262 262309 78322 264830
rect 79550 264830 79652 264890
rect 80470 264830 80604 264890
rect 81758 264830 81828 264890
rect 83046 264830 83188 264890
rect 83966 264830 84276 264890
rect 85438 264830 85500 264890
rect 86528 264890 86588 265106
rect 87616 264890 87676 265106
rect 88296 264890 88356 265106
rect 88704 264890 88764 265106
rect 90064 264890 90124 265106
rect 86528 264830 86602 264890
rect 87616 264830 87706 264890
rect 88296 264830 88442 264890
rect 88704 264830 88810 264890
rect 79550 262853 79610 264830
rect 80470 263533 80530 264830
rect 80467 263532 80533 263533
rect 80467 263468 80468 263532
rect 80532 263468 80533 263532
rect 80467 263467 80533 263468
rect 81758 263261 81818 264830
rect 83046 263397 83106 264830
rect 83043 263396 83109 263397
rect 83043 263332 83044 263396
rect 83108 263332 83109 263396
rect 83043 263331 83109 263332
rect 81755 263260 81821 263261
rect 81755 263196 81756 263260
rect 81820 263196 81821 263260
rect 81755 263195 81821 263196
rect 81234 262894 81854 263000
rect 83966 262989 84026 264830
rect 85438 263261 85498 264830
rect 85435 263260 85501 263261
rect 85435 263196 85436 263260
rect 85500 263196 85501 263260
rect 85435 263195 85501 263196
rect 83963 262988 84029 262989
rect 83963 262924 83964 262988
rect 84028 262924 84029 262988
rect 83963 262923 84029 262924
rect 79547 262852 79613 262853
rect 79547 262788 79548 262852
rect 79612 262788 79613 262852
rect 79547 262787 79613 262788
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 78259 262308 78325 262309
rect 78259 262244 78260 262308
rect 78324 262244 78325 262308
rect 78259 262243 78325 262244
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 240308 78134 258618
rect 81234 240308 81854 262338
rect 84954 249554 85574 263000
rect 86542 262581 86602 264830
rect 87646 262989 87706 264830
rect 88382 263533 88442 264830
rect 88379 263532 88445 263533
rect 88379 263468 88380 263532
rect 88444 263468 88445 263532
rect 88379 263467 88445 263468
rect 88750 262989 88810 264830
rect 90038 264830 90124 264890
rect 90744 264890 90804 265106
rect 91288 264890 91348 265106
rect 92376 264890 92436 265106
rect 93464 264893 93524 265106
rect 93461 264892 93527 264893
rect 90744 264830 90834 264890
rect 91288 264830 91386 264890
rect 92376 264830 92490 264890
rect 90038 263533 90098 264830
rect 90774 263533 90834 264830
rect 91326 263533 91386 264830
rect 92430 263533 92490 264830
rect 93461 264828 93462 264892
rect 93526 264828 93527 264892
rect 93600 264890 93660 265106
rect 94552 264890 94612 265106
rect 93600 264830 93778 264890
rect 93461 264827 93527 264828
rect 93718 263533 93778 264830
rect 94454 264830 94612 264890
rect 95912 264890 95972 265106
rect 96048 264890 96108 265106
rect 97000 264890 97060 265106
rect 98088 264890 98148 265106
rect 98496 264890 98556 265106
rect 99448 264890 99508 265106
rect 95912 264830 95986 264890
rect 96048 264830 96170 264890
rect 97000 264830 97090 264890
rect 98088 264830 98194 264890
rect 98496 264830 98562 264890
rect 90035 263532 90101 263533
rect 90035 263468 90036 263532
rect 90100 263468 90101 263532
rect 90035 263467 90101 263468
rect 90771 263532 90837 263533
rect 90771 263468 90772 263532
rect 90836 263468 90837 263532
rect 90771 263467 90837 263468
rect 91323 263532 91389 263533
rect 91323 263468 91324 263532
rect 91388 263468 91389 263532
rect 91323 263467 91389 263468
rect 92427 263532 92493 263533
rect 92427 263468 92428 263532
rect 92492 263468 92493 263532
rect 92427 263467 92493 263468
rect 93715 263532 93781 263533
rect 93715 263468 93716 263532
rect 93780 263468 93781 263532
rect 93715 263467 93781 263468
rect 87643 262988 87709 262989
rect 87643 262924 87644 262988
rect 87708 262924 87709 262988
rect 87643 262923 87709 262924
rect 88747 262988 88813 262989
rect 88747 262924 88748 262988
rect 88812 262924 88813 262988
rect 88747 262923 88813 262924
rect 86539 262580 86605 262581
rect 86539 262516 86540 262580
rect 86604 262516 86605 262580
rect 86539 262515 86605 262516
rect 84954 249318 84986 249554
rect 85222 249318 85306 249554
rect 85542 249318 85574 249554
rect 84954 249234 85574 249318
rect 84954 248998 84986 249234
rect 85222 248998 85306 249234
rect 85542 248998 85574 249234
rect 84954 240308 85574 248998
rect 91794 254514 92414 263000
rect 94454 262717 94514 264830
rect 95926 263261 95986 264830
rect 96110 263533 96170 264830
rect 96107 263532 96173 263533
rect 96107 263468 96108 263532
rect 96172 263468 96173 263532
rect 96107 263467 96173 263468
rect 95923 263260 95989 263261
rect 95923 263196 95924 263260
rect 95988 263196 95989 263260
rect 95923 263195 95989 263196
rect 94451 262716 94517 262717
rect 94451 262652 94452 262716
rect 94516 262652 94517 262716
rect 94451 262651 94517 262652
rect 91794 254278 91826 254514
rect 92062 254278 92146 254514
rect 92382 254278 92414 254514
rect 91794 254194 92414 254278
rect 91794 253958 91826 254194
rect 92062 253958 92146 254194
rect 92382 253958 92414 254194
rect 91794 240308 92414 253958
rect 95514 241174 96134 263000
rect 97030 262309 97090 264830
rect 98134 262309 98194 264830
rect 98502 263533 98562 264830
rect 99422 264830 99508 264890
rect 100672 264890 100732 265106
rect 101080 264890 101140 265106
rect 100672 264830 100770 264890
rect 98499 263532 98565 263533
rect 98499 263468 98500 263532
rect 98564 263468 98565 263532
rect 98499 263467 98565 263468
rect 99422 263261 99482 264830
rect 99419 263260 99485 263261
rect 99419 263196 99420 263260
rect 99484 263196 99485 263260
rect 99419 263195 99485 263196
rect 97027 262308 97093 262309
rect 97027 262244 97028 262308
rect 97092 262244 97093 262308
rect 97027 262243 97093 262244
rect 98131 262308 98197 262309
rect 98131 262244 98132 262308
rect 98196 262244 98197 262308
rect 98131 262243 98197 262244
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 240308 96134 240618
rect 99234 244894 99854 263000
rect 100710 262989 100770 264830
rect 101078 264830 101140 264890
rect 101760 264890 101820 265106
rect 102848 264890 102908 265106
rect 103528 264890 103588 265106
rect 103936 264890 103996 265106
rect 101760 264830 101874 264890
rect 101078 263533 101138 264830
rect 101075 263532 101141 263533
rect 101075 263468 101076 263532
rect 101140 263468 101141 263532
rect 101075 263467 101141 263468
rect 100707 262988 100773 262989
rect 100707 262924 100708 262988
rect 100772 262924 100773 262988
rect 100707 262923 100773 262924
rect 101814 262717 101874 264830
rect 102734 264830 102908 264890
rect 103286 264830 103588 264890
rect 103838 264830 103996 264890
rect 105296 264890 105356 265106
rect 105976 264890 106036 265106
rect 105296 264830 105370 264890
rect 102734 262717 102794 264830
rect 103286 263533 103346 264830
rect 103283 263532 103349 263533
rect 103283 263468 103284 263532
rect 103348 263468 103349 263532
rect 103283 263467 103349 263468
rect 103838 263125 103898 264830
rect 103835 263124 103901 263125
rect 103835 263060 103836 263124
rect 103900 263060 103901 263124
rect 103835 263059 103901 263060
rect 101811 262716 101877 262717
rect 101811 262652 101812 262716
rect 101876 262652 101877 262716
rect 101811 262651 101877 262652
rect 102731 262716 102797 262717
rect 102731 262652 102732 262716
rect 102796 262652 102797 262716
rect 102731 262651 102797 262652
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 240308 99854 244338
rect 102954 248614 103574 263000
rect 105310 262717 105370 264830
rect 105862 264830 106036 264890
rect 106384 264890 106444 265106
rect 107608 264890 107668 265106
rect 108288 264890 108348 265106
rect 108696 264890 108756 265106
rect 109784 264890 109844 265106
rect 111008 264893 111068 265106
rect 106384 264830 106474 264890
rect 105862 263533 105922 264830
rect 105859 263532 105925 263533
rect 105859 263468 105860 263532
rect 105924 263468 105925 263532
rect 105859 263467 105925 263468
rect 105307 262716 105373 262717
rect 105307 262652 105308 262716
rect 105372 262652 105373 262716
rect 105307 262651 105373 262652
rect 106414 262445 106474 264830
rect 107518 264830 107668 264890
rect 108254 264830 108348 264890
rect 108622 264830 108756 264890
rect 109726 264830 109844 264890
rect 111005 264892 111071 264893
rect 106411 262444 106477 262445
rect 106411 262380 106412 262444
rect 106476 262380 106477 262444
rect 106411 262379 106477 262380
rect 107518 262309 107578 264830
rect 108254 263533 108314 264830
rect 108251 263532 108317 263533
rect 108251 263468 108252 263532
rect 108316 263468 108317 263532
rect 108251 263467 108317 263468
rect 108622 262717 108682 264830
rect 109726 263533 109786 264830
rect 111005 264828 111006 264892
rect 111070 264828 111071 264892
rect 111144 264890 111204 265106
rect 112232 264890 112292 265106
rect 111144 264830 111258 264890
rect 111005 264827 111071 264828
rect 109723 263532 109789 263533
rect 109723 263468 109724 263532
rect 109788 263468 109789 263532
rect 109723 263467 109789 263468
rect 108619 262716 108685 262717
rect 108619 262652 108620 262716
rect 108684 262652 108685 262716
rect 108619 262651 108685 262652
rect 107515 262308 107581 262309
rect 107515 262244 107516 262308
rect 107580 262244 107581 262308
rect 107515 262243 107581 262244
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 240308 103574 248058
rect 109794 255454 110414 263000
rect 111198 262309 111258 264830
rect 112118 264830 112292 264890
rect 113320 264890 113380 265106
rect 113592 264890 113652 265106
rect 114408 264890 114468 265106
rect 113320 264830 113466 264890
rect 112118 262853 112178 264830
rect 113406 263397 113466 264830
rect 113590 264830 113652 264890
rect 114326 264830 114468 264890
rect 115768 264890 115828 265106
rect 116040 264890 116100 265106
rect 116992 264890 117052 265106
rect 118080 264890 118140 265106
rect 118488 264890 118548 265106
rect 119168 264890 119228 265106
rect 115768 264830 115858 264890
rect 113590 263533 113650 264830
rect 113587 263532 113653 263533
rect 113587 263468 113588 263532
rect 113652 263468 113653 263532
rect 113587 263467 113653 263468
rect 113403 263396 113469 263397
rect 113403 263332 113404 263396
rect 113468 263332 113469 263396
rect 113403 263331 113469 263332
rect 112115 262852 112181 262853
rect 112115 262788 112116 262852
rect 112180 262788 112181 262852
rect 112115 262787 112181 262788
rect 111195 262308 111261 262309
rect 111195 262244 111196 262308
rect 111260 262244 111261 262308
rect 111195 262243 111261 262244
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 240308 110414 254898
rect 113514 259174 114134 263000
rect 114326 262309 114386 264830
rect 115798 262581 115858 264830
rect 115982 264830 116100 264890
rect 116902 264830 117052 264890
rect 118006 264830 118140 264890
rect 118374 264830 118548 264890
rect 119110 264830 119228 264890
rect 120936 264890 120996 265106
rect 123520 264890 123580 265106
rect 125968 264893 126028 265106
rect 128280 264893 128340 265106
rect 131000 264893 131060 265106
rect 133448 264893 133508 265106
rect 135896 264893 135956 265106
rect 138480 264893 138540 265106
rect 125965 264892 126031 264893
rect 120936 264830 121010 264890
rect 123520 264830 123586 264890
rect 115982 263533 116042 264830
rect 116902 263533 116962 264830
rect 118006 264213 118066 264830
rect 118003 264212 118069 264213
rect 118003 264148 118004 264212
rect 118068 264148 118069 264212
rect 118003 264147 118069 264148
rect 118374 263533 118434 264830
rect 115979 263532 116045 263533
rect 115979 263468 115980 263532
rect 116044 263468 116045 263532
rect 115979 263467 116045 263468
rect 116899 263532 116965 263533
rect 116899 263468 116900 263532
rect 116964 263468 116965 263532
rect 116899 263467 116965 263468
rect 118371 263532 118437 263533
rect 118371 263468 118372 263532
rect 118436 263468 118437 263532
rect 118371 263467 118437 263468
rect 117234 262894 117854 263000
rect 119110 262989 119170 264830
rect 120950 263533 121010 264830
rect 123526 263533 123586 264830
rect 125965 264828 125966 264892
rect 126030 264828 126031 264892
rect 128280 264892 128373 264893
rect 128280 264830 128308 264892
rect 125965 264827 126031 264828
rect 128307 264828 128308 264830
rect 128372 264828 128373 264892
rect 128307 264827 128373 264828
rect 130997 264892 131063 264893
rect 130997 264828 130998 264892
rect 131062 264828 131063 264892
rect 130997 264827 131063 264828
rect 133445 264892 133511 264893
rect 133445 264828 133446 264892
rect 133510 264828 133511 264892
rect 133445 264827 133511 264828
rect 135893 264892 135959 264893
rect 135893 264828 135894 264892
rect 135958 264828 135959 264892
rect 135893 264827 135959 264828
rect 138477 264892 138543 264893
rect 138477 264828 138478 264892
rect 138542 264828 138543 264892
rect 138477 264827 138543 264828
rect 140928 264757 140988 265106
rect 143512 264757 143572 265106
rect 145960 264757 146020 265106
rect 148544 264757 148604 265106
rect 150992 264890 151052 265106
rect 150942 264830 151052 264890
rect 153440 264890 153500 265106
rect 155888 264890 155948 265106
rect 158472 264890 158532 265106
rect 160920 264890 160980 265106
rect 153440 264830 153578 264890
rect 155888 264830 155970 264890
rect 158472 264830 158546 264890
rect 140925 264756 140991 264757
rect 140925 264692 140926 264756
rect 140990 264692 140991 264756
rect 140925 264691 140991 264692
rect 143509 264756 143575 264757
rect 143509 264692 143510 264756
rect 143574 264692 143575 264756
rect 143509 264691 143575 264692
rect 145957 264756 146023 264757
rect 145957 264692 145958 264756
rect 146022 264692 146023 264756
rect 145957 264691 146023 264692
rect 148541 264756 148607 264757
rect 148541 264692 148542 264756
rect 148606 264692 148607 264756
rect 148541 264691 148607 264692
rect 150942 263533 151002 264830
rect 120947 263532 121013 263533
rect 120947 263468 120948 263532
rect 121012 263468 121013 263532
rect 120947 263467 121013 263468
rect 123523 263532 123589 263533
rect 123523 263468 123524 263532
rect 123588 263468 123589 263532
rect 123523 263467 123589 263468
rect 150939 263532 151005 263533
rect 150939 263468 150940 263532
rect 151004 263468 151005 263532
rect 150939 263467 151005 263468
rect 153518 263397 153578 264830
rect 155910 263533 155970 264830
rect 158486 263533 158546 264830
rect 160878 264830 160980 264890
rect 163368 264890 163428 265106
rect 165952 264890 166012 265106
rect 183224 264890 183284 265106
rect 163368 264830 163514 264890
rect 165952 264830 166090 264890
rect 160878 263533 160938 264830
rect 163454 263533 163514 264830
rect 166030 263533 166090 264830
rect 183142 264830 183284 264890
rect 183360 264890 183420 265106
rect 183360 264830 183570 264890
rect 155907 263532 155973 263533
rect 155907 263468 155908 263532
rect 155972 263468 155973 263532
rect 155907 263467 155973 263468
rect 158483 263532 158549 263533
rect 158483 263468 158484 263532
rect 158548 263468 158549 263532
rect 158483 263467 158549 263468
rect 160875 263532 160941 263533
rect 160875 263468 160876 263532
rect 160940 263468 160941 263532
rect 160875 263467 160941 263468
rect 163451 263532 163517 263533
rect 163451 263468 163452 263532
rect 163516 263468 163517 263532
rect 163451 263467 163517 263468
rect 166027 263532 166093 263533
rect 166027 263468 166028 263532
rect 166092 263468 166093 263532
rect 166027 263467 166093 263468
rect 153515 263396 153581 263397
rect 153515 263332 153516 263396
rect 153580 263332 153581 263396
rect 153515 263331 153581 263332
rect 119107 262988 119173 262989
rect 119107 262924 119108 262988
rect 119172 262924 119173 262988
rect 119107 262923 119173 262924
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 115795 262580 115861 262581
rect 115795 262516 115796 262580
rect 115860 262516 115861 262580
rect 115795 262515 115861 262516
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 114323 262308 114389 262309
rect 114323 262244 114324 262308
rect 114388 262244 114389 262308
rect 114323 262243 114389 262244
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 240308 114134 258618
rect 117234 240308 117854 262338
rect 120954 249554 121574 263000
rect 120954 249318 120986 249554
rect 121222 249318 121306 249554
rect 121542 249318 121574 249554
rect 120954 249234 121574 249318
rect 120954 248998 120986 249234
rect 121222 248998 121306 249234
rect 121542 248998 121574 249234
rect 120954 240308 121574 248998
rect 127794 254514 128414 263000
rect 127794 254278 127826 254514
rect 128062 254278 128146 254514
rect 128382 254278 128414 254514
rect 127794 254194 128414 254278
rect 127794 253958 127826 254194
rect 128062 253958 128146 254194
rect 128382 253958 128414 254194
rect 127794 240308 128414 253958
rect 131514 241174 132134 263000
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 240308 132134 240618
rect 135234 244894 135854 263000
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 240308 135854 244338
rect 138954 248614 139574 263000
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 240308 139574 248058
rect 145794 255454 146414 263000
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 240308 146414 254898
rect 149514 259174 150134 263000
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 240308 150134 258618
rect 153234 262894 153854 263000
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 240308 153854 262338
rect 156954 249554 157574 263000
rect 156954 249318 156986 249554
rect 157222 249318 157306 249554
rect 157542 249318 157574 249554
rect 156954 249234 157574 249318
rect 156954 248998 156986 249234
rect 157222 248998 157306 249234
rect 157542 248998 157574 249234
rect 156954 240308 157574 248998
rect 163794 254514 164414 263000
rect 163794 254278 163826 254514
rect 164062 254278 164146 254514
rect 164382 254278 164414 254514
rect 163794 254194 164414 254278
rect 163794 253958 163826 254194
rect 164062 253958 164146 254194
rect 164382 253958 164414 254194
rect 163794 240308 164414 253958
rect 167514 241174 168134 263000
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 240308 168134 240618
rect 171234 244894 171854 263000
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 240308 171854 244338
rect 174954 248614 175574 263000
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 240308 175574 248058
rect 181794 255454 182414 263000
rect 183142 262445 183202 264830
rect 183139 262444 183205 262445
rect 183139 262380 183140 262444
rect 183204 262380 183205 262444
rect 183139 262379 183205 262380
rect 183510 262309 183570 264830
rect 196574 264757 196634 492491
rect 197859 492420 197925 492421
rect 197859 492356 197860 492420
rect 197924 492356 197925 492420
rect 197859 492355 197925 492356
rect 196755 491740 196821 491741
rect 196755 491676 196756 491740
rect 196820 491676 196821 491740
rect 196755 491675 196821 491676
rect 196758 264893 196818 491675
rect 196755 264892 196821 264893
rect 196755 264828 196756 264892
rect 196820 264828 196821 264892
rect 196755 264827 196821 264828
rect 196571 264756 196637 264757
rect 196571 264692 196572 264756
rect 196636 264692 196637 264756
rect 196571 264691 196637 264692
rect 183507 262308 183573 262309
rect 183507 262244 183508 262308
rect 183572 262244 183573 262308
rect 183507 262243 183573 262244
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 240308 182414 254898
rect 185514 259174 186134 263000
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 240308 186134 258618
rect 189234 262894 189854 263000
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 240308 189854 262338
rect 192954 249554 193574 263000
rect 192954 249318 192986 249554
rect 193222 249318 193306 249554
rect 193542 249318 193574 249554
rect 192954 249234 193574 249318
rect 192954 248998 192986 249234
rect 193222 248998 193306 249234
rect 193542 248998 193574 249234
rect 192954 240308 193574 248998
rect 178539 240276 178605 240277
rect 178539 240212 178540 240276
rect 178604 240212 178605 240276
rect 178539 240211 178605 240212
rect 179643 240276 179709 240277
rect 179643 240212 179644 240276
rect 179708 240212 179709 240276
rect 179643 240211 179709 240212
rect 190867 240276 190933 240277
rect 190867 240212 190868 240276
rect 190932 240212 190933 240276
rect 190867 240211 190933 240212
rect 178542 238770 178602 240211
rect 59862 238710 60290 238770
rect 178464 238710 178602 238770
rect 179646 238770 179706 240211
rect 190870 238770 190930 240211
rect 179646 238710 179748 238770
rect 59862 154730 59922 238710
rect 178464 238202 178524 238710
rect 179688 238202 179748 238710
rect 190840 238710 190930 238770
rect 190840 238202 190900 238710
rect 60272 237454 60620 237486
rect 60272 237218 60328 237454
rect 60564 237218 60620 237454
rect 60272 237134 60620 237218
rect 60272 236898 60328 237134
rect 60564 236898 60620 237134
rect 60272 236866 60620 236898
rect 196000 237454 196348 237486
rect 196000 237218 196056 237454
rect 196292 237218 196348 237454
rect 196000 237134 196348 237218
rect 196000 236898 196056 237134
rect 196292 236898 196348 237134
rect 196000 236866 196348 236898
rect 60952 219454 61300 219486
rect 60952 219218 61008 219454
rect 61244 219218 61300 219454
rect 60952 219134 61300 219218
rect 60952 218898 61008 219134
rect 61244 218898 61300 219134
rect 60952 218866 61300 218898
rect 195320 219454 195668 219486
rect 195320 219218 195376 219454
rect 195612 219218 195668 219454
rect 195320 219134 195668 219218
rect 195320 218898 195376 219134
rect 195612 218898 195668 219134
rect 195320 218866 195668 218898
rect 60272 201454 60620 201486
rect 60272 201218 60328 201454
rect 60564 201218 60620 201454
rect 60272 201134 60620 201218
rect 60272 200898 60328 201134
rect 60564 200898 60620 201134
rect 60272 200866 60620 200898
rect 196000 201454 196348 201486
rect 196000 201218 196056 201454
rect 196292 201218 196348 201454
rect 196000 201134 196348 201218
rect 196000 200898 196056 201134
rect 196292 200898 196348 201134
rect 196000 200866 196348 200898
rect 60952 183454 61300 183486
rect 60952 183218 61008 183454
rect 61244 183218 61300 183454
rect 60952 183134 61300 183218
rect 60952 182898 61008 183134
rect 61244 182898 61300 183134
rect 60952 182866 61300 182898
rect 195320 183454 195668 183486
rect 195320 183218 195376 183454
rect 195612 183218 195668 183454
rect 195320 183134 195668 183218
rect 195320 182898 195376 183134
rect 195612 182898 195668 183134
rect 195320 182866 195668 182898
rect 60272 165454 60620 165486
rect 60272 165218 60328 165454
rect 60564 165218 60620 165454
rect 60272 165134 60620 165218
rect 60272 164898 60328 165134
rect 60564 164898 60620 165134
rect 60272 164866 60620 164898
rect 196000 165454 196348 165486
rect 196000 165218 196056 165454
rect 196292 165218 196348 165454
rect 196000 165134 196348 165218
rect 196000 164898 196056 165134
rect 196292 164898 196348 165134
rect 196000 164866 196348 164898
rect 59862 154670 60290 154730
rect 59514 133174 60134 153000
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 130308 60134 132618
rect 60230 128370 60290 154670
rect 76056 154590 76116 155040
rect 76054 154530 76116 154590
rect 77144 154590 77204 155040
rect 78232 154590 78292 155040
rect 79592 154590 79652 155040
rect 80544 154590 80604 155040
rect 77144 154530 77218 154590
rect 78232 154530 78322 154590
rect 76054 153101 76114 154530
rect 76051 153100 76117 153101
rect 76051 153036 76052 153100
rect 76116 153036 76117 153100
rect 76051 153035 76117 153036
rect 63234 136894 63854 153000
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 130308 63854 136338
rect 66954 140614 67574 153000
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 130308 67574 140058
rect 73794 147454 74414 153000
rect 77158 152557 77218 154530
rect 78262 153101 78322 154530
rect 79550 154530 79652 154590
rect 80470 154530 80604 154590
rect 81768 154590 81828 155040
rect 83128 154590 83188 155040
rect 84216 154590 84276 155040
rect 85440 154590 85500 155040
rect 81768 154530 82002 154590
rect 79550 153101 79610 154530
rect 78259 153100 78325 153101
rect 78259 153036 78260 153100
rect 78324 153036 78325 153100
rect 78259 153035 78325 153036
rect 79547 153100 79613 153101
rect 79547 153036 79548 153100
rect 79612 153036 79613 153100
rect 79547 153035 79613 153036
rect 77155 152556 77221 152557
rect 77155 152492 77156 152556
rect 77220 152492 77221 152556
rect 77155 152491 77221 152492
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 130308 74414 146898
rect 77514 151174 78134 153000
rect 80470 152013 80530 154530
rect 81942 153101 82002 154530
rect 83046 154530 83188 154590
rect 83966 154530 84276 154590
rect 85438 154530 85500 154590
rect 86528 154590 86588 155040
rect 87616 154590 87676 155040
rect 88296 154590 88356 155040
rect 88704 154590 88764 155040
rect 90064 154590 90124 155040
rect 86528 154530 86602 154590
rect 87616 154530 87706 154590
rect 88296 154530 88442 154590
rect 88704 154530 88810 154590
rect 83046 153101 83106 154530
rect 81939 153100 82005 153101
rect 81939 153036 81940 153100
rect 82004 153036 82005 153100
rect 81939 153035 82005 153036
rect 83043 153100 83109 153101
rect 83043 153036 83044 153100
rect 83108 153036 83109 153100
rect 83043 153035 83109 153036
rect 80467 152012 80533 152013
rect 80467 151948 80468 152012
rect 80532 151948 80533 152012
rect 80467 151947 80533 151948
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 130308 78134 150618
rect 81234 137834 81854 153000
rect 83966 152010 84026 154530
rect 85438 153237 85498 154530
rect 85435 153236 85501 153237
rect 85435 153172 85436 153236
rect 85500 153172 85501 153236
rect 85435 153171 85501 153172
rect 86542 153101 86602 154530
rect 87646 153101 87706 154530
rect 86539 153100 86605 153101
rect 86539 153036 86540 153100
rect 86604 153036 86605 153100
rect 86539 153035 86605 153036
rect 87643 153100 87709 153101
rect 87643 153036 87644 153100
rect 87708 153036 87709 153100
rect 87643 153035 87709 153036
rect 84147 152012 84213 152013
rect 84147 152010 84148 152012
rect 83966 151950 84148 152010
rect 84147 151948 84148 151950
rect 84212 151948 84213 152012
rect 84147 151947 84213 151948
rect 81234 137598 81266 137834
rect 81502 137598 81586 137834
rect 81822 137598 81854 137834
rect 81234 137514 81854 137598
rect 81234 137278 81266 137514
rect 81502 137278 81586 137514
rect 81822 137278 81854 137514
rect 81234 130308 81854 137278
rect 84954 141554 85574 153000
rect 88382 152421 88442 154530
rect 88750 153101 88810 154530
rect 90038 154530 90124 154590
rect 90744 154590 90804 155040
rect 91288 154590 91348 155040
rect 92376 154590 92436 155040
rect 93464 154590 93524 155040
rect 90744 154530 90834 154590
rect 91288 154530 91386 154590
rect 90038 153101 90098 154530
rect 88747 153100 88813 153101
rect 88747 153036 88748 153100
rect 88812 153036 88813 153100
rect 88747 153035 88813 153036
rect 90035 153100 90101 153101
rect 90035 153036 90036 153100
rect 90100 153036 90101 153100
rect 90035 153035 90101 153036
rect 90774 152421 90834 154530
rect 91326 153101 91386 154530
rect 91510 154530 92436 154590
rect 93350 154530 93524 154590
rect 93600 154590 93660 155040
rect 94552 154590 94612 155040
rect 93600 154530 93778 154590
rect 91323 153100 91389 153101
rect 91323 153036 91324 153100
rect 91388 153036 91389 153100
rect 91323 153035 91389 153036
rect 91510 152829 91570 154530
rect 93350 153101 93410 154530
rect 93347 153100 93413 153101
rect 93347 153036 93348 153100
rect 93412 153036 93413 153100
rect 93347 153035 93413 153036
rect 91507 152828 91573 152829
rect 91507 152764 91508 152828
rect 91572 152764 91573 152828
rect 91507 152763 91573 152764
rect 88379 152420 88445 152421
rect 88379 152356 88380 152420
rect 88444 152356 88445 152420
rect 88379 152355 88445 152356
rect 90771 152420 90837 152421
rect 90771 152356 90772 152420
rect 90836 152356 90837 152420
rect 90771 152355 90837 152356
rect 84954 141318 84986 141554
rect 85222 141318 85306 141554
rect 85542 141318 85574 141554
rect 84954 141234 85574 141318
rect 84954 140998 84986 141234
rect 85222 140998 85306 141234
rect 85542 140998 85574 141234
rect 84954 130308 85574 140998
rect 91794 146514 92414 153000
rect 93718 152557 93778 154530
rect 94454 154530 94612 154590
rect 95912 154590 95972 155040
rect 96048 154733 96108 155040
rect 96045 154732 96111 154733
rect 96045 154668 96046 154732
rect 96110 154668 96111 154732
rect 96045 154667 96111 154668
rect 97000 154590 97060 155040
rect 98088 154590 98148 155040
rect 98496 154590 98556 155040
rect 99448 154590 99508 155040
rect 100672 154730 100732 155040
rect 100672 154670 100770 154730
rect 95912 154530 95986 154590
rect 97000 154530 97090 154590
rect 98088 154530 98194 154590
rect 98496 154530 98562 154590
rect 94454 153101 94514 154530
rect 95926 153237 95986 154530
rect 95923 153236 95989 153237
rect 95923 153172 95924 153236
rect 95988 153172 95989 153236
rect 95923 153171 95989 153172
rect 97030 153101 97090 154530
rect 98134 153101 98194 154530
rect 98502 154189 98562 154530
rect 99422 154530 99508 154590
rect 98499 154188 98565 154189
rect 98499 154124 98500 154188
rect 98564 154124 98565 154188
rect 98499 154123 98565 154124
rect 99422 153237 99482 154530
rect 99419 153236 99485 153237
rect 99419 153172 99420 153236
rect 99484 153172 99485 153236
rect 99419 153171 99485 153172
rect 100710 153101 100770 154670
rect 101080 154590 101140 155040
rect 101078 154530 101140 154590
rect 101760 154590 101820 155040
rect 102848 154590 102908 155040
rect 101760 154530 101874 154590
rect 101078 154189 101138 154530
rect 101075 154188 101141 154189
rect 101075 154124 101076 154188
rect 101140 154124 101141 154188
rect 101075 154123 101141 154124
rect 94451 153100 94517 153101
rect 94451 153036 94452 153100
rect 94516 153036 94517 153100
rect 94451 153035 94517 153036
rect 97027 153100 97093 153101
rect 97027 153036 97028 153100
rect 97092 153036 97093 153100
rect 97027 153035 97093 153036
rect 98131 153100 98197 153101
rect 98131 153036 98132 153100
rect 98196 153036 98197 153100
rect 98131 153035 98197 153036
rect 100707 153100 100773 153101
rect 100707 153036 100708 153100
rect 100772 153036 100773 153100
rect 100707 153035 100773 153036
rect 93715 152556 93781 152557
rect 93715 152492 93716 152556
rect 93780 152492 93781 152556
rect 93715 152491 93781 152492
rect 91794 146278 91826 146514
rect 92062 146278 92146 146514
rect 92382 146278 92414 146514
rect 91794 146194 92414 146278
rect 91794 145958 91826 146194
rect 92062 145958 92146 146194
rect 92382 145958 92414 146194
rect 91794 130308 92414 145958
rect 95514 133174 96134 153000
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 130308 96134 132618
rect 99234 136894 99854 153000
rect 101814 152829 101874 154530
rect 102734 154530 102908 154590
rect 103528 154590 103588 155040
rect 103936 154590 103996 155040
rect 103528 154530 103714 154590
rect 102734 153101 102794 154530
rect 102731 153100 102797 153101
rect 102731 153036 102732 153100
rect 102796 153036 102797 153100
rect 102731 153035 102797 153036
rect 101811 152828 101877 152829
rect 101811 152764 101812 152828
rect 101876 152764 101877 152828
rect 101811 152763 101877 152764
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 130308 99854 136338
rect 102954 140614 103574 153000
rect 103654 152826 103714 154530
rect 103838 154530 103996 154590
rect 105296 154590 105356 155040
rect 105976 154590 106036 155040
rect 105296 154530 105370 154590
rect 103838 153101 103898 154530
rect 103835 153100 103901 153101
rect 103835 153036 103836 153100
rect 103900 153036 103901 153100
rect 103835 153035 103901 153036
rect 103835 152828 103901 152829
rect 103835 152826 103836 152828
rect 103654 152766 103836 152826
rect 103835 152764 103836 152766
rect 103900 152764 103901 152828
rect 103835 152763 103901 152764
rect 105310 152149 105370 154530
rect 105862 154530 106036 154590
rect 106384 154590 106444 155040
rect 107608 154590 107668 155040
rect 108288 154590 108348 155040
rect 106384 154530 106474 154590
rect 105862 154189 105922 154530
rect 105859 154188 105925 154189
rect 105859 154124 105860 154188
rect 105924 154124 105925 154188
rect 105859 154123 105925 154124
rect 106414 153101 106474 154530
rect 107518 154530 107668 154590
rect 108254 154530 108348 154590
rect 108696 154590 108756 155040
rect 109784 154590 109844 155040
rect 108696 154530 108866 154590
rect 106411 153100 106477 153101
rect 106411 153036 106412 153100
rect 106476 153036 106477 153100
rect 106411 153035 106477 153036
rect 107518 152829 107578 154530
rect 108254 154189 108314 154530
rect 108251 154188 108317 154189
rect 108251 154124 108252 154188
rect 108316 154124 108317 154188
rect 108251 154123 108317 154124
rect 108806 153101 108866 154530
rect 109542 154530 109844 154590
rect 111008 154590 111068 155040
rect 111144 154590 111204 155040
rect 112232 154590 112292 155040
rect 113320 154733 113380 155040
rect 113317 154732 113383 154733
rect 113317 154668 113318 154732
rect 113382 154668 113383 154732
rect 113317 154667 113383 154668
rect 113592 154590 113652 155040
rect 111008 154530 111074 154590
rect 111144 154530 111258 154590
rect 108803 153100 108869 153101
rect 108803 153036 108804 153100
rect 108868 153036 108869 153100
rect 108803 153035 108869 153036
rect 109542 152829 109602 154530
rect 111014 153101 111074 154530
rect 111198 153101 111258 154530
rect 112118 154530 112292 154590
rect 113222 154530 113652 154590
rect 114408 154590 114468 155040
rect 115768 154590 115828 155040
rect 116040 154590 116100 155040
rect 114408 154530 114570 154590
rect 115768 154530 115858 154590
rect 112118 153101 112178 154530
rect 111011 153100 111077 153101
rect 111011 153036 111012 153100
rect 111076 153036 111077 153100
rect 111011 153035 111077 153036
rect 111195 153100 111261 153101
rect 111195 153036 111196 153100
rect 111260 153036 111261 153100
rect 111195 153035 111261 153036
rect 112115 153100 112181 153101
rect 112115 153036 112116 153100
rect 112180 153036 112181 153100
rect 112115 153035 112181 153036
rect 107515 152828 107581 152829
rect 107515 152764 107516 152828
rect 107580 152764 107581 152828
rect 107515 152763 107581 152764
rect 109539 152828 109605 152829
rect 109539 152764 109540 152828
rect 109604 152764 109605 152828
rect 109539 152763 109605 152764
rect 105307 152148 105373 152149
rect 105307 152084 105308 152148
rect 105372 152084 105373 152148
rect 105307 152083 105373 152084
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 130308 103574 140058
rect 109794 147454 110414 153000
rect 113222 152829 113282 154530
rect 114510 153101 114570 154530
rect 115798 153101 115858 154530
rect 115982 154530 116100 154590
rect 116992 154590 117052 155040
rect 118080 154590 118140 155040
rect 118488 154590 118548 155040
rect 119168 154590 119228 155040
rect 120936 154590 120996 155040
rect 123520 154730 123580 155040
rect 122974 154670 123580 154730
rect 122974 154590 123034 154670
rect 125968 154590 126028 155040
rect 128280 154730 128340 155040
rect 128280 154670 128554 154730
rect 116992 154530 117146 154590
rect 114507 153100 114573 153101
rect 114507 153036 114508 153100
rect 114572 153036 114573 153100
rect 114507 153035 114573 153036
rect 115795 153100 115861 153101
rect 115795 153036 115796 153100
rect 115860 153036 115861 153100
rect 115795 153035 115861 153036
rect 113219 152828 113285 152829
rect 113219 152764 113220 152828
rect 113284 152764 113285 152828
rect 113219 152763 113285 152764
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 130308 110414 146898
rect 113514 151174 114134 153000
rect 115982 152557 116042 154530
rect 117086 153101 117146 154530
rect 118006 154530 118140 154590
rect 118374 154530 118548 154590
rect 119110 154530 119228 154590
rect 120766 154530 120996 154590
rect 122606 154530 123034 154590
rect 125918 154530 126028 154590
rect 117083 153100 117149 153101
rect 117083 153036 117084 153100
rect 117148 153036 117149 153100
rect 117083 153035 117149 153036
rect 115979 152556 116045 152557
rect 115979 152492 115980 152556
rect 116044 152492 116045 152556
rect 115979 152491 116045 152492
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 130308 114134 150618
rect 117234 137834 117854 153000
rect 118006 152829 118066 154530
rect 118374 153101 118434 154530
rect 119110 153101 119170 154530
rect 118371 153100 118437 153101
rect 118371 153036 118372 153100
rect 118436 153036 118437 153100
rect 118371 153035 118437 153036
rect 119107 153100 119173 153101
rect 119107 153036 119108 153100
rect 119172 153036 119173 153100
rect 119107 153035 119173 153036
rect 120766 152829 120826 154530
rect 118003 152828 118069 152829
rect 118003 152764 118004 152828
rect 118068 152764 118069 152828
rect 118003 152763 118069 152764
rect 120763 152828 120829 152829
rect 120763 152764 120764 152828
rect 120828 152764 120829 152828
rect 120763 152763 120829 152764
rect 117234 137598 117266 137834
rect 117502 137598 117586 137834
rect 117822 137598 117854 137834
rect 117234 137514 117854 137598
rect 117234 137278 117266 137514
rect 117502 137278 117586 137514
rect 117822 137278 117854 137514
rect 117234 130308 117854 137278
rect 120954 141554 121574 153000
rect 122606 152829 122666 154530
rect 125918 153101 125978 154530
rect 128494 153101 128554 154670
rect 131000 154590 131060 155040
rect 133448 154730 133508 155040
rect 135896 154730 135956 155040
rect 138480 154730 138540 155040
rect 140928 154730 140988 155040
rect 133448 154670 133522 154730
rect 135896 154670 136098 154730
rect 130886 154530 131060 154590
rect 130886 153101 130946 154530
rect 133462 153101 133522 154670
rect 136038 153101 136098 154670
rect 138430 154670 138540 154730
rect 140822 154670 140988 154730
rect 143512 154730 143572 155040
rect 145960 154730 146020 155040
rect 148544 154730 148604 155040
rect 150992 154730 151052 155040
rect 153440 154730 153500 155040
rect 143512 154670 143642 154730
rect 145960 154670 146034 154730
rect 148544 154670 148610 154730
rect 138430 154325 138490 154670
rect 138427 154324 138493 154325
rect 138427 154260 138428 154324
rect 138492 154260 138493 154324
rect 138427 154259 138493 154260
rect 140822 154189 140882 154670
rect 143582 154189 143642 154670
rect 140819 154188 140885 154189
rect 140819 154124 140820 154188
rect 140884 154124 140885 154188
rect 140819 154123 140885 154124
rect 143579 154188 143645 154189
rect 143579 154124 143580 154188
rect 143644 154124 143645 154188
rect 143579 154123 143645 154124
rect 145974 154053 146034 154670
rect 148550 154461 148610 154670
rect 150942 154670 151052 154730
rect 153334 154670 153500 154730
rect 155888 154730 155948 155040
rect 158472 154730 158532 155040
rect 160920 154730 160980 155040
rect 163368 154733 163428 155040
rect 165952 154733 166012 155040
rect 155888 154670 155970 154730
rect 158472 154670 158546 154730
rect 148547 154460 148613 154461
rect 148547 154396 148548 154460
rect 148612 154396 148613 154460
rect 148547 154395 148613 154396
rect 150942 154053 151002 154670
rect 145971 154052 146037 154053
rect 145971 153988 145972 154052
rect 146036 153988 146037 154052
rect 145971 153987 146037 153988
rect 150939 154052 151005 154053
rect 150939 153988 150940 154052
rect 151004 153988 151005 154052
rect 150939 153987 151005 153988
rect 153334 153917 153394 154670
rect 153331 153916 153397 153917
rect 153331 153852 153332 153916
rect 153396 153852 153397 153916
rect 153331 153851 153397 153852
rect 155910 153101 155970 154670
rect 125915 153100 125981 153101
rect 125915 153036 125916 153100
rect 125980 153036 125981 153100
rect 125915 153035 125981 153036
rect 128491 153100 128557 153101
rect 128491 153036 128492 153100
rect 128556 153036 128557 153100
rect 128491 153035 128557 153036
rect 130883 153100 130949 153101
rect 130883 153036 130884 153100
rect 130948 153036 130949 153100
rect 130883 153035 130949 153036
rect 133459 153100 133525 153101
rect 133459 153036 133460 153100
rect 133524 153036 133525 153100
rect 133459 153035 133525 153036
rect 136035 153100 136101 153101
rect 136035 153036 136036 153100
rect 136100 153036 136101 153100
rect 136035 153035 136101 153036
rect 155907 153100 155973 153101
rect 155907 153036 155908 153100
rect 155972 153036 155973 153100
rect 155907 153035 155973 153036
rect 122603 152828 122669 152829
rect 122603 152764 122604 152828
rect 122668 152764 122669 152828
rect 122603 152763 122669 152764
rect 120954 141318 120986 141554
rect 121222 141318 121306 141554
rect 121542 141318 121574 141554
rect 120954 141234 121574 141318
rect 120954 140998 120986 141234
rect 121222 140998 121306 141234
rect 121542 140998 121574 141234
rect 120954 130308 121574 140998
rect 127794 146514 128414 153000
rect 127794 146278 127826 146514
rect 128062 146278 128146 146514
rect 128382 146278 128414 146514
rect 127794 146194 128414 146278
rect 127794 145958 127826 146194
rect 128062 145958 128146 146194
rect 128382 145958 128414 146194
rect 127794 130308 128414 145958
rect 131514 133174 132134 153000
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 130308 132134 132618
rect 135234 136894 135854 153000
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 130308 135854 136338
rect 138954 140614 139574 153000
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 130308 139574 140058
rect 145794 147454 146414 153000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 130308 146414 146898
rect 149514 151174 150134 153000
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 130308 150134 150618
rect 153234 137834 153854 153000
rect 153234 137598 153266 137834
rect 153502 137598 153586 137834
rect 153822 137598 153854 137834
rect 153234 137514 153854 137598
rect 153234 137278 153266 137514
rect 153502 137278 153586 137514
rect 153822 137278 153854 137514
rect 153234 130308 153854 137278
rect 156954 141554 157574 153000
rect 158486 152965 158546 154670
rect 160878 154670 160980 154730
rect 163365 154732 163431 154733
rect 158483 152964 158549 152965
rect 158483 152900 158484 152964
rect 158548 152900 158549 152964
rect 158483 152899 158549 152900
rect 160878 152693 160938 154670
rect 163365 154668 163366 154732
rect 163430 154668 163431 154732
rect 163365 154667 163431 154668
rect 165949 154732 166015 154733
rect 165949 154668 165950 154732
rect 166014 154668 166015 154732
rect 183224 154730 183284 155040
rect 165949 154667 166015 154668
rect 183142 154670 183284 154730
rect 183360 154730 183420 155040
rect 183360 154670 183570 154730
rect 160875 152692 160941 152693
rect 160875 152628 160876 152692
rect 160940 152628 160941 152692
rect 160875 152627 160941 152628
rect 156954 141318 156986 141554
rect 157222 141318 157306 141554
rect 157542 141318 157574 141554
rect 156954 141234 157574 141318
rect 156954 140998 156986 141234
rect 157222 140998 157306 141234
rect 157542 140998 157574 141234
rect 156954 130308 157574 140998
rect 163794 146514 164414 153000
rect 163794 146278 163826 146514
rect 164062 146278 164146 146514
rect 164382 146278 164414 146514
rect 163794 146194 164414 146278
rect 163794 145958 163826 146194
rect 164062 145958 164146 146194
rect 164382 145958 164414 146194
rect 163794 130308 164414 145958
rect 167514 133174 168134 153000
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 130308 168134 132618
rect 171234 136894 171854 153000
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 130308 171854 136338
rect 174954 140614 175574 153000
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 130308 175574 140058
rect 181794 147454 182414 153000
rect 183142 152829 183202 154670
rect 183139 152828 183205 152829
rect 183139 152764 183140 152828
rect 183204 152764 183205 152828
rect 183139 152763 183205 152764
rect 183510 152557 183570 154670
rect 183507 152556 183573 152557
rect 183507 152492 183508 152556
rect 183572 152492 183573 152556
rect 183507 152491 183573 152492
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 130308 182414 146898
rect 185514 151174 186134 153000
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 130308 186134 150618
rect 189234 137834 189854 153000
rect 189234 137598 189266 137834
rect 189502 137598 189586 137834
rect 189822 137598 189854 137834
rect 189234 137514 189854 137598
rect 189234 137278 189266 137514
rect 189502 137278 189586 137514
rect 189822 137278 189854 137514
rect 189234 130308 189854 137278
rect 192954 141554 193574 153000
rect 192954 141318 192986 141554
rect 193222 141318 193306 141554
rect 193542 141318 193574 141554
rect 192954 141234 193574 141318
rect 192954 140998 192986 141234
rect 193222 140998 193306 141234
rect 193542 140998 193574 141234
rect 190867 130388 190933 130389
rect 190867 130324 190868 130388
rect 190932 130324 190933 130388
rect 190867 130323 190933 130324
rect 178539 129844 178605 129845
rect 178539 129780 178540 129844
rect 178604 129780 178605 129844
rect 178539 129779 178605 129780
rect 179643 129844 179709 129845
rect 179643 129780 179644 129844
rect 179708 129780 179709 129844
rect 179643 129779 179709 129780
rect 178542 128890 178602 129779
rect 59862 128310 60290 128370
rect 178464 128830 178602 128890
rect 179646 128890 179706 129779
rect 190870 128890 190930 130323
rect 192954 130308 193574 140998
rect 179646 128830 179748 128890
rect 59862 43890 59922 128310
rect 178464 128202 178524 128830
rect 179688 128202 179748 128830
rect 190840 128830 190930 128890
rect 190840 128202 190900 128830
rect 60952 111454 61300 111486
rect 60952 111218 61008 111454
rect 61244 111218 61300 111454
rect 60952 111134 61300 111218
rect 60952 110898 61008 111134
rect 61244 110898 61300 111134
rect 60952 110866 61300 110898
rect 195320 111454 195668 111486
rect 195320 111218 195376 111454
rect 195612 111218 195668 111454
rect 195320 111134 195668 111218
rect 195320 110898 195376 111134
rect 195612 110898 195668 111134
rect 195320 110866 195668 110898
rect 60272 93454 60620 93486
rect 60272 93218 60328 93454
rect 60564 93218 60620 93454
rect 60272 93134 60620 93218
rect 60272 92898 60328 93134
rect 60564 92898 60620 93134
rect 60272 92866 60620 92898
rect 196000 93454 196348 93486
rect 196000 93218 196056 93454
rect 196292 93218 196348 93454
rect 196000 93134 196348 93218
rect 196000 92898 196056 93134
rect 196292 92898 196348 93134
rect 196000 92866 196348 92898
rect 60952 75454 61300 75486
rect 60952 75218 61008 75454
rect 61244 75218 61300 75454
rect 60952 75134 61300 75218
rect 60952 74898 61008 75134
rect 61244 74898 61300 75134
rect 60952 74866 61300 74898
rect 195320 75454 195668 75486
rect 195320 75218 195376 75454
rect 195612 75218 195668 75454
rect 195320 75134 195668 75218
rect 195320 74898 195376 75134
rect 195612 74898 195668 75134
rect 195320 74866 195668 74898
rect 60272 57454 60620 57486
rect 60272 57218 60328 57454
rect 60564 57218 60620 57454
rect 60272 57134 60620 57218
rect 60272 56898 60328 57134
rect 60564 56898 60620 57134
rect 60272 56866 60620 56898
rect 196000 57454 196348 57486
rect 196000 57218 196056 57454
rect 196292 57218 196348 57454
rect 196000 57134 196348 57218
rect 196000 56898 196056 57134
rect 196292 56898 196348 57134
rect 196000 56866 196348 56898
rect 76056 44570 76116 45106
rect 77144 44845 77204 45106
rect 77141 44844 77207 44845
rect 77141 44780 77142 44844
rect 77206 44780 77207 44844
rect 77141 44779 77207 44780
rect 76054 44510 76116 44570
rect 78232 44570 78292 45106
rect 79592 44570 79652 45106
rect 80544 44842 80604 45106
rect 78232 44510 78322 44570
rect 59862 43830 60290 43890
rect 59307 43620 59373 43621
rect 59307 43556 59308 43620
rect 59372 43556 59373 43620
rect 59307 43555 59373 43556
rect 59123 43348 59189 43349
rect 59123 43284 59124 43348
rect 59188 43284 59189 43348
rect 59123 43283 59189 43284
rect 58939 42260 59005 42261
rect 58939 42196 58940 42260
rect 59004 42196 59005 42260
rect 58939 42195 59005 42196
rect 58755 42124 58821 42125
rect 58755 42060 58756 42124
rect 58820 42060 58821 42124
rect 58755 42059 58821 42060
rect 58571 41988 58637 41989
rect 58571 41924 58572 41988
rect 58636 41924 58637 41988
rect 58571 41923 58637 41924
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 43000
rect 60230 42669 60290 43830
rect 60227 42668 60293 42669
rect 60227 42604 60228 42668
rect 60292 42604 60293 42668
rect 60227 42603 60293 42604
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 43000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 43000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 43000
rect 76054 42805 76114 44510
rect 76051 42804 76117 42805
rect 76051 42740 76052 42804
rect 76116 42740 76117 42804
rect 76051 42739 76117 42740
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 43000
rect 78262 42805 78322 44510
rect 79550 44510 79652 44570
rect 80470 44782 80604 44842
rect 78259 42804 78325 42805
rect 78259 42740 78260 42804
rect 78324 42740 78325 42804
rect 78259 42739 78325 42740
rect 79550 41853 79610 44510
rect 80470 42805 80530 44782
rect 81768 44570 81828 45106
rect 83128 44845 83188 45106
rect 84216 44845 84276 45106
rect 83125 44844 83191 44845
rect 83125 44780 83126 44844
rect 83190 44780 83191 44844
rect 83125 44779 83191 44780
rect 84213 44844 84279 44845
rect 84213 44780 84214 44844
rect 84278 44780 84279 44844
rect 84213 44779 84279 44780
rect 85440 44570 85500 45106
rect 81768 44510 82002 44570
rect 80467 42804 80533 42805
rect 80467 42740 80468 42804
rect 80532 42740 80533 42804
rect 80467 42739 80533 42740
rect 79547 41852 79613 41853
rect 79547 41788 79548 41852
rect 79612 41788 79613 41852
rect 79547 41787 79613 41788
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 43000
rect 81942 41853 82002 44510
rect 85438 44510 85500 44570
rect 86528 44570 86588 45106
rect 87616 44570 87676 45106
rect 88296 44570 88356 45106
rect 88704 44570 88764 45106
rect 90064 44570 90124 45106
rect 86528 44510 86602 44570
rect 87616 44510 87706 44570
rect 88296 44510 88442 44570
rect 88704 44510 88810 44570
rect 85438 43213 85498 44510
rect 85435 43212 85501 43213
rect 85435 43148 85436 43212
rect 85500 43148 85501 43212
rect 85435 43147 85501 43148
rect 81939 41852 82005 41853
rect 81939 41788 81940 41852
rect 82004 41788 82005 41852
rect 81939 41787 82005 41788
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 43000
rect 86542 42805 86602 44510
rect 87646 42805 87706 44510
rect 88382 42805 88442 44510
rect 88750 42805 88810 44510
rect 90038 44510 90124 44570
rect 90744 44570 90804 45106
rect 91288 44570 91348 45106
rect 92376 44570 92436 45106
rect 93464 44570 93524 45106
rect 90744 44510 90834 44570
rect 91288 44510 91386 44570
rect 92376 44510 92490 44570
rect 86539 42804 86605 42805
rect 86539 42740 86540 42804
rect 86604 42740 86605 42804
rect 86539 42739 86605 42740
rect 87643 42804 87709 42805
rect 87643 42740 87644 42804
rect 87708 42740 87709 42804
rect 87643 42739 87709 42740
rect 88379 42804 88445 42805
rect 88379 42740 88380 42804
rect 88444 42740 88445 42804
rect 88379 42739 88445 42740
rect 88747 42804 88813 42805
rect 88747 42740 88748 42804
rect 88812 42740 88813 42804
rect 88747 42739 88813 42740
rect 90038 41853 90098 44510
rect 90774 42805 90834 44510
rect 91326 42805 91386 44510
rect 92430 43213 92490 44510
rect 93350 44510 93524 44570
rect 93600 44570 93660 45106
rect 94552 44845 94612 45106
rect 94549 44844 94615 44845
rect 94549 44780 94550 44844
rect 94614 44780 94615 44844
rect 94549 44779 94615 44780
rect 95912 44570 95972 45106
rect 96048 44570 96108 45106
rect 97000 44845 97060 45106
rect 98088 44845 98148 45106
rect 96997 44844 97063 44845
rect 96997 44780 96998 44844
rect 97062 44780 97063 44844
rect 96997 44779 97063 44780
rect 98085 44844 98151 44845
rect 98085 44780 98086 44844
rect 98150 44780 98151 44844
rect 98085 44779 98151 44780
rect 98496 44570 98556 45106
rect 99448 44709 99508 45106
rect 100672 44842 100732 45106
rect 100672 44782 100770 44842
rect 100710 44709 100770 44782
rect 99445 44708 99511 44709
rect 99445 44644 99446 44708
rect 99510 44644 99511 44708
rect 99445 44643 99511 44644
rect 100707 44708 100773 44709
rect 100707 44644 100708 44708
rect 100772 44644 100773 44708
rect 100707 44643 100773 44644
rect 101080 44570 101140 45106
rect 101760 44709 101820 45106
rect 102848 44709 102908 45106
rect 101757 44708 101823 44709
rect 101757 44644 101758 44708
rect 101822 44644 101823 44708
rect 101757 44643 101823 44644
rect 102845 44708 102911 44709
rect 102845 44644 102846 44708
rect 102910 44644 102911 44708
rect 102845 44643 102911 44644
rect 93600 44510 93778 44570
rect 95912 44510 95986 44570
rect 96048 44510 96354 44570
rect 98496 44510 98562 44570
rect 92427 43212 92493 43213
rect 92427 43148 92428 43212
rect 92492 43148 92493 43212
rect 92427 43147 92493 43148
rect 90771 42804 90837 42805
rect 90771 42740 90772 42804
rect 90836 42740 90837 42804
rect 90771 42739 90837 42740
rect 91323 42804 91389 42805
rect 91323 42740 91324 42804
rect 91388 42740 91389 42804
rect 91323 42739 91389 42740
rect 90035 41852 90101 41853
rect 90035 41788 90036 41852
rect 90100 41788 90101 41852
rect 90035 41787 90101 41788
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 43000
rect 93350 42805 93410 44510
rect 93718 42805 93778 44510
rect 95926 43213 95986 44510
rect 95923 43212 95989 43213
rect 95923 43148 95924 43212
rect 95988 43148 95989 43212
rect 95923 43147 95989 43148
rect 93347 42804 93413 42805
rect 93347 42740 93348 42804
rect 93412 42740 93413 42804
rect 93347 42739 93413 42740
rect 93715 42804 93781 42805
rect 93715 42740 93716 42804
rect 93780 42740 93781 42804
rect 93715 42739 93781 42740
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 43000
rect 96294 42805 96354 44510
rect 96291 42804 96357 42805
rect 96291 42740 96292 42804
rect 96356 42740 96357 42804
rect 96291 42739 96357 42740
rect 98502 41989 98562 44510
rect 101078 44510 101140 44570
rect 103528 44570 103588 45106
rect 103936 44709 103996 45106
rect 103933 44708 103999 44709
rect 103933 44644 103934 44708
rect 103998 44644 103999 44708
rect 103933 44643 103999 44644
rect 105296 44570 105356 45106
rect 105976 44570 106036 45106
rect 103528 44510 103898 44570
rect 105296 44510 105370 44570
rect 101078 43349 101138 44510
rect 101075 43348 101141 43349
rect 101075 43284 101076 43348
rect 101140 43284 101141 43348
rect 101075 43283 101141 43284
rect 98499 41988 98565 41989
rect 98499 41924 98500 41988
rect 98564 41924 98565 41988
rect 98499 41923 98565 41924
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 43000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 43000
rect 103838 42125 103898 44510
rect 105310 43485 105370 44510
rect 105862 44510 106036 44570
rect 106384 44570 106444 45106
rect 107608 44570 107668 45106
rect 108288 44573 108348 45106
rect 106384 44510 106474 44570
rect 105307 43484 105373 43485
rect 105307 43420 105308 43484
rect 105372 43420 105373 43484
rect 105307 43419 105373 43420
rect 105862 42261 105922 44510
rect 106414 42805 106474 44510
rect 107518 44510 107668 44570
rect 108285 44572 108351 44573
rect 107518 42805 107578 44510
rect 108285 44508 108286 44572
rect 108350 44508 108351 44572
rect 108696 44570 108756 45106
rect 109784 44570 109844 45106
rect 108285 44507 108351 44508
rect 108622 44510 108756 44570
rect 109542 44510 109844 44570
rect 111008 44570 111068 45106
rect 111144 44570 111204 45106
rect 112232 44570 112292 45106
rect 113320 44573 113380 45106
rect 111008 44510 111074 44570
rect 111144 44510 111258 44570
rect 108622 42805 108682 44510
rect 106411 42804 106477 42805
rect 106411 42740 106412 42804
rect 106476 42740 106477 42804
rect 106411 42739 106477 42740
rect 107515 42804 107581 42805
rect 107515 42740 107516 42804
rect 107580 42740 107581 42804
rect 107515 42739 107581 42740
rect 108619 42804 108685 42805
rect 108619 42740 108620 42804
rect 108684 42740 108685 42804
rect 108619 42739 108685 42740
rect 109542 42261 109602 44510
rect 111014 43757 111074 44510
rect 111011 43756 111077 43757
rect 111011 43692 111012 43756
rect 111076 43692 111077 43756
rect 111011 43691 111077 43692
rect 105859 42260 105925 42261
rect 105859 42196 105860 42260
rect 105924 42196 105925 42260
rect 105859 42195 105925 42196
rect 109539 42260 109605 42261
rect 109539 42196 109540 42260
rect 109604 42196 109605 42260
rect 109539 42195 109605 42196
rect 103835 42124 103901 42125
rect 103835 42060 103836 42124
rect 103900 42060 103901 42124
rect 103835 42059 103901 42060
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 43000
rect 111198 42261 111258 44510
rect 112118 44510 112292 44570
rect 113317 44572 113383 44573
rect 112118 42805 112178 44510
rect 113317 44508 113318 44572
rect 113382 44508 113383 44572
rect 113592 44570 113652 45106
rect 114408 44570 114468 45106
rect 113317 44507 113383 44508
rect 113590 44510 113652 44570
rect 114326 44510 114468 44570
rect 115768 44570 115828 45106
rect 116040 44570 116100 45106
rect 116992 44570 117052 45106
rect 118080 44570 118140 45106
rect 118488 44570 118548 45106
rect 119168 44570 119228 45106
rect 120936 44570 120996 45106
rect 115768 44510 115858 44570
rect 113590 43890 113650 44510
rect 113222 43830 113650 43890
rect 113222 42805 113282 43830
rect 112115 42804 112181 42805
rect 112115 42740 112116 42804
rect 112180 42740 112181 42804
rect 112115 42739 112181 42740
rect 113219 42804 113285 42805
rect 113219 42740 113220 42804
rect 113284 42740 113285 42804
rect 113219 42739 113285 42740
rect 111195 42260 111261 42261
rect 111195 42196 111196 42260
rect 111260 42196 111261 42260
rect 111195 42195 111261 42196
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 43000
rect 114326 42805 114386 44510
rect 115798 42805 115858 44510
rect 115982 44510 116100 44570
rect 116902 44510 117052 44570
rect 118006 44510 118140 44570
rect 118374 44510 118548 44570
rect 119110 44510 119228 44570
rect 120766 44510 120996 44570
rect 123520 44570 123580 45106
rect 125968 44570 126028 45106
rect 123520 44510 123586 44570
rect 115982 43757 116042 44510
rect 115979 43756 116045 43757
rect 115979 43692 115980 43756
rect 116044 43692 116045 43756
rect 115979 43691 116045 43692
rect 116902 42805 116962 44510
rect 114323 42804 114389 42805
rect 114323 42740 114324 42804
rect 114388 42740 114389 42804
rect 114323 42739 114389 42740
rect 115795 42804 115861 42805
rect 115795 42740 115796 42804
rect 115860 42740 115861 42804
rect 115795 42739 115861 42740
rect 116899 42804 116965 42805
rect 116899 42740 116900 42804
rect 116964 42740 116965 42804
rect 116899 42739 116965 42740
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 43000
rect 118006 42397 118066 44510
rect 118374 42805 118434 44510
rect 119110 42805 119170 44510
rect 118371 42804 118437 42805
rect 118371 42740 118372 42804
rect 118436 42740 118437 42804
rect 118371 42739 118437 42740
rect 119107 42804 119173 42805
rect 119107 42740 119108 42804
rect 119172 42740 119173 42804
rect 119107 42739 119173 42740
rect 120766 42533 120826 44510
rect 123526 43621 123586 44510
rect 125918 44510 126028 44570
rect 128280 44570 128340 45106
rect 131000 44570 131060 45106
rect 128280 44510 128370 44570
rect 123523 43620 123589 43621
rect 123523 43556 123524 43620
rect 123588 43556 123589 43620
rect 123523 43555 123589 43556
rect 120763 42532 120829 42533
rect 120763 42468 120764 42532
rect 120828 42468 120829 42532
rect 120763 42467 120829 42468
rect 118003 42396 118069 42397
rect 118003 42332 118004 42396
rect 118068 42332 118069 42396
rect 118003 42331 118069 42332
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 43000
rect 125918 42669 125978 44510
rect 128310 43213 128370 44510
rect 130886 44510 131060 44570
rect 133448 44570 133508 45106
rect 135896 44570 135956 45106
rect 138480 44570 138540 45106
rect 140928 44573 140988 45106
rect 143512 44709 143572 45106
rect 145960 44709 146020 45106
rect 143509 44708 143575 44709
rect 143509 44644 143510 44708
rect 143574 44644 143575 44708
rect 143509 44643 143575 44644
rect 145957 44708 146023 44709
rect 145957 44644 145958 44708
rect 146022 44644 146023 44708
rect 145957 44643 146023 44644
rect 133448 44510 133522 44570
rect 135896 44510 136098 44570
rect 128307 43212 128373 43213
rect 128307 43148 128308 43212
rect 128372 43148 128373 43212
rect 128307 43147 128373 43148
rect 125915 42668 125981 42669
rect 125915 42604 125916 42668
rect 125980 42604 125981 42668
rect 125915 42603 125981 42604
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 43000
rect 130886 41581 130946 44510
rect 130883 41580 130949 41581
rect 130883 41516 130884 41580
rect 130948 41516 130949 41580
rect 130883 41515 130949 41516
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 43000
rect 133462 42805 133522 44510
rect 133459 42804 133525 42805
rect 133459 42740 133460 42804
rect 133524 42740 133525 42804
rect 133459 42739 133525 42740
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 43000
rect 136038 42805 136098 44510
rect 138430 44510 138540 44570
rect 140925 44572 140991 44573
rect 138430 44437 138490 44510
rect 140925 44508 140926 44572
rect 140990 44508 140991 44572
rect 148544 44570 148604 45106
rect 150992 44570 151052 45106
rect 153440 44570 153500 45106
rect 148544 44510 148610 44570
rect 140925 44507 140991 44508
rect 138427 44436 138493 44437
rect 138427 44372 138428 44436
rect 138492 44372 138493 44436
rect 138427 44371 138493 44372
rect 148550 43893 148610 44510
rect 150942 44510 151052 44570
rect 153334 44510 153500 44570
rect 155888 44570 155948 45106
rect 158472 44570 158532 45106
rect 160920 44570 160980 45106
rect 163368 44570 163428 45106
rect 165952 44570 166012 45106
rect 183224 44570 183284 45106
rect 155888 44510 155970 44570
rect 158472 44510 158546 44570
rect 150942 44029 151002 44510
rect 153334 44165 153394 44510
rect 153331 44164 153397 44165
rect 153331 44100 153332 44164
rect 153396 44100 153397 44164
rect 153331 44099 153397 44100
rect 150939 44028 151005 44029
rect 150939 43964 150940 44028
rect 151004 43964 151005 44028
rect 150939 43963 151005 43964
rect 148547 43892 148613 43893
rect 148547 43828 148548 43892
rect 148612 43828 148613 43892
rect 148547 43827 148613 43828
rect 136035 42804 136101 42805
rect 136035 42740 136036 42804
rect 136100 42740 136101 42804
rect 136035 42739 136101 42740
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 43000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 43000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 43000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 43000
rect 155910 42805 155970 44510
rect 158486 44165 158546 44510
rect 160878 44510 160980 44570
rect 163270 44510 163428 44570
rect 165846 44510 166012 44570
rect 183142 44510 183284 44570
rect 183360 44570 183420 45106
rect 183360 44510 183570 44570
rect 160878 44165 160938 44510
rect 158483 44164 158549 44165
rect 158483 44100 158484 44164
rect 158548 44100 158549 44164
rect 158483 44099 158549 44100
rect 160875 44164 160941 44165
rect 160875 44100 160876 44164
rect 160940 44100 160941 44164
rect 160875 44099 160941 44100
rect 155907 42804 155973 42805
rect 155907 42740 155908 42804
rect 155972 42740 155973 42804
rect 155907 42739 155973 42740
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 43000
rect 163270 41445 163330 44510
rect 163267 41444 163333 41445
rect 163267 41380 163268 41444
rect 163332 41380 163333 41444
rect 163267 41379 163333 41380
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 43000
rect 165846 42533 165906 44510
rect 165843 42532 165909 42533
rect 165843 42468 165844 42532
rect 165908 42468 165909 42532
rect 165843 42467 165909 42468
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 43000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 43000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 43000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 43000
rect 183142 42669 183202 44510
rect 183510 42805 183570 44510
rect 197862 43757 197922 492355
rect 198043 491740 198109 491741
rect 198043 491676 198044 491740
rect 198108 491676 198109 491740
rect 198043 491675 198109 491676
rect 198046 375325 198106 491675
rect 198411 491604 198477 491605
rect 198411 491540 198412 491604
rect 198476 491540 198477 491604
rect 198411 491539 198477 491540
rect 198043 375324 198109 375325
rect 198043 375260 198044 375324
rect 198108 375260 198109 375324
rect 198043 375259 198109 375260
rect 198414 44301 198474 491539
rect 198595 491332 198661 491333
rect 198595 491268 198596 491332
rect 198660 491268 198661 491332
rect 198595 491267 198661 491268
rect 198411 44300 198477 44301
rect 198411 44236 198412 44300
rect 198476 44236 198477 44300
rect 198411 44235 198477 44236
rect 198598 43893 198658 491267
rect 199794 489454 200414 493000
rect 201355 492284 201421 492285
rect 201355 492220 201356 492284
rect 201420 492220 201421 492284
rect 201355 492219 201421 492220
rect 202643 492284 202709 492285
rect 202643 492220 202644 492284
rect 202708 492220 202709 492284
rect 202643 492219 202709 492220
rect 201171 492148 201237 492149
rect 201171 492084 201172 492148
rect 201236 492084 201237 492148
rect 201171 492083 201237 492084
rect 200619 491468 200685 491469
rect 200619 491404 200620 491468
rect 200684 491404 200685 491468
rect 200619 491403 200685 491404
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199147 487796 199213 487797
rect 199147 487732 199148 487796
rect 199212 487732 199213 487796
rect 199147 487731 199213 487732
rect 198779 462908 198845 462909
rect 198779 462844 198780 462908
rect 198844 462844 198845 462908
rect 198779 462843 198845 462844
rect 198782 263397 198842 462843
rect 198963 461412 199029 461413
rect 198963 461348 198964 461412
rect 199028 461348 199029 461412
rect 198963 461347 199029 461348
rect 198966 350573 199026 461347
rect 199150 388517 199210 487731
rect 199331 463452 199397 463453
rect 199331 463388 199332 463452
rect 199396 463388 199397 463452
rect 199331 463387 199397 463388
rect 199147 388516 199213 388517
rect 199147 388452 199148 388516
rect 199212 388452 199213 388516
rect 199147 388451 199213 388452
rect 198963 350572 199029 350573
rect 198963 350508 198964 350572
rect 199028 350508 199029 350572
rect 198963 350507 199029 350508
rect 198779 263396 198845 263397
rect 198779 263332 198780 263396
rect 198844 263332 198845 263396
rect 198779 263331 198845 263332
rect 199334 262173 199394 463387
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199515 388516 199581 388517
rect 199515 388452 199516 388516
rect 199580 388452 199581 388516
rect 199515 388451 199581 388452
rect 199518 366349 199578 388451
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199515 366348 199581 366349
rect 199515 366284 199516 366348
rect 199580 366284 199581 366348
rect 199515 366283 199581 366284
rect 199794 362514 200414 380898
rect 199794 362278 199826 362514
rect 200062 362278 200146 362514
rect 200382 362278 200414 362514
rect 199794 362194 200414 362278
rect 199794 361958 199826 362194
rect 200062 361958 200146 362194
rect 200382 361958 200414 362194
rect 199794 345454 200414 361958
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199331 262172 199397 262173
rect 199331 262108 199332 262172
rect 199396 262108 199397 262172
rect 199331 262107 199397 262108
rect 199794 254514 200414 272898
rect 199794 254278 199826 254514
rect 200062 254278 200146 254514
rect 200382 254278 200414 254514
rect 199794 254194 200414 254278
rect 199794 253958 199826 254194
rect 200062 253958 200146 254194
rect 200382 253958 200414 254194
rect 199794 237454 200414 253958
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 146514 200414 164898
rect 199794 146278 199826 146514
rect 200062 146278 200146 146514
rect 200382 146278 200414 146514
rect 199794 146194 200414 146278
rect 199794 145958 199826 146194
rect 200062 145958 200146 146194
rect 200382 145958 200414 146194
rect 199794 129454 200414 145958
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 198595 43892 198661 43893
rect 198595 43828 198596 43892
rect 198660 43828 198661 43892
rect 198595 43827 198661 43828
rect 197859 43756 197925 43757
rect 197859 43692 197860 43756
rect 197924 43692 197925 43756
rect 197859 43691 197925 43692
rect 183507 42804 183573 42805
rect 183507 42740 183508 42804
rect 183572 42740 183573 42804
rect 183507 42739 183573 42740
rect 183139 42668 183205 42669
rect 183139 42604 183140 42668
rect 183204 42604 183205 42668
rect 183139 42603 183205 42604
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 43000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 43000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 43000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 56898
rect 200622 43349 200682 491403
rect 200803 479500 200869 479501
rect 200803 479436 200804 479500
rect 200868 479436 200869 479500
rect 200803 479435 200869 479436
rect 200619 43348 200685 43349
rect 200619 43284 200620 43348
rect 200684 43284 200685 43348
rect 200619 43283 200685 43284
rect 200806 41717 200866 479435
rect 201174 44437 201234 492083
rect 201171 44436 201237 44437
rect 201171 44372 201172 44436
rect 201236 44372 201237 44436
rect 201171 44371 201237 44372
rect 201358 43621 201418 492219
rect 202275 467124 202341 467125
rect 202275 467060 202276 467124
rect 202340 467060 202341 467124
rect 202275 467059 202341 467060
rect 202091 463180 202157 463181
rect 202091 463116 202092 463180
rect 202156 463116 202157 463180
rect 202091 463115 202157 463116
rect 202094 55045 202154 463115
rect 202278 152149 202338 467059
rect 202459 461684 202525 461685
rect 202459 461620 202460 461684
rect 202524 461620 202525 461684
rect 202459 461619 202525 461620
rect 202462 154461 202522 461619
rect 202459 154460 202525 154461
rect 202459 154396 202460 154460
rect 202524 154396 202525 154460
rect 202459 154395 202525 154396
rect 202275 152148 202341 152149
rect 202275 152084 202276 152148
rect 202340 152084 202341 152148
rect 202275 152083 202341 152084
rect 202091 55044 202157 55045
rect 202091 54980 202092 55044
rect 202156 54980 202157 55044
rect 202091 54979 202157 54980
rect 202646 44029 202706 492219
rect 203514 476114 204134 493000
rect 206875 492148 206941 492149
rect 206875 492084 206876 492148
rect 206940 492084 206941 492148
rect 206875 492083 206941 492084
rect 204851 492012 204917 492013
rect 204851 491948 204852 492012
rect 204916 491948 204917 492012
rect 204851 491947 204917 491948
rect 203514 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 204134 476114
rect 203514 475794 204134 475878
rect 203514 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 204134 475794
rect 203195 461548 203261 461549
rect 203195 461484 203196 461548
rect 203260 461484 203261 461548
rect 203195 461483 203261 461484
rect 203011 460460 203077 460461
rect 203011 460396 203012 460460
rect 203076 460396 203077 460460
rect 203011 460395 203077 460396
rect 203014 154189 203074 460395
rect 203011 154188 203077 154189
rect 203011 154124 203012 154188
rect 203076 154124 203077 154188
rect 203011 154123 203077 154124
rect 203198 152557 203258 461483
rect 203514 457174 204134 475558
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 366234 204134 384618
rect 203514 365998 203546 366234
rect 203782 365998 203866 366234
rect 204102 365998 204134 366234
rect 203514 365914 204134 365998
rect 203514 365678 203546 365914
rect 203782 365678 203866 365914
rect 204102 365678 204134 365914
rect 203514 349174 204134 365678
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203195 152556 203261 152557
rect 203195 152492 203196 152556
rect 203260 152492 203261 152556
rect 203195 152491 203261 152492
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 202643 44028 202709 44029
rect 202643 43964 202644 44028
rect 202708 43964 202709 44028
rect 202643 43963 202709 43964
rect 201355 43620 201421 43621
rect 201355 43556 201356 43620
rect 201420 43556 201421 43620
rect 201355 43555 201421 43556
rect 200803 41716 200869 41717
rect 200803 41652 200804 41716
rect 200868 41652 200869 41716
rect 200803 41651 200869 41652
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 60618
rect 204854 43485 204914 491947
rect 205035 491876 205101 491877
rect 205035 491812 205036 491876
rect 205100 491812 205101 491876
rect 205035 491811 205101 491812
rect 205038 44709 205098 491811
rect 205219 491740 205285 491741
rect 205219 491676 205220 491740
rect 205284 491676 205285 491740
rect 205219 491675 205285 491676
rect 205035 44708 205101 44709
rect 205035 44644 205036 44708
rect 205100 44644 205101 44708
rect 205035 44643 205101 44644
rect 205222 44573 205282 491675
rect 206507 489156 206573 489157
rect 206507 489092 206508 489156
rect 206572 489092 206573 489156
rect 206507 489091 206573 489092
rect 206139 483716 206205 483717
rect 206139 483652 206140 483716
rect 206204 483652 206205 483716
rect 206139 483651 206205 483652
rect 205403 459372 205469 459373
rect 205403 459308 205404 459372
rect 205468 459308 205469 459372
rect 205403 459307 205469 459308
rect 205406 151741 205466 459307
rect 205403 151740 205469 151741
rect 205403 151676 205404 151740
rect 205468 151676 205469 151740
rect 205403 151675 205469 151676
rect 205219 44572 205285 44573
rect 205219 44508 205220 44572
rect 205284 44508 205285 44572
rect 205219 44507 205285 44508
rect 204851 43484 204917 43485
rect 204851 43420 204852 43484
rect 204916 43420 204917 43484
rect 204851 43419 204917 43420
rect 206142 42261 206202 483651
rect 206323 478140 206389 478141
rect 206323 478076 206324 478140
rect 206388 478076 206389 478140
rect 206323 478075 206389 478076
rect 206326 53141 206386 478075
rect 206510 152965 206570 489091
rect 206507 152964 206573 152965
rect 206507 152900 206508 152964
rect 206572 152900 206573 152964
rect 206507 152899 206573 152900
rect 206323 53140 206389 53141
rect 206323 53076 206324 53140
rect 206388 53076 206389 53140
rect 206323 53075 206389 53076
rect 206878 44165 206938 492083
rect 207234 477954 207854 493000
rect 210371 486572 210437 486573
rect 210371 486508 210372 486572
rect 210436 486508 210437 486572
rect 210371 486507 210437 486508
rect 208899 486436 208965 486437
rect 208899 486372 208900 486436
rect 208964 486372 208965 486436
rect 208899 486371 208965 486372
rect 207234 477718 207266 477954
rect 207502 477718 207586 477954
rect 207822 477718 207854 477954
rect 207234 477634 207854 477718
rect 207234 477398 207266 477634
rect 207502 477398 207586 477634
rect 207822 477398 207854 477634
rect 207234 460894 207854 477398
rect 208347 476780 208413 476781
rect 208347 476716 208348 476780
rect 208412 476716 208413 476780
rect 208347 476715 208413 476716
rect 207979 472564 208045 472565
rect 207979 472500 207980 472564
rect 208044 472500 208045 472564
rect 207979 472499 208045 472500
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 206875 44164 206941 44165
rect 206875 44100 206876 44164
rect 206940 44100 206941 44164
rect 206875 44099 206941 44100
rect 206139 42260 206205 42261
rect 206139 42196 206140 42260
rect 206204 42196 206205 42260
rect 206139 42195 206205 42196
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 64338
rect 207982 42125 208042 472499
rect 208163 459236 208229 459237
rect 208163 459172 208164 459236
rect 208228 459172 208229 459236
rect 208163 459171 208229 459172
rect 208166 154325 208226 459171
rect 208350 372605 208410 476715
rect 208531 474060 208597 474061
rect 208531 473996 208532 474060
rect 208596 473996 208597 474060
rect 208531 473995 208597 473996
rect 208347 372604 208413 372605
rect 208347 372540 208348 372604
rect 208412 372540 208413 372604
rect 208347 372539 208413 372540
rect 208534 371245 208594 473995
rect 208531 371244 208597 371245
rect 208531 371180 208532 371244
rect 208596 371180 208597 371244
rect 208531 371179 208597 371180
rect 208163 154324 208229 154325
rect 208163 154260 208164 154324
rect 208228 154260 208229 154324
rect 208163 154259 208229 154260
rect 207979 42124 208045 42125
rect 207979 42060 207980 42124
rect 208044 42060 208045 42124
rect 207979 42059 208045 42060
rect 208902 41989 208962 486371
rect 209819 460324 209885 460325
rect 209819 460260 209820 460324
rect 209884 460260 209885 460324
rect 209819 460259 209885 460260
rect 209822 369205 209882 460259
rect 209819 369204 209885 369205
rect 209819 369140 209820 369204
rect 209884 369140 209885 369204
rect 209819 369139 209885 369140
rect 210374 42533 210434 486507
rect 210954 464614 211574 493000
rect 213315 492556 213381 492557
rect 213315 492492 213316 492556
rect 213380 492492 213381 492556
rect 213315 492491 213381 492492
rect 217363 492556 217429 492557
rect 217363 492492 217364 492556
rect 217428 492492 217429 492556
rect 217363 492491 217429 492492
rect 211659 491604 211725 491605
rect 211659 491540 211660 491604
rect 211724 491540 211725 491604
rect 211659 491539 211725 491540
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 211662 369205 211722 491539
rect 212579 468484 212645 468485
rect 212579 468420 212580 468484
rect 212644 468420 212645 468484
rect 212579 468419 212645 468420
rect 212582 383670 212642 468419
rect 213131 458964 213197 458965
rect 213131 458900 213132 458964
rect 213196 458900 213197 458964
rect 213131 458899 213197 458900
rect 212582 383610 212826 383670
rect 212766 373829 212826 383610
rect 212763 373828 212829 373829
rect 212763 373764 212764 373828
rect 212828 373764 212829 373828
rect 212763 373763 212829 373764
rect 211659 369204 211725 369205
rect 211659 369140 211660 369204
rect 211724 369140 211725 369204
rect 211659 369139 211725 369140
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 213134 153917 213194 458899
rect 213318 369205 213378 492491
rect 213867 490516 213933 490517
rect 213867 490452 213868 490516
rect 213932 490452 213933 490516
rect 213867 490451 213933 490452
rect 213870 369205 213930 490451
rect 217179 478276 217245 478277
rect 217179 478212 217180 478276
rect 217244 478212 217245 478276
rect 217179 478211 217245 478212
rect 214419 475420 214485 475421
rect 214419 475356 214420 475420
rect 214484 475356 214485 475420
rect 214419 475355 214485 475356
rect 213315 369204 213381 369205
rect 213315 369140 213316 369204
rect 213380 369140 213381 369204
rect 213315 369139 213381 369140
rect 213867 369204 213933 369205
rect 213867 369140 213868 369204
rect 213932 369140 213933 369204
rect 213867 369139 213933 369140
rect 213131 153916 213197 153917
rect 213131 153852 213132 153916
rect 213196 153852 213197 153916
rect 213131 153851 213197 153852
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210371 42532 210437 42533
rect 210371 42468 210372 42532
rect 210436 42468 210437 42532
rect 210371 42467 210437 42468
rect 208899 41988 208965 41989
rect 208899 41924 208900 41988
rect 208964 41924 208965 41988
rect 208899 41923 208965 41924
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 68058
rect 214422 42397 214482 475355
rect 214603 469980 214669 469981
rect 214603 469916 214604 469980
rect 214668 469916 214669 469980
rect 214603 469915 214669 469916
rect 214606 152693 214666 469915
rect 215339 469844 215405 469845
rect 215339 469780 215340 469844
rect 215404 469780 215405 469844
rect 215339 469779 215405 469780
rect 215342 369885 215402 469779
rect 216075 463044 216141 463045
rect 216075 462980 216076 463044
rect 216140 462980 216141 463044
rect 216075 462979 216141 462980
rect 215891 458828 215957 458829
rect 215891 458764 215892 458828
rect 215956 458764 215957 458828
rect 215891 458763 215957 458764
rect 215339 369884 215405 369885
rect 215339 369820 215340 369884
rect 215404 369820 215405 369884
rect 215339 369819 215405 369820
rect 214603 152692 214669 152693
rect 214603 152628 214604 152692
rect 214668 152628 214669 152692
rect 214603 152627 214669 152628
rect 215894 42669 215954 458763
rect 216078 154053 216138 462979
rect 216995 459644 217061 459645
rect 216995 459580 216996 459644
rect 217060 459580 217061 459644
rect 216995 459579 217061 459580
rect 216627 372876 216693 372877
rect 216627 372812 216628 372876
rect 216692 372812 216693 372876
rect 216627 372811 216693 372812
rect 216630 370565 216690 372811
rect 216811 372740 216877 372741
rect 216811 372676 216812 372740
rect 216876 372676 216877 372740
rect 216811 372675 216877 372676
rect 216814 371109 216874 372675
rect 216998 371653 217058 459579
rect 216995 371652 217061 371653
rect 216995 371588 216996 371652
rect 217060 371588 217061 371652
rect 216995 371587 217061 371588
rect 216811 371108 216877 371109
rect 216811 371044 216812 371108
rect 216876 371044 216877 371108
rect 216811 371043 216877 371044
rect 216627 370564 216693 370565
rect 216627 370500 216628 370564
rect 216692 370500 216693 370564
rect 216627 370499 216693 370500
rect 217182 263125 217242 478211
rect 217366 373829 217426 492491
rect 217547 492420 217613 492421
rect 217547 492356 217548 492420
rect 217612 492356 217613 492420
rect 217547 492355 217613 492356
rect 217550 374237 217610 492355
rect 217794 471454 218414 493000
rect 219939 492556 220005 492557
rect 219939 492492 219940 492556
rect 220004 492492 220005 492556
rect 219939 492491 220005 492492
rect 219203 491876 219269 491877
rect 219203 491812 219204 491876
rect 219268 491812 219269 491876
rect 219203 491811 219269 491812
rect 219019 475556 219085 475557
rect 219019 475492 219020 475556
rect 219084 475492 219085 475556
rect 219019 475491 219085 475492
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 460308 218414 470898
rect 218651 460188 218717 460189
rect 218651 460124 218652 460188
rect 218716 460124 218717 460188
rect 218651 460123 218717 460124
rect 217547 374236 217613 374237
rect 217547 374172 217548 374236
rect 217612 374172 217613 374236
rect 217547 374171 217613 374172
rect 217363 373828 217429 373829
rect 217363 373764 217364 373828
rect 217428 373764 217429 373828
rect 217363 373763 217429 373764
rect 217366 373421 217426 373763
rect 217363 373420 217429 373421
rect 217363 373356 217364 373420
rect 217428 373356 217429 373420
rect 217363 373355 217429 373356
rect 217794 363454 218414 373000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 350308 218414 362898
rect 217179 263124 217245 263125
rect 217179 263060 217180 263124
rect 217244 263060 217245 263124
rect 217179 263059 217245 263060
rect 217794 255454 218414 263000
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 240308 218414 254898
rect 217547 240276 217613 240277
rect 217547 240212 217548 240276
rect 217612 240212 217613 240276
rect 217547 240211 217613 240212
rect 216075 154052 216141 154053
rect 216075 153988 216076 154052
rect 216140 153988 216141 154052
rect 216075 153987 216141 153988
rect 217550 130933 217610 240211
rect 218654 153101 218714 460123
rect 218835 350436 218901 350437
rect 218835 350372 218836 350436
rect 218900 350372 218901 350436
rect 218835 350371 218901 350372
rect 218651 153100 218717 153101
rect 218651 153036 218652 153100
rect 218716 153036 218717 153100
rect 218651 153035 218717 153036
rect 217794 147454 218414 153000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217547 130932 217613 130933
rect 217547 130868 217548 130932
rect 217612 130868 217613 130932
rect 217547 130867 217613 130868
rect 215891 42668 215957 42669
rect 215891 42604 215892 42668
rect 215956 42604 215957 42668
rect 215891 42603 215957 42604
rect 214419 42396 214485 42397
rect 214419 42332 214420 42396
rect 214484 42332 214485 42396
rect 214419 42331 214485 42332
rect 217550 39949 217610 130867
rect 217794 130308 218414 146898
rect 218838 44845 218898 350371
rect 219022 263669 219082 475491
rect 219019 263668 219085 263669
rect 219019 263604 219020 263668
rect 219084 263604 219085 263668
rect 219019 263603 219085 263604
rect 219206 44845 219266 491811
rect 218835 44844 218901 44845
rect 218835 44780 218836 44844
rect 218900 44780 218901 44844
rect 218835 44779 218901 44780
rect 219203 44844 219269 44845
rect 219203 44780 219204 44844
rect 219268 44780 219269 44844
rect 219203 44779 219269 44780
rect 217547 39948 217613 39949
rect 217547 39884 217548 39948
rect 217612 39884 217613 39948
rect 217547 39883 217613 39884
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 43000
rect 219942 41309 220002 492491
rect 221514 475174 222134 493000
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 460308 222134 474618
rect 225234 478894 225854 493000
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 460308 225854 478338
rect 228954 482614 229574 493000
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 460308 229574 482058
rect 235794 489454 236414 493000
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 460308 236414 488898
rect 239514 476114 240134 493000
rect 239514 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 240134 476114
rect 239514 475794 240134 475878
rect 239514 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 240134 475794
rect 239514 460308 240134 475558
rect 243234 477954 243854 493000
rect 243234 477718 243266 477954
rect 243502 477718 243586 477954
rect 243822 477718 243854 477954
rect 243234 477634 243854 477718
rect 243234 477398 243266 477634
rect 243502 477398 243586 477634
rect 243822 477398 243854 477634
rect 243234 460308 243854 477398
rect 246954 464614 247574 493000
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 460308 247574 464058
rect 253794 471454 254414 493000
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 460308 254414 470898
rect 257514 475174 258134 493000
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 460308 258134 474618
rect 261234 478894 261854 493000
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 460308 261854 478338
rect 264954 482614 265574 493000
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 460308 265574 482058
rect 271794 489454 272414 493000
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 460308 272414 488898
rect 275514 476114 276134 493000
rect 275514 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 275514 475794 276134 475878
rect 275514 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 275514 460308 276134 475558
rect 279234 477954 279854 493000
rect 279234 477718 279266 477954
rect 279502 477718 279586 477954
rect 279822 477718 279854 477954
rect 279234 477634 279854 477718
rect 279234 477398 279266 477634
rect 279502 477398 279586 477634
rect 279822 477398 279854 477634
rect 279234 460308 279854 477398
rect 282954 464614 283574 493000
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 460308 283574 464058
rect 289794 471454 290414 493000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 460308 290414 470898
rect 293514 475174 294134 493000
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 460308 294134 474618
rect 297234 478894 297854 493000
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 460308 297854 478338
rect 300954 482614 301574 493000
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 460308 301574 482058
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 460308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 460308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 648033 319574 680058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 648033 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 648033 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 648033 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 648033 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 648033 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 648033 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 648033 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 648033 355574 680058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 648033 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 648033 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 648033 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 648033 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 648033 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 648033 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 648033 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 648033 391574 680058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 648033 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 648033 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 648033 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 648033 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 648033 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 648033 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 648033 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 648033 427574 680058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 339568 633454 339888 633486
rect 339568 633218 339610 633454
rect 339846 633218 339888 633454
rect 339568 633134 339888 633218
rect 339568 632898 339610 633134
rect 339846 632898 339888 633134
rect 339568 632866 339888 632898
rect 370288 633454 370608 633486
rect 370288 633218 370330 633454
rect 370566 633218 370608 633454
rect 370288 633134 370608 633218
rect 370288 632898 370330 633134
rect 370566 632898 370608 633134
rect 370288 632866 370608 632898
rect 401008 633454 401328 633486
rect 401008 633218 401050 633454
rect 401286 633218 401328 633454
rect 401008 633134 401328 633218
rect 401008 632898 401050 633134
rect 401286 632898 401328 633134
rect 401008 632866 401328 632898
rect 430619 622164 430685 622165
rect 430619 622100 430620 622164
rect 430684 622100 430685 622164
rect 430619 622099 430685 622100
rect 324208 615454 324528 615486
rect 324208 615218 324250 615454
rect 324486 615218 324528 615454
rect 324208 615134 324528 615218
rect 324208 614898 324250 615134
rect 324486 614898 324528 615134
rect 324208 614866 324528 614898
rect 354928 615454 355248 615486
rect 354928 615218 354970 615454
rect 355206 615218 355248 615454
rect 354928 615134 355248 615218
rect 354928 614898 354970 615134
rect 355206 614898 355248 615134
rect 354928 614866 355248 614898
rect 385648 615454 385968 615486
rect 385648 615218 385690 615454
rect 385926 615218 385968 615454
rect 385648 615134 385968 615218
rect 385648 614898 385690 615134
rect 385926 614898 385968 615134
rect 385648 614866 385968 614898
rect 416368 615454 416688 615486
rect 416368 615218 416410 615454
rect 416646 615218 416688 615454
rect 416368 615134 416688 615218
rect 416368 614898 416410 615134
rect 416646 614898 416688 615134
rect 416368 614866 416688 614898
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 339568 597454 339888 597486
rect 339568 597218 339610 597454
rect 339846 597218 339888 597454
rect 339568 597134 339888 597218
rect 339568 596898 339610 597134
rect 339846 596898 339888 597134
rect 339568 596866 339888 596898
rect 370288 597454 370608 597486
rect 370288 597218 370330 597454
rect 370566 597218 370608 597454
rect 370288 597134 370608 597218
rect 370288 596898 370330 597134
rect 370566 596898 370608 597134
rect 370288 596866 370608 596898
rect 401008 597454 401328 597486
rect 401008 597218 401050 597454
rect 401286 597218 401328 597454
rect 401008 597134 401328 597218
rect 401008 596898 401050 597134
rect 401286 596898 401328 597134
rect 401008 596866 401328 596898
rect 324208 579454 324528 579486
rect 324208 579218 324250 579454
rect 324486 579218 324528 579454
rect 324208 579134 324528 579218
rect 324208 578898 324250 579134
rect 324486 578898 324528 579134
rect 324208 578866 324528 578898
rect 354928 579454 355248 579486
rect 354928 579218 354970 579454
rect 355206 579218 355248 579454
rect 354928 579134 355248 579218
rect 354928 578898 354970 579134
rect 355206 578898 355248 579134
rect 354928 578866 355248 578898
rect 385648 579454 385968 579486
rect 385648 579218 385690 579454
rect 385926 579218 385968 579454
rect 385648 579134 385968 579218
rect 385648 578898 385690 579134
rect 385926 578898 385968 579134
rect 385648 578866 385968 578898
rect 416368 579454 416688 579486
rect 416368 579218 416410 579454
rect 416646 579218 416688 579454
rect 416368 579134 416688 579218
rect 416368 578898 416410 579134
rect 416646 578898 416688 579134
rect 416368 578866 416688 578898
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 339568 561454 339888 561486
rect 339568 561218 339610 561454
rect 339846 561218 339888 561454
rect 339568 561134 339888 561218
rect 339568 560898 339610 561134
rect 339846 560898 339888 561134
rect 339568 560866 339888 560898
rect 370288 561454 370608 561486
rect 370288 561218 370330 561454
rect 370566 561218 370608 561454
rect 370288 561134 370608 561218
rect 370288 560898 370330 561134
rect 370566 560898 370608 561134
rect 370288 560866 370608 560898
rect 401008 561454 401328 561486
rect 401008 561218 401050 561454
rect 401286 561218 401328 561454
rect 401008 561134 401328 561218
rect 401008 560898 401050 561134
rect 401286 560898 401328 561134
rect 401008 560866 401328 560898
rect 324208 543454 324528 543486
rect 324208 543218 324250 543454
rect 324486 543218 324528 543454
rect 324208 543134 324528 543218
rect 324208 542898 324250 543134
rect 324486 542898 324528 543134
rect 324208 542866 324528 542898
rect 354928 543454 355248 543486
rect 354928 543218 354970 543454
rect 355206 543218 355248 543454
rect 354928 543134 355248 543218
rect 354928 542898 354970 543134
rect 355206 542898 355248 543134
rect 354928 542866 355248 542898
rect 385648 543454 385968 543486
rect 385648 543218 385690 543454
rect 385926 543218 385968 543454
rect 385648 543134 385968 543218
rect 385648 542898 385690 543134
rect 385926 542898 385968 543134
rect 385648 542866 385968 542898
rect 416368 543454 416688 543486
rect 416368 543218 416410 543454
rect 416646 543218 416688 543454
rect 416368 543134 416688 543218
rect 416368 542898 416410 543134
rect 416646 542898 416688 543134
rect 416368 542866 416688 542898
rect 430622 535533 430682 622099
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 430803 607884 430869 607885
rect 430803 607820 430804 607884
rect 430868 607820 430869 607884
rect 430803 607819 430869 607820
rect 430619 535532 430685 535533
rect 430619 535468 430620 535532
rect 430684 535468 430685 535532
rect 430619 535467 430685 535468
rect 430806 535397 430866 607819
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 430803 535396 430869 535397
rect 430803 535332 430804 535396
rect 430868 535332 430869 535396
rect 430803 535331 430869 535332
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460308 315854 496338
rect 318954 500614 319574 533000
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 460308 319574 464058
rect 325794 507454 326414 533000
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 460308 326414 470898
rect 329514 511174 330134 533000
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 460308 330134 474618
rect 333234 514894 333854 533000
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 460308 333854 478338
rect 336954 518614 337574 533000
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 460308 337574 482058
rect 343794 525454 344414 533000
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 339723 461276 339789 461277
rect 339723 461212 339724 461276
rect 339788 461212 339789 461276
rect 339723 461211 339789 461212
rect 338251 461004 338317 461005
rect 338251 460940 338252 461004
rect 338316 460950 338317 461004
rect 338316 460940 338498 460950
rect 338251 460939 338498 460940
rect 338254 460890 338498 460939
rect 338438 458690 338498 460890
rect 339726 458690 339786 461211
rect 343794 460308 344414 488898
rect 347514 529174 348134 533000
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 460308 348134 492618
rect 351234 532894 351854 533000
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350947 461004 351013 461005
rect 350947 460940 350948 461004
rect 351012 460940 351013 461004
rect 350947 460939 351013 460940
rect 350950 458690 351010 460939
rect 351234 460308 351854 496338
rect 354954 500614 355574 533000
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 361794 507454 362414 533000
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 357939 492556 358005 492557
rect 357939 492492 357940 492556
rect 358004 492492 358005 492556
rect 357939 492491 358005 492492
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 460308 355574 464058
rect 338438 458630 338524 458690
rect 338464 458202 338524 458630
rect 339688 458630 339786 458690
rect 350840 458630 351010 458690
rect 339688 458202 339748 458630
rect 350840 458202 350900 458630
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 220952 399454 221300 399486
rect 220952 399218 221008 399454
rect 221244 399218 221300 399454
rect 220952 399134 221300 399218
rect 220952 398898 221008 399134
rect 221244 398898 221300 399134
rect 220952 398866 221300 398898
rect 355320 399454 355668 399486
rect 355320 399218 355376 399454
rect 355612 399218 355668 399454
rect 355320 399134 355668 399218
rect 355320 398898 355376 399134
rect 355612 398898 355668 399134
rect 355320 398866 355668 398898
rect 220272 381454 220620 381486
rect 220272 381218 220328 381454
rect 220564 381218 220620 381454
rect 220272 381134 220620 381218
rect 220272 380898 220328 381134
rect 220564 380898 220620 381134
rect 220272 380866 220620 380898
rect 356000 381454 356348 381486
rect 356000 381218 356056 381454
rect 356292 381218 356348 381454
rect 356000 381134 356348 381218
rect 356000 380898 356056 381134
rect 356292 380898 356348 381134
rect 356000 380866 356348 380898
rect 263731 375052 263797 375053
rect 235950 374990 236086 375050
rect 236502 374990 237174 375050
rect 238158 374990 238262 375050
rect 239078 374990 239622 375050
rect 235950 373285 236010 374990
rect 236502 373693 236562 374990
rect 236499 373692 236565 373693
rect 236499 373628 236500 373692
rect 236564 373628 236565 373692
rect 236499 373627 236565 373628
rect 235947 373284 236013 373285
rect 235947 373220 235948 373284
rect 236012 373220 236013 373284
rect 235947 373219 236013 373220
rect 221514 367174 222134 373000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 350308 222134 366618
rect 225234 370894 225854 373000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 350308 225854 370338
rect 228954 357554 229574 373000
rect 228954 357318 228986 357554
rect 229222 357318 229306 357554
rect 229542 357318 229574 357554
rect 228954 357234 229574 357318
rect 228954 356998 228986 357234
rect 229222 356998 229306 357234
rect 229542 356998 229574 357234
rect 228954 350308 229574 356998
rect 235794 362514 236414 373000
rect 238158 372605 238218 374990
rect 239078 372605 239138 374990
rect 238155 372604 238221 372605
rect 238155 372540 238156 372604
rect 238220 372540 238221 372604
rect 238155 372539 238221 372540
rect 239075 372604 239141 372605
rect 239075 372540 239076 372604
rect 239140 372540 239141 372604
rect 239075 372539 239141 372540
rect 235794 362278 235826 362514
rect 236062 362278 236146 362514
rect 236382 362278 236414 362514
rect 235794 362194 236414 362278
rect 235794 361958 235826 362194
rect 236062 361958 236146 362194
rect 236382 361958 236414 362194
rect 235794 350308 236414 361958
rect 239514 366234 240134 373000
rect 240550 372061 240610 375050
rect 241654 374990 241798 375050
rect 242942 374990 243158 375050
rect 240547 372060 240613 372061
rect 240547 371996 240548 372060
rect 240612 371996 240613 372060
rect 240547 371995 240613 371996
rect 241654 371925 241714 374990
rect 242942 373693 243002 374990
rect 244230 374509 244290 375050
rect 244782 374990 245470 375050
rect 245886 374990 246558 375050
rect 247174 374990 247646 375050
rect 247910 374990 248326 375050
rect 244227 374508 244293 374509
rect 244227 374444 244228 374508
rect 244292 374444 244293 374508
rect 244227 374443 244293 374444
rect 242939 373692 243005 373693
rect 242939 373628 242940 373692
rect 243004 373628 243005 373692
rect 242939 373627 243005 373628
rect 241651 371924 241717 371925
rect 241651 371860 241652 371924
rect 241716 371860 241717 371924
rect 241651 371859 241717 371860
rect 241654 371653 241714 371859
rect 241651 371652 241717 371653
rect 241651 371588 241652 371652
rect 241716 371588 241717 371652
rect 241651 371587 241717 371588
rect 239514 365998 239546 366234
rect 239782 365998 239866 366234
rect 240102 365998 240134 366234
rect 239514 365914 240134 365998
rect 239514 365678 239546 365914
rect 239782 365678 239866 365914
rect 240102 365678 240134 365914
rect 239514 350308 240134 365678
rect 243234 352894 243854 373000
rect 244782 372605 244842 374990
rect 244779 372604 244845 372605
rect 244779 372540 244780 372604
rect 244844 372540 244845 372604
rect 244779 372539 244845 372540
rect 245886 371925 245946 374990
rect 247174 373149 247234 374990
rect 247171 373148 247237 373149
rect 247171 373084 247172 373148
rect 247236 373084 247237 373148
rect 247171 373083 247237 373084
rect 245883 371924 245949 371925
rect 245883 371860 245884 371924
rect 245948 371860 245949 371924
rect 245883 371859 245949 371860
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 350308 243854 352338
rect 246954 356614 247574 373000
rect 247910 371517 247970 374990
rect 248704 374509 248764 375020
rect 250064 374509 250124 375020
rect 250302 374990 250774 375050
rect 251222 374990 251318 375050
rect 251958 374990 252406 375050
rect 252878 374990 253494 375050
rect 248701 374508 248767 374509
rect 248701 374444 248702 374508
rect 248766 374444 248767 374508
rect 248701 374443 248767 374444
rect 250061 374508 250127 374509
rect 250061 374444 250062 374508
rect 250126 374444 250127 374508
rect 250061 374443 250127 374444
rect 250302 371517 250362 374990
rect 251222 371653 251282 374990
rect 251958 372605 252018 374990
rect 252878 372605 252938 374990
rect 251955 372604 252021 372605
rect 251955 372540 251956 372604
rect 252020 372540 252021 372604
rect 251955 372539 252021 372540
rect 252875 372604 252941 372605
rect 252875 372540 252876 372604
rect 252940 372540 252941 372604
rect 252875 372539 252941 372540
rect 251219 371652 251285 371653
rect 251219 371588 251220 371652
rect 251284 371588 251285 371652
rect 251219 371587 251285 371588
rect 253614 371517 253674 375050
rect 253982 374990 254582 375050
rect 255454 374990 255942 375050
rect 256078 374990 256250 375050
rect 253982 373285 254042 374990
rect 255454 373285 255514 374990
rect 253979 373284 254045 373285
rect 253979 373220 253980 373284
rect 254044 373220 254045 373284
rect 253979 373219 254045 373220
rect 255451 373284 255517 373285
rect 255451 373220 255452 373284
rect 255516 373220 255517 373284
rect 255451 373219 255517 373220
rect 247907 371516 247973 371517
rect 247907 371452 247908 371516
rect 247972 371452 247973 371516
rect 247907 371451 247973 371452
rect 250299 371516 250365 371517
rect 250299 371452 250300 371516
rect 250364 371452 250365 371516
rect 250299 371451 250365 371452
rect 253611 371516 253677 371517
rect 253611 371452 253612 371516
rect 253676 371452 253677 371516
rect 253611 371451 253677 371452
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 350308 247574 356058
rect 253794 363454 254414 373000
rect 256190 371517 256250 374990
rect 256742 374990 257030 375050
rect 258118 374990 258274 375050
rect 256742 373285 256802 374990
rect 258214 374010 258274 374990
rect 258030 373965 258274 374010
rect 258027 373964 258274 373965
rect 258027 373900 258028 373964
rect 258092 373950 258274 373964
rect 258398 374990 258526 375050
rect 259478 374990 259562 375050
rect 258092 373900 258093 373950
rect 258027 373899 258093 373900
rect 256739 373284 256805 373285
rect 256739 373220 256740 373284
rect 256804 373220 256805 373284
rect 256739 373219 256805 373220
rect 256187 371516 256253 371517
rect 256187 371452 256188 371516
rect 256252 371452 256253 371516
rect 256187 371451 256253 371452
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 350308 254414 362898
rect 257514 367174 258134 373000
rect 258398 371653 258458 374990
rect 259502 372605 259562 374990
rect 260054 374990 260702 375050
rect 260974 374990 261110 375050
rect 261342 374990 261790 375050
rect 262262 374990 262878 375050
rect 260054 372605 260114 374990
rect 259499 372604 259565 372605
rect 259499 372540 259500 372604
rect 259564 372540 259565 372604
rect 259499 372539 259565 372540
rect 260051 372604 260117 372605
rect 260051 372540 260052 372604
rect 260116 372540 260117 372604
rect 260051 372539 260117 372540
rect 258395 371652 258461 371653
rect 258395 371588 258396 371652
rect 258460 371588 258461 371652
rect 258395 371587 258461 371588
rect 260974 371517 261034 374990
rect 261342 373149 261402 374990
rect 261339 373148 261405 373149
rect 261339 373084 261340 373148
rect 261404 373084 261405 373148
rect 261339 373083 261405 373084
rect 260971 371516 261037 371517
rect 260971 371452 260972 371516
rect 261036 371452 261037 371516
rect 260971 371451 261037 371452
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 350308 258134 366618
rect 261234 370894 261854 373000
rect 262262 372605 262322 374990
rect 262259 372604 262325 372605
rect 262259 372540 262260 372604
rect 262324 372540 262325 372604
rect 262259 372539 262325 372540
rect 263550 371517 263610 375050
rect 263731 374988 263732 375052
rect 263796 375050 263797 375052
rect 315251 375052 315317 375053
rect 263796 374990 263966 375050
rect 265022 374990 265326 375050
rect 265758 374990 266006 375050
rect 266310 374990 266414 375050
rect 267046 374990 267638 375050
rect 267782 374990 268318 375050
rect 268518 374990 268726 375050
rect 269254 374990 269814 375050
rect 270910 374990 271038 375050
rect 263796 374988 263797 374990
rect 263731 374987 263797 374988
rect 265022 373149 265082 374990
rect 265019 373148 265085 373149
rect 265019 373084 265020 373148
rect 265084 373084 265085 373148
rect 265019 373083 265085 373084
rect 263547 371516 263613 371517
rect 263547 371452 263548 371516
rect 263612 371452 263613 371516
rect 263547 371451 263613 371452
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 350308 261854 370338
rect 264954 357554 265574 373000
rect 265758 371517 265818 374990
rect 266310 374101 266370 374990
rect 266307 374100 266373 374101
rect 266307 374036 266308 374100
rect 266372 374036 266373 374100
rect 266307 374035 266373 374036
rect 267046 372605 267106 374990
rect 267043 372604 267109 372605
rect 267043 372540 267044 372604
rect 267108 372540 267109 372604
rect 267043 372539 267109 372540
rect 267782 371517 267842 374990
rect 268518 373829 268578 374990
rect 268515 373828 268581 373829
rect 268515 373764 268516 373828
rect 268580 373764 268581 373828
rect 268515 373763 268581 373764
rect 269254 373421 269314 374990
rect 269251 373420 269317 373421
rect 269251 373356 269252 373420
rect 269316 373356 269317 373420
rect 269251 373355 269317 373356
rect 265755 371516 265821 371517
rect 265755 371452 265756 371516
rect 265820 371452 265821 371516
rect 265755 371451 265821 371452
rect 267779 371516 267845 371517
rect 267779 371452 267780 371516
rect 267844 371452 267845 371516
rect 267779 371451 267845 371452
rect 270910 371381 270970 374990
rect 271144 374509 271204 375020
rect 272262 374990 272626 375050
rect 271141 374508 271207 374509
rect 271141 374444 271142 374508
rect 271206 374444 271207 374508
rect 271141 374443 271207 374444
rect 270907 371380 270973 371381
rect 270907 371316 270908 371380
rect 270972 371316 270973 371380
rect 270907 371315 270973 371316
rect 264954 357318 264986 357554
rect 265222 357318 265306 357554
rect 265542 357318 265574 357554
rect 264954 357234 265574 357318
rect 264954 356998 264986 357234
rect 265222 356998 265306 357234
rect 265542 356998 265574 357234
rect 264954 350308 265574 356998
rect 271794 362514 272414 373000
rect 272566 372605 272626 374990
rect 272563 372604 272629 372605
rect 272563 372540 272564 372604
rect 272628 372540 272629 372604
rect 272563 372539 272629 372540
rect 273302 372197 273362 375050
rect 273622 374990 273730 375050
rect 273299 372196 273365 372197
rect 273299 372132 273300 372196
rect 273364 372132 273365 372196
rect 273299 372131 273365 372132
rect 273670 371381 273730 374990
rect 273854 374990 274438 375050
rect 273854 372605 273914 374990
rect 275768 374509 275828 375020
rect 276070 374990 276306 375050
rect 275765 374508 275831 374509
rect 275765 374444 275766 374508
rect 275830 374444 275831 374508
rect 275765 374443 275831 374444
rect 273851 372604 273917 372605
rect 273851 372540 273852 372604
rect 273916 372540 273917 372604
rect 273851 372539 273917 372540
rect 273667 371380 273733 371381
rect 273667 371316 273668 371380
rect 273732 371316 273733 371380
rect 273667 371315 273733 371316
rect 271794 362278 271826 362514
rect 272062 362278 272146 362514
rect 272382 362278 272414 362514
rect 271794 362194 272414 362278
rect 271794 361958 271826 362194
rect 272062 361958 272146 362194
rect 272382 361958 272414 362194
rect 271794 350308 272414 361958
rect 275514 366234 276134 373000
rect 276246 371381 276306 374990
rect 276430 374990 277022 375050
rect 277534 374990 278110 375050
rect 278270 374990 278518 375050
rect 279006 374990 279198 375050
rect 280294 374990 280966 375050
rect 283550 374990 283850 375050
rect 276430 371789 276490 374990
rect 277534 372333 277594 374990
rect 277531 372332 277597 372333
rect 277531 372268 277532 372332
rect 277596 372268 277597 372332
rect 277531 372267 277597 372268
rect 276427 371788 276493 371789
rect 276427 371724 276428 371788
rect 276492 371724 276493 371788
rect 276427 371723 276493 371724
rect 277534 371517 277594 372267
rect 277531 371516 277597 371517
rect 277531 371452 277532 371516
rect 277596 371452 277597 371516
rect 277531 371451 277597 371452
rect 278270 371381 278330 374990
rect 279006 372469 279066 374990
rect 279003 372468 279069 372469
rect 279003 372404 279004 372468
rect 279068 372404 279069 372468
rect 279003 372403 279069 372404
rect 276243 371380 276309 371381
rect 276243 371316 276244 371380
rect 276308 371316 276309 371380
rect 276243 371315 276309 371316
rect 278267 371380 278333 371381
rect 278267 371316 278268 371380
rect 278332 371316 278333 371380
rect 278267 371315 278333 371316
rect 275514 365998 275546 366234
rect 275782 365998 275866 366234
rect 276102 365998 276134 366234
rect 275514 365914 276134 365998
rect 275514 365678 275546 365914
rect 275782 365678 275866 365914
rect 276102 365678 276134 365914
rect 275514 350308 276134 365678
rect 279234 352894 279854 373000
rect 280294 371381 280354 374990
rect 280291 371380 280357 371381
rect 280291 371316 280292 371380
rect 280356 371316 280357 371380
rect 280291 371315 280357 371316
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 350308 279854 352338
rect 282954 356614 283574 373000
rect 283790 371381 283850 374990
rect 285814 374990 285998 375050
rect 287654 374990 288310 375050
rect 290598 374990 291030 375050
rect 292806 374990 293478 375050
rect 295382 374990 295926 375050
rect 298142 374990 298510 375050
rect 285814 371381 285874 374990
rect 287654 371381 287714 374990
rect 283787 371380 283853 371381
rect 283787 371316 283788 371380
rect 283852 371316 283853 371380
rect 283787 371315 283853 371316
rect 285811 371380 285877 371381
rect 285811 371316 285812 371380
rect 285876 371316 285877 371380
rect 285811 371315 285877 371316
rect 287651 371380 287717 371381
rect 287651 371316 287652 371380
rect 287716 371316 287717 371380
rect 287651 371315 287717 371316
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 350308 283574 356058
rect 289794 363454 290414 373000
rect 290598 371381 290658 374990
rect 292806 372197 292866 374990
rect 292803 372196 292869 372197
rect 292803 372132 292804 372196
rect 292868 372132 292869 372196
rect 292803 372131 292869 372132
rect 290595 371380 290661 371381
rect 290595 371316 290596 371380
rect 290660 371316 290661 371380
rect 290595 371315 290661 371316
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 350308 290414 362898
rect 293514 367174 294134 373000
rect 295382 371381 295442 374990
rect 295379 371380 295445 371381
rect 295379 371316 295380 371380
rect 295444 371316 295445 371380
rect 295379 371315 295445 371316
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 350308 294134 366618
rect 297234 370894 297854 373000
rect 298142 371381 298202 374990
rect 300902 373149 300962 375050
rect 302926 374990 303542 375050
rect 305318 374990 305990 375050
rect 308574 374990 308690 375050
rect 300899 373148 300965 373149
rect 300899 373084 300900 373148
rect 300964 373084 300965 373148
rect 300899 373083 300965 373084
rect 298139 371380 298205 371381
rect 298139 371316 298140 371380
rect 298204 371316 298205 371380
rect 298139 371315 298205 371316
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 350308 297854 370338
rect 300954 357554 301574 373000
rect 302926 371789 302986 374990
rect 302923 371788 302989 371789
rect 302923 371724 302924 371788
rect 302988 371724 302989 371788
rect 302923 371723 302989 371724
rect 305318 371381 305378 374990
rect 305315 371380 305381 371381
rect 305315 371316 305316 371380
rect 305380 371316 305381 371380
rect 305315 371315 305381 371316
rect 300954 357318 300986 357554
rect 301222 357318 301306 357554
rect 301542 357318 301574 357554
rect 300954 357234 301574 357318
rect 300954 356998 300986 357234
rect 301222 356998 301306 357234
rect 301542 356998 301574 357234
rect 300954 350308 301574 356998
rect 307794 362514 308414 373000
rect 308630 371381 308690 374990
rect 310654 374990 311022 375050
rect 310654 371381 310714 374990
rect 308627 371380 308693 371381
rect 308627 371316 308628 371380
rect 308692 371316 308693 371380
rect 308627 371315 308693 371316
rect 310651 371380 310717 371381
rect 310651 371316 310652 371380
rect 310716 371316 310717 371380
rect 310651 371315 310717 371316
rect 307794 362278 307826 362514
rect 308062 362278 308146 362514
rect 308382 362278 308414 362514
rect 307794 362194 308414 362278
rect 307794 361958 307826 362194
rect 308062 361958 308146 362194
rect 308382 361958 308414 362194
rect 307794 350308 308414 361958
rect 311514 366234 312134 373000
rect 313414 371381 313474 375050
rect 315251 374988 315252 375052
rect 315316 375050 315317 375052
rect 315316 374990 315918 375050
rect 317830 374990 318502 375050
rect 315316 374988 315317 374990
rect 315251 374987 315317 374988
rect 317830 374781 317890 374990
rect 317827 374780 317893 374781
rect 317827 374716 317828 374780
rect 317892 374716 317893 374780
rect 317827 374715 317893 374716
rect 320920 374509 320980 375020
rect 322982 374990 323398 375050
rect 325982 374990 326722 375050
rect 320917 374508 320983 374509
rect 320917 374444 320918 374508
rect 320982 374444 320983 374508
rect 320917 374443 320983 374444
rect 313411 371380 313477 371381
rect 313411 371316 313412 371380
rect 313476 371316 313477 371380
rect 313411 371315 313477 371316
rect 311514 365998 311546 366234
rect 311782 365998 311866 366234
rect 312102 365998 312134 366234
rect 311514 365914 312134 365998
rect 311514 365678 311546 365914
rect 311782 365678 311866 365914
rect 312102 365678 312134 365914
rect 311514 350308 312134 365678
rect 315234 352894 315854 373000
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 350308 315854 352338
rect 318954 356614 319574 373000
rect 322982 371381 323042 374990
rect 322979 371380 323045 371381
rect 322979 371316 322980 371380
rect 323044 371316 323045 371380
rect 322979 371315 323045 371316
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 350308 319574 356058
rect 325794 363454 326414 373000
rect 326662 372605 326722 374990
rect 326659 372604 326725 372605
rect 326659 372540 326660 372604
rect 326724 372540 326725 372604
rect 326659 372539 326725 372540
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 350308 326414 362898
rect 329514 367174 330134 373000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 350308 330134 366618
rect 333234 370894 333854 373000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 350308 333854 370338
rect 336954 357554 337574 373000
rect 343222 372197 343282 375050
rect 343390 374990 343466 375050
rect 343406 372197 343466 374990
rect 343219 372196 343285 372197
rect 343219 372132 343220 372196
rect 343284 372132 343285 372196
rect 343219 372131 343285 372132
rect 343403 372196 343469 372197
rect 343403 372132 343404 372196
rect 343468 372132 343469 372196
rect 343403 372131 343469 372132
rect 336954 357318 336986 357554
rect 337222 357318 337306 357554
rect 337542 357318 337574 357554
rect 336954 357234 337574 357318
rect 336954 356998 336986 357234
rect 337222 356998 337306 357234
rect 337542 356998 337574 357234
rect 336954 350308 337574 356998
rect 343794 362514 344414 373000
rect 343794 362278 343826 362514
rect 344062 362278 344146 362514
rect 344382 362278 344414 362514
rect 343794 362194 344414 362278
rect 343794 361958 343826 362194
rect 344062 361958 344146 362194
rect 344382 361958 344414 362194
rect 338435 350572 338501 350573
rect 338435 350508 338436 350572
rect 338500 350508 338501 350572
rect 338435 350507 338501 350508
rect 339723 350572 339789 350573
rect 339723 350508 339724 350572
rect 339788 350508 339789 350572
rect 339723 350507 339789 350508
rect 338438 348530 338498 350507
rect 339726 348530 339786 350507
rect 343794 350308 344414 361958
rect 347514 366234 348134 373000
rect 347514 365998 347546 366234
rect 347782 365998 347866 366234
rect 348102 365998 348134 366234
rect 347514 365914 348134 365998
rect 347514 365678 347546 365914
rect 347782 365678 347866 365914
rect 348102 365678 348134 365914
rect 347514 350308 348134 365678
rect 351234 352894 351854 373000
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 350947 350572 351013 350573
rect 350947 350508 350948 350572
rect 351012 350508 351013 350572
rect 350947 350507 351013 350508
rect 350950 348530 351010 350507
rect 351234 350308 351854 352338
rect 354954 356614 355574 373000
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 350308 355574 356058
rect 338438 348470 338524 348530
rect 338464 348202 338524 348470
rect 339688 348470 339786 348530
rect 350840 348470 351010 348530
rect 339688 348202 339748 348470
rect 350840 348202 350900 348470
rect 220272 345454 220620 345486
rect 220272 345218 220328 345454
rect 220564 345218 220620 345454
rect 220272 345134 220620 345218
rect 220272 344898 220328 345134
rect 220564 344898 220620 345134
rect 220272 344866 220620 344898
rect 356000 345454 356348 345486
rect 356000 345218 356056 345454
rect 356292 345218 356348 345454
rect 356000 345134 356348 345218
rect 356000 344898 356056 345134
rect 356292 344898 356348 345134
rect 356000 344866 356348 344898
rect 220952 327454 221300 327486
rect 220952 327218 221008 327454
rect 221244 327218 221300 327454
rect 220952 327134 221300 327218
rect 220952 326898 221008 327134
rect 221244 326898 221300 327134
rect 220952 326866 221300 326898
rect 355320 327454 355668 327486
rect 355320 327218 355376 327454
rect 355612 327218 355668 327454
rect 355320 327134 355668 327218
rect 355320 326898 355376 327134
rect 355612 326898 355668 327134
rect 355320 326866 355668 326898
rect 220272 309454 220620 309486
rect 220272 309218 220328 309454
rect 220564 309218 220620 309454
rect 220272 309134 220620 309218
rect 220272 308898 220328 309134
rect 220564 308898 220620 309134
rect 220272 308866 220620 308898
rect 356000 309454 356348 309486
rect 356000 309218 356056 309454
rect 356292 309218 356348 309454
rect 356000 309134 356348 309218
rect 356000 308898 356056 309134
rect 356292 308898 356348 309134
rect 356000 308866 356348 308898
rect 220952 291454 221300 291486
rect 220952 291218 221008 291454
rect 221244 291218 221300 291454
rect 220952 291134 221300 291218
rect 220952 290898 221008 291134
rect 221244 290898 221300 291134
rect 220952 290866 221300 290898
rect 355320 291454 355668 291486
rect 355320 291218 355376 291454
rect 355612 291218 355668 291454
rect 355320 291134 355668 291218
rect 355320 290898 355376 291134
rect 355612 290898 355668 291134
rect 355320 290866 355668 290898
rect 220272 273454 220620 273486
rect 220272 273218 220328 273454
rect 220564 273218 220620 273454
rect 220272 273134 220620 273218
rect 220272 272898 220328 273134
rect 220564 272898 220620 273134
rect 220272 272866 220620 272898
rect 356000 273454 356348 273486
rect 356000 273218 356056 273454
rect 356292 273218 356348 273454
rect 356000 273134 356348 273218
rect 356000 272898 356056 273134
rect 356292 272898 356348 273134
rect 356000 272866 356348 272898
rect 236056 264890 236116 265106
rect 237144 264890 237204 265106
rect 238232 264890 238292 265106
rect 235950 264830 236116 264890
rect 237054 264830 237204 264890
rect 238158 264830 238292 264890
rect 239592 264890 239652 265106
rect 240544 264890 240604 265106
rect 241768 264890 241828 265106
rect 243128 264890 243188 265106
rect 239592 264830 239690 264890
rect 240544 264830 240610 264890
rect 235950 263533 236010 264830
rect 235947 263532 236013 263533
rect 235947 263468 235948 263532
rect 236012 263468 236013 263532
rect 235947 263467 236013 263468
rect 221514 259174 222134 263000
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 240308 222134 258618
rect 225234 262894 225854 263000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 240308 225854 262338
rect 228954 249554 229574 263000
rect 228954 249318 228986 249554
rect 229222 249318 229306 249554
rect 229542 249318 229574 249554
rect 228954 249234 229574 249318
rect 228954 248998 228986 249234
rect 229222 248998 229306 249234
rect 229542 248998 229574 249234
rect 228954 240308 229574 248998
rect 235794 254514 236414 263000
rect 237054 262989 237114 264830
rect 237051 262988 237117 262989
rect 237051 262924 237052 262988
rect 237116 262924 237117 262988
rect 237051 262923 237117 262924
rect 238158 262309 238218 264830
rect 239630 263533 239690 264830
rect 239627 263532 239693 263533
rect 239627 263468 239628 263532
rect 239692 263468 239693 263532
rect 239627 263467 239693 263468
rect 238155 262308 238221 262309
rect 238155 262244 238156 262308
rect 238220 262244 238221 262308
rect 238155 262243 238221 262244
rect 235794 254278 235826 254514
rect 236062 254278 236146 254514
rect 236382 254278 236414 254514
rect 235794 254194 236414 254278
rect 235794 253958 235826 254194
rect 236062 253958 236146 254194
rect 236382 253958 236414 254194
rect 235794 240308 236414 253958
rect 239514 241174 240134 263000
rect 240550 262309 240610 264830
rect 241654 264830 241828 264890
rect 243126 264830 243188 264890
rect 244216 264890 244276 265106
rect 245440 264890 245500 265106
rect 246528 264890 246588 265106
rect 247616 264890 247676 265106
rect 248296 264890 248356 265106
rect 248704 264890 248764 265106
rect 244216 264830 244290 264890
rect 241654 262309 241714 264830
rect 243126 263533 243186 264830
rect 243123 263532 243189 263533
rect 243123 263468 243124 263532
rect 243188 263468 243189 263532
rect 243123 263467 243189 263468
rect 240547 262308 240613 262309
rect 240547 262244 240548 262308
rect 240612 262244 240613 262308
rect 240547 262243 240613 262244
rect 241651 262308 241717 262309
rect 241651 262244 241652 262308
rect 241716 262244 241717 262308
rect 241651 262243 241717 262244
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 240308 240134 240618
rect 243234 244894 243854 263000
rect 244230 262989 244290 264830
rect 245334 264830 245500 264890
rect 246438 264830 246588 264890
rect 247542 264830 247676 264890
rect 248278 264830 248356 264890
rect 248646 264830 248764 264890
rect 250064 264890 250124 265106
rect 250483 265028 250549 265029
rect 250483 264964 250484 265028
rect 250548 264964 250549 265028
rect 250483 264963 250549 264964
rect 250486 264890 250546 264963
rect 250744 264890 250804 265106
rect 251288 264890 251348 265106
rect 252376 264890 252436 265106
rect 253464 264890 253524 265106
rect 250064 264830 250178 264890
rect 250486 264830 250804 264890
rect 251222 264830 251348 264890
rect 252326 264830 252436 264890
rect 253430 264830 253524 264890
rect 253600 264890 253660 265106
rect 254552 264890 254612 265106
rect 255912 264890 255972 265106
rect 253600 264830 253674 264890
rect 244227 262988 244293 262989
rect 244227 262924 244228 262988
rect 244292 262924 244293 262988
rect 244227 262923 244293 262924
rect 245334 262309 245394 264830
rect 246438 262309 246498 264830
rect 247542 263533 247602 264830
rect 248278 263533 248338 264830
rect 247539 263532 247605 263533
rect 247539 263468 247540 263532
rect 247604 263468 247605 263532
rect 247539 263467 247605 263468
rect 248275 263532 248341 263533
rect 248275 263468 248276 263532
rect 248340 263468 248341 263532
rect 248275 263467 248341 263468
rect 245331 262308 245397 262309
rect 245331 262244 245332 262308
rect 245396 262244 245397 262308
rect 245331 262243 245397 262244
rect 246435 262308 246501 262309
rect 246435 262244 246436 262308
rect 246500 262244 246501 262308
rect 246435 262243 246501 262244
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 240308 243854 244338
rect 246954 248614 247574 263000
rect 248646 262309 248706 264830
rect 250118 262309 250178 264830
rect 251222 262309 251282 264830
rect 252326 262445 252386 264830
rect 252323 262444 252389 262445
rect 252323 262380 252324 262444
rect 252388 262380 252389 262444
rect 252323 262379 252389 262380
rect 253430 262309 253490 264830
rect 253614 263533 253674 264830
rect 254534 264830 254612 264890
rect 255822 264830 255972 264890
rect 256048 264890 256108 265106
rect 257000 264890 257060 265106
rect 256048 264830 256250 264890
rect 253611 263532 253677 263533
rect 253611 263468 253612 263532
rect 253676 263468 253677 263532
rect 253611 263467 253677 263468
rect 248643 262308 248709 262309
rect 248643 262244 248644 262308
rect 248708 262244 248709 262308
rect 248643 262243 248709 262244
rect 250115 262308 250181 262309
rect 250115 262244 250116 262308
rect 250180 262244 250181 262308
rect 250115 262243 250181 262244
rect 251219 262308 251285 262309
rect 251219 262244 251220 262308
rect 251284 262244 251285 262308
rect 251219 262243 251285 262244
rect 253427 262308 253493 262309
rect 253427 262244 253428 262308
rect 253492 262244 253493 262308
rect 253427 262243 253493 262244
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 240308 247574 248058
rect 253794 255454 254414 263000
rect 254534 262309 254594 264830
rect 255822 262309 255882 264830
rect 256190 263533 256250 264830
rect 256926 264830 257060 264890
rect 258088 264890 258148 265106
rect 258496 264890 258556 265106
rect 258088 264830 258274 264890
rect 256187 263532 256253 263533
rect 256187 263468 256188 263532
rect 256252 263468 256253 263532
rect 256187 263467 256253 263468
rect 256926 262309 256986 264830
rect 258214 263533 258274 264830
rect 258398 264830 258556 264890
rect 259448 264890 259508 265106
rect 260672 264890 260732 265106
rect 261080 264890 261140 265106
rect 261760 264890 261820 265106
rect 262848 264890 262908 265106
rect 259448 264830 259562 264890
rect 258211 263532 258277 263533
rect 258211 263468 258212 263532
rect 258276 263468 258277 263532
rect 258211 263467 258277 263468
rect 254531 262308 254597 262309
rect 254531 262244 254532 262308
rect 254596 262244 254597 262308
rect 254531 262243 254597 262244
rect 255819 262308 255885 262309
rect 255819 262244 255820 262308
rect 255884 262244 255885 262308
rect 255819 262243 255885 262244
rect 256923 262308 256989 262309
rect 256923 262244 256924 262308
rect 256988 262244 256989 262308
rect 256923 262243 256989 262244
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 240308 254414 254898
rect 257514 259174 258134 263000
rect 258398 262989 258458 264830
rect 258395 262988 258461 262989
rect 258395 262924 258396 262988
rect 258460 262924 258461 262988
rect 258395 262923 258461 262924
rect 259502 262309 259562 264830
rect 260606 264830 260732 264890
rect 260974 264830 261140 264890
rect 261710 264830 261820 264890
rect 262814 264830 262908 264890
rect 263528 264890 263588 265106
rect 263936 264890 263996 265106
rect 265296 264890 265356 265106
rect 265976 264890 266036 265106
rect 266384 264890 266444 265106
rect 267608 264890 267668 265106
rect 263528 264830 263610 264890
rect 260606 262445 260666 264830
rect 260974 262989 261034 264830
rect 261710 263533 261770 264830
rect 262814 263533 262874 264830
rect 263550 263533 263610 264830
rect 263918 264830 263996 264890
rect 265206 264830 265356 264890
rect 265942 264830 266036 264890
rect 266310 264830 266444 264890
rect 267598 264830 267668 264890
rect 268288 264890 268348 265106
rect 268696 264890 268756 265106
rect 269784 264890 269844 265106
rect 271008 264890 271068 265106
rect 268288 264830 268394 264890
rect 268696 264830 268762 264890
rect 269784 264830 269866 264890
rect 261707 263532 261773 263533
rect 261707 263468 261708 263532
rect 261772 263468 261773 263532
rect 261707 263467 261773 263468
rect 262811 263532 262877 263533
rect 262811 263468 262812 263532
rect 262876 263468 262877 263532
rect 262811 263467 262877 263468
rect 263547 263532 263613 263533
rect 263547 263468 263548 263532
rect 263612 263468 263613 263532
rect 263547 263467 263613 263468
rect 260971 262988 261037 262989
rect 260971 262924 260972 262988
rect 261036 262924 261037 262988
rect 260971 262923 261037 262924
rect 261234 262894 261854 263000
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 260603 262444 260669 262445
rect 260603 262380 260604 262444
rect 260668 262380 260669 262444
rect 260603 262379 260669 262380
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 259499 262308 259565 262309
rect 259499 262244 259500 262308
rect 259564 262244 259565 262308
rect 259499 262243 259565 262244
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 240308 258134 258618
rect 261234 240308 261854 262338
rect 263918 262309 263978 264830
rect 265206 263533 265266 264830
rect 265942 263533 266002 264830
rect 265203 263532 265269 263533
rect 265203 263468 265204 263532
rect 265268 263468 265269 263532
rect 265203 263467 265269 263468
rect 265939 263532 266005 263533
rect 265939 263468 265940 263532
rect 266004 263468 266005 263532
rect 265939 263467 266005 263468
rect 263915 262308 263981 262309
rect 263915 262244 263916 262308
rect 263980 262244 263981 262308
rect 263915 262243 263981 262244
rect 264954 249554 265574 263000
rect 266310 262309 266370 264830
rect 267598 262445 267658 264830
rect 268334 263533 268394 264830
rect 268331 263532 268397 263533
rect 268331 263468 268332 263532
rect 268396 263468 268397 263532
rect 268331 263467 268397 263468
rect 267595 262444 267661 262445
rect 267595 262380 267596 262444
rect 267660 262380 267661 262444
rect 267595 262379 267661 262380
rect 268702 262309 268762 264830
rect 269806 263533 269866 264830
rect 270910 264830 271068 264890
rect 271144 264890 271204 265106
rect 272232 264890 272292 265106
rect 273320 264890 273380 265106
rect 273592 264890 273652 265106
rect 274219 265028 274285 265029
rect 274219 264964 274220 265028
rect 274284 264964 274285 265028
rect 274219 264963 274285 264964
rect 271144 264830 271338 264890
rect 270910 263533 270970 264830
rect 271278 263533 271338 264830
rect 272198 264830 272292 264890
rect 273302 264830 273380 264890
rect 273486 264830 273652 264890
rect 274222 264890 274282 264963
rect 274408 264890 274468 265106
rect 274222 264830 274468 264890
rect 275768 264890 275828 265106
rect 276040 264890 276100 265106
rect 276992 264890 277052 265106
rect 275768 264830 275938 264890
rect 276040 264830 276122 264890
rect 272198 263533 272258 264830
rect 273302 263533 273362 264830
rect 269803 263532 269869 263533
rect 269803 263468 269804 263532
rect 269868 263468 269869 263532
rect 269803 263467 269869 263468
rect 270907 263532 270973 263533
rect 270907 263468 270908 263532
rect 270972 263468 270973 263532
rect 270907 263467 270973 263468
rect 271275 263532 271341 263533
rect 271275 263468 271276 263532
rect 271340 263468 271341 263532
rect 271275 263467 271341 263468
rect 272195 263532 272261 263533
rect 272195 263468 272196 263532
rect 272260 263468 272261 263532
rect 272195 263467 272261 263468
rect 273299 263532 273365 263533
rect 273299 263468 273300 263532
rect 273364 263468 273365 263532
rect 273299 263467 273365 263468
rect 266307 262308 266373 262309
rect 266307 262244 266308 262308
rect 266372 262244 266373 262308
rect 266307 262243 266373 262244
rect 268699 262308 268765 262309
rect 268699 262244 268700 262308
rect 268764 262244 268765 262308
rect 268699 262243 268765 262244
rect 264954 249318 264986 249554
rect 265222 249318 265306 249554
rect 265542 249318 265574 249554
rect 264954 249234 265574 249318
rect 264954 248998 264986 249234
rect 265222 248998 265306 249234
rect 265542 248998 265574 249234
rect 264954 240308 265574 248998
rect 271794 254514 272414 263000
rect 273486 262989 273546 264830
rect 275878 263533 275938 264830
rect 276062 263533 276122 264830
rect 276982 264830 277052 264890
rect 278080 264890 278140 265106
rect 278488 264890 278548 265106
rect 278080 264830 278146 264890
rect 275875 263532 275941 263533
rect 275875 263468 275876 263532
rect 275940 263468 275941 263532
rect 275875 263467 275941 263468
rect 276059 263532 276125 263533
rect 276059 263468 276060 263532
rect 276124 263468 276125 263532
rect 276059 263467 276125 263468
rect 273483 262988 273549 262989
rect 273483 262924 273484 262988
rect 273548 262924 273549 262988
rect 273483 262923 273549 262924
rect 271794 254278 271826 254514
rect 272062 254278 272146 254514
rect 272382 254278 272414 254514
rect 271794 254194 272414 254278
rect 271794 253958 271826 254194
rect 272062 253958 272146 254194
rect 272382 253958 272414 254194
rect 271794 240308 272414 253958
rect 275514 241174 276134 263000
rect 276982 262309 277042 264830
rect 278086 262309 278146 264830
rect 278454 264830 278548 264890
rect 279168 264890 279228 265106
rect 280936 264890 280996 265106
rect 283520 264890 283580 265106
rect 279168 264830 279250 264890
rect 278454 263125 278514 264830
rect 279190 263533 279250 264830
rect 280846 264830 280996 264890
rect 283422 264830 283580 264890
rect 285968 264890 286028 265106
rect 288280 264890 288340 265106
rect 291000 264890 291060 265106
rect 285968 264830 286058 264890
rect 280846 264349 280906 264830
rect 283422 264349 283482 264830
rect 285998 264349 286058 264830
rect 288206 264830 288340 264890
rect 290966 264830 291060 264890
rect 288206 264349 288266 264830
rect 290966 264349 291026 264830
rect 293448 264621 293508 265106
rect 295896 264890 295956 265106
rect 298480 264890 298540 265106
rect 300928 264890 300988 265106
rect 303512 264890 303572 265106
rect 305960 264890 306020 265106
rect 308544 264890 308604 265106
rect 295896 264830 295994 264890
rect 298480 264830 298570 264890
rect 293445 264620 293511 264621
rect 293445 264556 293446 264620
rect 293510 264556 293511 264620
rect 293445 264555 293511 264556
rect 280843 264348 280909 264349
rect 280843 264284 280844 264348
rect 280908 264284 280909 264348
rect 280843 264283 280909 264284
rect 283419 264348 283485 264349
rect 283419 264284 283420 264348
rect 283484 264284 283485 264348
rect 283419 264283 283485 264284
rect 285995 264348 286061 264349
rect 285995 264284 285996 264348
rect 286060 264284 286061 264348
rect 285995 264283 286061 264284
rect 288203 264348 288269 264349
rect 288203 264284 288204 264348
rect 288268 264284 288269 264348
rect 288203 264283 288269 264284
rect 290963 264348 291029 264349
rect 290963 264284 290964 264348
rect 291028 264284 291029 264348
rect 290963 264283 291029 264284
rect 295934 264213 295994 264830
rect 298510 264349 298570 264830
rect 300902 264830 300988 264890
rect 303478 264830 303572 264890
rect 305870 264830 306020 264890
rect 308446 264830 308604 264890
rect 300902 264485 300962 264830
rect 300899 264484 300965 264485
rect 300899 264420 300900 264484
rect 300964 264420 300965 264484
rect 300899 264419 300965 264420
rect 298507 264348 298573 264349
rect 298507 264284 298508 264348
rect 298572 264284 298573 264348
rect 298507 264283 298573 264284
rect 295931 264212 295997 264213
rect 295931 264148 295932 264212
rect 295996 264148 295997 264212
rect 295931 264147 295997 264148
rect 279187 263532 279253 263533
rect 279187 263468 279188 263532
rect 279252 263468 279253 263532
rect 279187 263467 279253 263468
rect 278451 263124 278517 263125
rect 278451 263060 278452 263124
rect 278516 263060 278517 263124
rect 278451 263059 278517 263060
rect 276979 262308 277045 262309
rect 276979 262244 276980 262308
rect 277044 262244 277045 262308
rect 276979 262243 277045 262244
rect 278083 262308 278149 262309
rect 278083 262244 278084 262308
rect 278148 262244 278149 262308
rect 278083 262243 278149 262244
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 240308 276134 240618
rect 279234 244894 279854 263000
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 240308 279854 244338
rect 282954 248614 283574 263000
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 240308 283574 248058
rect 289794 255454 290414 263000
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 240308 290414 254898
rect 293514 259174 294134 263000
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 240308 294134 258618
rect 297234 262894 297854 263000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 240308 297854 262338
rect 300954 249554 301574 263000
rect 303478 262309 303538 264830
rect 305870 263533 305930 264830
rect 308446 263533 308506 264830
rect 310992 264757 311052 265106
rect 313440 264890 313500 265106
rect 315888 264890 315948 265106
rect 318472 264893 318532 265106
rect 313414 264830 313500 264890
rect 315806 264830 315948 264890
rect 318469 264892 318535 264893
rect 310989 264756 311055 264757
rect 310989 264692 310990 264756
rect 311054 264692 311055 264756
rect 310989 264691 311055 264692
rect 305867 263532 305933 263533
rect 305867 263468 305868 263532
rect 305932 263468 305933 263532
rect 305867 263467 305933 263468
rect 308443 263532 308509 263533
rect 308443 263468 308444 263532
rect 308508 263468 308509 263532
rect 308443 263467 308509 263468
rect 313414 263261 313474 264830
rect 315806 263261 315866 264830
rect 318469 264828 318470 264892
rect 318534 264828 318535 264892
rect 320920 264890 320980 265106
rect 323368 264890 323428 265106
rect 325952 264890 326012 265106
rect 343224 264890 343284 265106
rect 320920 264830 321018 264890
rect 318469 264827 318535 264828
rect 320958 263397 321018 264830
rect 323350 264830 323428 264890
rect 325926 264830 326012 264890
rect 343222 264830 343284 264890
rect 343360 264890 343420 265106
rect 343360 264830 343466 264890
rect 323350 263533 323410 264830
rect 325926 263533 325986 264830
rect 343222 263533 343282 264830
rect 323347 263532 323413 263533
rect 323347 263468 323348 263532
rect 323412 263468 323413 263532
rect 323347 263467 323413 263468
rect 325923 263532 325989 263533
rect 325923 263468 325924 263532
rect 325988 263468 325989 263532
rect 325923 263467 325989 263468
rect 343219 263532 343285 263533
rect 343219 263468 343220 263532
rect 343284 263468 343285 263532
rect 343219 263467 343285 263468
rect 320955 263396 321021 263397
rect 320955 263332 320956 263396
rect 321020 263332 321021 263396
rect 320955 263331 321021 263332
rect 313411 263260 313477 263261
rect 313411 263196 313412 263260
rect 313476 263196 313477 263260
rect 313411 263195 313477 263196
rect 315803 263260 315869 263261
rect 315803 263196 315804 263260
rect 315868 263196 315869 263260
rect 315803 263195 315869 263196
rect 343406 263125 343466 264830
rect 343403 263124 343469 263125
rect 343403 263060 343404 263124
rect 343468 263060 343469 263124
rect 343403 263059 343469 263060
rect 303475 262308 303541 262309
rect 303475 262244 303476 262308
rect 303540 262244 303541 262308
rect 303475 262243 303541 262244
rect 300954 249318 300986 249554
rect 301222 249318 301306 249554
rect 301542 249318 301574 249554
rect 300954 249234 301574 249318
rect 300954 248998 300986 249234
rect 301222 248998 301306 249234
rect 301542 248998 301574 249234
rect 300954 240308 301574 248998
rect 307794 254514 308414 263000
rect 307794 254278 307826 254514
rect 308062 254278 308146 254514
rect 308382 254278 308414 254514
rect 307794 254194 308414 254278
rect 307794 253958 307826 254194
rect 308062 253958 308146 254194
rect 308382 253958 308414 254194
rect 307794 240308 308414 253958
rect 311514 241174 312134 263000
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 240308 312134 240618
rect 315234 244894 315854 263000
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 240308 315854 244338
rect 318954 248614 319574 263000
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 240308 319574 248058
rect 325794 255454 326414 263000
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 240308 326414 254898
rect 329514 259174 330134 263000
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 240308 330134 258618
rect 333234 262894 333854 263000
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 240308 333854 262338
rect 336954 249554 337574 263000
rect 336954 249318 336986 249554
rect 337222 249318 337306 249554
rect 337542 249318 337574 249554
rect 336954 249234 337574 249318
rect 336954 248998 336986 249234
rect 337222 248998 337306 249234
rect 337542 248998 337574 249234
rect 336954 240308 337574 248998
rect 343794 254514 344414 263000
rect 343794 254278 343826 254514
rect 344062 254278 344146 254514
rect 344382 254278 344414 254514
rect 343794 254194 344414 254278
rect 343794 253958 343826 254194
rect 344062 253958 344146 254194
rect 344382 253958 344414 254194
rect 343794 240308 344414 253958
rect 347514 241174 348134 263000
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 240308 348134 240618
rect 351234 244894 351854 263000
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 240308 351854 244338
rect 354954 248614 355574 263000
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 240308 355574 248058
rect 338435 240276 338501 240277
rect 338435 240212 338436 240276
rect 338500 240212 338501 240276
rect 338435 240211 338501 240212
rect 339723 240276 339789 240277
rect 339723 240212 339724 240276
rect 339788 240212 339789 240276
rect 339723 240211 339789 240212
rect 350947 240276 351013 240277
rect 350947 240212 350948 240276
rect 351012 240212 351013 240276
rect 350947 240211 351013 240212
rect 338438 238770 338498 240211
rect 339726 238770 339786 240211
rect 350950 238770 351010 240211
rect 338438 238710 338524 238770
rect 338464 238202 338524 238710
rect 339688 238710 339786 238770
rect 350840 238710 351010 238770
rect 339688 238202 339748 238710
rect 350840 238202 350900 238710
rect 220272 237454 220620 237486
rect 220272 237218 220328 237454
rect 220564 237218 220620 237454
rect 220272 237134 220620 237218
rect 220272 236898 220328 237134
rect 220564 236898 220620 237134
rect 220272 236866 220620 236898
rect 356000 237454 356348 237486
rect 356000 237218 356056 237454
rect 356292 237218 356348 237454
rect 356000 237134 356348 237218
rect 356000 236898 356056 237134
rect 356292 236898 356348 237134
rect 356000 236866 356348 236898
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 201454 220620 201486
rect 220272 201218 220328 201454
rect 220564 201218 220620 201454
rect 220272 201134 220620 201218
rect 220272 200898 220328 201134
rect 220564 200898 220620 201134
rect 220272 200866 220620 200898
rect 356000 201454 356348 201486
rect 356000 201218 356056 201454
rect 356292 201218 356348 201454
rect 356000 201134 356348 201218
rect 356000 200898 356056 201134
rect 356292 200898 356348 201134
rect 356000 200866 356348 200898
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 220272 165454 220620 165486
rect 220272 165218 220328 165454
rect 220564 165218 220620 165454
rect 220272 165134 220620 165218
rect 220272 164898 220328 165134
rect 220564 164898 220620 165134
rect 220272 164866 220620 164898
rect 356000 165454 356348 165486
rect 356000 165218 356056 165454
rect 356292 165218 356348 165454
rect 356000 165134 356348 165218
rect 356000 164898 356056 165134
rect 356292 164898 356348 165134
rect 356000 164866 356348 164898
rect 236056 154590 236116 155040
rect 237144 154590 237204 155040
rect 238232 154590 238292 155040
rect 239592 154730 239652 155040
rect 238894 154670 239652 154730
rect 238894 154590 238954 154670
rect 236056 154530 236194 154590
rect 236134 153237 236194 154530
rect 237054 154530 237204 154590
rect 238158 154530 238292 154590
rect 238526 154530 238954 154590
rect 240544 154590 240604 155040
rect 241768 154590 241828 155040
rect 243128 154590 243188 155040
rect 244216 154730 244276 155040
rect 244216 154670 244290 154730
rect 240544 154530 240610 154590
rect 236131 153236 236197 153237
rect 236131 153172 236132 153236
rect 236196 153172 236197 153236
rect 236131 153171 236197 153172
rect 221514 151174 222134 153000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 130308 222134 150618
rect 225234 137834 225854 153000
rect 225234 137598 225266 137834
rect 225502 137598 225586 137834
rect 225822 137598 225854 137834
rect 225234 137514 225854 137598
rect 225234 137278 225266 137514
rect 225502 137278 225586 137514
rect 225822 137278 225854 137514
rect 225234 130308 225854 137278
rect 228954 141554 229574 153000
rect 228954 141318 228986 141554
rect 229222 141318 229306 141554
rect 229542 141318 229574 141554
rect 228954 141234 229574 141318
rect 228954 140998 228986 141234
rect 229222 140998 229306 141234
rect 229542 140998 229574 141234
rect 228954 130308 229574 140998
rect 235794 146514 236414 153000
rect 237054 152421 237114 154530
rect 238158 153101 238218 154530
rect 238155 153100 238221 153101
rect 238155 153036 238156 153100
rect 238220 153036 238221 153100
rect 238155 153035 238221 153036
rect 237051 152420 237117 152421
rect 237051 152356 237052 152420
rect 237116 152356 237117 152420
rect 237051 152355 237117 152356
rect 238526 152010 238586 154530
rect 240550 153101 240610 154530
rect 241654 154530 241828 154590
rect 242942 154530 243188 154590
rect 241654 153101 241714 154530
rect 242942 153101 243002 154530
rect 244230 153101 244290 154670
rect 245440 154590 245500 155040
rect 246528 154590 246588 155040
rect 245334 154530 245500 154590
rect 246438 154530 246588 154590
rect 247616 154590 247676 155040
rect 248296 154590 248356 155040
rect 248704 154590 248764 155040
rect 247616 154530 247786 154590
rect 240547 153100 240613 153101
rect 240547 153036 240548 153100
rect 240612 153036 240613 153100
rect 240547 153035 240613 153036
rect 241651 153100 241717 153101
rect 241651 153036 241652 153100
rect 241716 153036 241717 153100
rect 241651 153035 241717 153036
rect 242939 153100 243005 153101
rect 242939 153036 242940 153100
rect 243004 153036 243005 153100
rect 242939 153035 243005 153036
rect 244227 153100 244293 153101
rect 244227 153036 244228 153100
rect 244292 153036 244293 153100
rect 244227 153035 244293 153036
rect 238707 152012 238773 152013
rect 238707 152010 238708 152012
rect 238526 151950 238708 152010
rect 238707 151948 238708 151950
rect 238772 151948 238773 152012
rect 238707 151947 238773 151948
rect 235794 146278 235826 146514
rect 236062 146278 236146 146514
rect 236382 146278 236414 146514
rect 235794 146194 236414 146278
rect 235794 145958 235826 146194
rect 236062 145958 236146 146194
rect 236382 145958 236414 146194
rect 235794 130308 236414 145958
rect 239514 133174 240134 153000
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 130308 240134 132618
rect 243234 136894 243854 153000
rect 245334 152421 245394 154530
rect 246438 153101 246498 154530
rect 247726 153101 247786 154530
rect 248278 154530 248356 154590
rect 248646 154530 248764 154590
rect 250064 154590 250124 155040
rect 250744 154590 250804 155040
rect 251288 154590 251348 155040
rect 252376 154590 252436 155040
rect 253464 154590 253524 155040
rect 250064 154530 250178 154590
rect 246435 153100 246501 153101
rect 246435 153036 246436 153100
rect 246500 153036 246501 153100
rect 246435 153035 246501 153036
rect 247723 153100 247789 153101
rect 247723 153036 247724 153100
rect 247788 153036 247789 153100
rect 247723 153035 247789 153036
rect 245331 152420 245397 152421
rect 245331 152356 245332 152420
rect 245396 152356 245397 152420
rect 245331 152355 245397 152356
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 130308 243854 136338
rect 246954 140614 247574 153000
rect 248278 152421 248338 154530
rect 248646 153101 248706 154530
rect 250118 153101 250178 154530
rect 250670 154530 250804 154590
rect 251222 154530 251348 154590
rect 252326 154530 252436 154590
rect 253430 154530 253524 154590
rect 253600 154590 253660 155040
rect 254552 154590 254612 155040
rect 255912 154590 255972 155040
rect 253600 154530 253674 154590
rect 250670 153101 250730 154530
rect 251222 153101 251282 154530
rect 248643 153100 248709 153101
rect 248643 153036 248644 153100
rect 248708 153036 248709 153100
rect 248643 153035 248709 153036
rect 250115 153100 250181 153101
rect 250115 153036 250116 153100
rect 250180 153036 250181 153100
rect 250115 153035 250181 153036
rect 250667 153100 250733 153101
rect 250667 153036 250668 153100
rect 250732 153036 250733 153100
rect 250667 153035 250733 153036
rect 251219 153100 251285 153101
rect 251219 153036 251220 153100
rect 251284 153036 251285 153100
rect 251219 153035 251285 153036
rect 252326 152421 252386 154530
rect 253430 153101 253490 154530
rect 253614 153101 253674 154530
rect 254534 154530 254612 154590
rect 255822 154530 255972 154590
rect 256048 154590 256108 155040
rect 257000 154590 257060 155040
rect 258088 154730 258148 155040
rect 258496 154730 258556 155040
rect 258088 154670 258274 154730
rect 256048 154530 256250 154590
rect 254534 153101 254594 154530
rect 255822 153101 255882 154530
rect 256190 153101 256250 154530
rect 256926 154530 257060 154590
rect 256926 153101 256986 154530
rect 258214 153101 258274 154670
rect 258398 154670 258556 154730
rect 259448 154730 259508 155040
rect 260672 154730 260732 155040
rect 259448 154670 259562 154730
rect 253427 153100 253493 153101
rect 253427 153036 253428 153100
rect 253492 153036 253493 153100
rect 253427 153035 253493 153036
rect 253611 153100 253677 153101
rect 253611 153036 253612 153100
rect 253676 153036 253677 153100
rect 253611 153035 253677 153036
rect 254531 153100 254597 153101
rect 254531 153036 254532 153100
rect 254596 153036 254597 153100
rect 254531 153035 254597 153036
rect 255819 153100 255885 153101
rect 255819 153036 255820 153100
rect 255884 153036 255885 153100
rect 255819 153035 255885 153036
rect 256187 153100 256253 153101
rect 256187 153036 256188 153100
rect 256252 153036 256253 153100
rect 256187 153035 256253 153036
rect 256923 153100 256989 153101
rect 256923 153036 256924 153100
rect 256988 153036 256989 153100
rect 256923 153035 256989 153036
rect 258211 153100 258277 153101
rect 258211 153036 258212 153100
rect 258276 153036 258277 153100
rect 258211 153035 258277 153036
rect 248275 152420 248341 152421
rect 248275 152356 248276 152420
rect 248340 152356 248341 152420
rect 248275 152355 248341 152356
rect 252323 152420 252389 152421
rect 252323 152356 252324 152420
rect 252388 152356 252389 152420
rect 252323 152355 252389 152356
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 130308 247574 140058
rect 253794 147454 254414 153000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 130308 254414 146898
rect 257514 151174 258134 153000
rect 258398 152557 258458 154670
rect 259502 153101 259562 154670
rect 260606 154670 260732 154730
rect 259499 153100 259565 153101
rect 259499 153036 259500 153100
rect 259564 153036 259565 153100
rect 259499 153035 259565 153036
rect 260606 152693 260666 154670
rect 261080 154597 261140 155040
rect 261760 154730 261820 155040
rect 262848 154730 262908 155040
rect 261710 154670 261820 154730
rect 262814 154670 262908 154730
rect 263528 154730 263588 155040
rect 263936 154730 263996 155040
rect 265296 154730 265356 155040
rect 265976 154730 266036 155040
rect 266384 154730 266444 155040
rect 267608 154730 267668 155040
rect 263528 154670 263610 154730
rect 261077 154596 261143 154597
rect 261077 154532 261078 154596
rect 261142 154532 261143 154596
rect 261077 154531 261143 154532
rect 261710 153237 261770 154670
rect 261707 153236 261773 153237
rect 261707 153172 261708 153236
rect 261772 153172 261773 153236
rect 261707 153171 261773 153172
rect 262814 153101 262874 154670
rect 262811 153100 262877 153101
rect 262811 153036 262812 153100
rect 262876 153036 262877 153100
rect 262811 153035 262877 153036
rect 260603 152692 260669 152693
rect 260603 152628 260604 152692
rect 260668 152628 260669 152692
rect 260603 152627 260669 152628
rect 258395 152556 258461 152557
rect 258395 152492 258396 152556
rect 258460 152492 258461 152556
rect 258395 152491 258461 152492
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 130308 258134 150618
rect 261234 137834 261854 153000
rect 263550 152421 263610 154670
rect 263918 154670 263996 154730
rect 265206 154670 265356 154730
rect 265942 154670 266036 154730
rect 266310 154670 266444 154730
rect 267598 154670 267668 154730
rect 263918 153101 263978 154670
rect 265206 153237 265266 154670
rect 265203 153236 265269 153237
rect 265203 153172 265204 153236
rect 265268 153172 265269 153236
rect 265203 153171 265269 153172
rect 263915 153100 263981 153101
rect 263915 153036 263916 153100
rect 263980 153036 263981 153100
rect 263915 153035 263981 153036
rect 263547 152420 263613 152421
rect 263547 152356 263548 152420
rect 263612 152356 263613 152420
rect 263547 152355 263613 152356
rect 261234 137598 261266 137834
rect 261502 137598 261586 137834
rect 261822 137598 261854 137834
rect 261234 137514 261854 137598
rect 261234 137278 261266 137514
rect 261502 137278 261586 137514
rect 261822 137278 261854 137514
rect 261234 130308 261854 137278
rect 264954 141554 265574 153000
rect 265942 152693 266002 154670
rect 266310 153101 266370 154670
rect 266307 153100 266373 153101
rect 266307 153036 266308 153100
rect 266372 153036 266373 153100
rect 266307 153035 266373 153036
rect 267598 152693 267658 154670
rect 268288 154590 268348 155040
rect 268696 154590 268756 155040
rect 269784 154590 269844 155040
rect 271008 154730 271068 155040
rect 270910 154670 271068 154730
rect 268288 154530 268394 154590
rect 268696 154530 268762 154590
rect 269784 154530 269866 154590
rect 268334 152693 268394 154530
rect 268702 153101 268762 154530
rect 269806 153101 269866 154530
rect 270910 153917 270970 154670
rect 271144 154590 271204 155040
rect 272232 154590 272292 155040
rect 273320 154590 273380 155040
rect 273592 154597 273652 155040
rect 271094 154530 271204 154590
rect 272198 154530 272292 154590
rect 273302 154530 273380 154590
rect 273589 154596 273655 154597
rect 273589 154532 273590 154596
rect 273654 154532 273655 154596
rect 274408 154590 274468 155040
rect 275768 154590 275828 155040
rect 273589 154531 273655 154532
rect 274406 154530 274468 154590
rect 275326 154530 275828 154590
rect 276040 154590 276100 155040
rect 276992 154590 277052 155040
rect 278080 154730 278140 155040
rect 277534 154670 278140 154730
rect 277534 154590 277594 154670
rect 278488 154590 278548 155040
rect 279168 154590 279228 155040
rect 280936 154590 280996 155040
rect 276040 154530 276306 154590
rect 270907 153916 270973 153917
rect 270907 153852 270908 153916
rect 270972 153852 270973 153916
rect 270907 153851 270973 153852
rect 271094 153101 271154 154530
rect 272198 153237 272258 154530
rect 272195 153236 272261 153237
rect 272195 153172 272196 153236
rect 272260 153172 272261 153236
rect 272195 153171 272261 153172
rect 268699 153100 268765 153101
rect 268699 153036 268700 153100
rect 268764 153036 268765 153100
rect 268699 153035 268765 153036
rect 269803 153100 269869 153101
rect 269803 153036 269804 153100
rect 269868 153036 269869 153100
rect 269803 153035 269869 153036
rect 271091 153100 271157 153101
rect 271091 153036 271092 153100
rect 271156 153036 271157 153100
rect 271091 153035 271157 153036
rect 265939 152692 266005 152693
rect 265939 152628 265940 152692
rect 266004 152628 266005 152692
rect 265939 152627 266005 152628
rect 267595 152692 267661 152693
rect 267595 152628 267596 152692
rect 267660 152628 267661 152692
rect 267595 152627 267661 152628
rect 268331 152692 268397 152693
rect 268331 152628 268332 152692
rect 268396 152628 268397 152692
rect 268331 152627 268397 152628
rect 264954 141318 264986 141554
rect 265222 141318 265306 141554
rect 265542 141318 265574 141554
rect 264954 141234 265574 141318
rect 264954 140998 264986 141234
rect 265222 140998 265306 141234
rect 265542 140998 265574 141234
rect 264954 130308 265574 140998
rect 271794 146514 272414 153000
rect 273302 152693 273362 154530
rect 274406 153101 274466 154530
rect 275326 153101 275386 154530
rect 274403 153100 274469 153101
rect 274403 153036 274404 153100
rect 274468 153036 274469 153100
rect 274403 153035 274469 153036
rect 275323 153100 275389 153101
rect 275323 153036 275324 153100
rect 275388 153036 275389 153100
rect 275323 153035 275389 153036
rect 273299 152692 273365 152693
rect 273299 152628 273300 152692
rect 273364 152628 273365 152692
rect 273299 152627 273365 152628
rect 271794 146278 271826 146514
rect 272062 146278 272146 146514
rect 272382 146278 272414 146514
rect 271794 146194 272414 146278
rect 271794 145958 271826 146194
rect 272062 145958 272146 146194
rect 272382 145958 272414 146194
rect 271794 130308 272414 145958
rect 275514 133174 276134 153000
rect 276246 152557 276306 154530
rect 276982 154530 277052 154590
rect 277166 154530 277594 154590
rect 278454 154530 278548 154590
rect 279006 154530 279228 154590
rect 280846 154530 280996 154590
rect 283520 154590 283580 155040
rect 285968 154590 286028 155040
rect 288280 154730 288340 155040
rect 291000 154730 291060 155040
rect 293448 154730 293508 155040
rect 288206 154670 288340 154730
rect 290966 154670 291060 154730
rect 293358 154670 293508 154730
rect 295896 154730 295956 155040
rect 298480 154730 298540 155040
rect 300928 154730 300988 155040
rect 303512 154730 303572 155040
rect 305960 154730 306020 155040
rect 295896 154670 295994 154730
rect 298480 154670 298570 154730
rect 283520 154530 283850 154590
rect 285968 154530 286058 154590
rect 276243 152556 276309 152557
rect 276243 152492 276244 152556
rect 276308 152492 276309 152556
rect 276243 152491 276309 152492
rect 276982 152013 277042 154530
rect 276979 152012 277045 152013
rect 276979 151948 276980 152012
rect 277044 151948 277045 152012
rect 277166 152010 277226 154530
rect 278454 153101 278514 154530
rect 279006 153101 279066 154530
rect 280846 153101 280906 154530
rect 283790 153101 283850 154530
rect 285998 153101 286058 154530
rect 288206 154189 288266 154670
rect 288203 154188 288269 154189
rect 288203 154124 288204 154188
rect 288268 154124 288269 154188
rect 288203 154123 288269 154124
rect 290966 153101 291026 154670
rect 293358 154189 293418 154670
rect 293355 154188 293421 154189
rect 293355 154124 293356 154188
rect 293420 154124 293421 154188
rect 293355 154123 293421 154124
rect 295934 153917 295994 154670
rect 298510 154053 298570 154670
rect 300902 154670 300988 154730
rect 303478 154670 303572 154730
rect 305870 154670 306020 154730
rect 298507 154052 298573 154053
rect 298507 153988 298508 154052
rect 298572 153988 298573 154052
rect 298507 153987 298573 153988
rect 295931 153916 295997 153917
rect 295931 153852 295932 153916
rect 295996 153852 295997 153916
rect 295931 153851 295997 153852
rect 300902 153237 300962 154670
rect 303478 154053 303538 154670
rect 305870 154189 305930 154670
rect 308544 154590 308604 155040
rect 308446 154530 308604 154590
rect 310992 154590 311052 155040
rect 313440 154590 313500 155040
rect 315888 154590 315948 155040
rect 310992 154530 311082 154590
rect 305867 154188 305933 154189
rect 305867 154124 305868 154188
rect 305932 154124 305933 154188
rect 305867 154123 305933 154124
rect 303475 154052 303541 154053
rect 303475 153988 303476 154052
rect 303540 153988 303541 154052
rect 303475 153987 303541 153988
rect 308446 153917 308506 154530
rect 308443 153916 308509 153917
rect 308443 153852 308444 153916
rect 308508 153852 308509 153916
rect 308443 153851 308509 153852
rect 300899 153236 300965 153237
rect 300899 153172 300900 153236
rect 300964 153172 300965 153236
rect 300899 153171 300965 153172
rect 278451 153100 278517 153101
rect 278451 153036 278452 153100
rect 278516 153036 278517 153100
rect 278451 153035 278517 153036
rect 279003 153100 279069 153101
rect 279003 153036 279004 153100
rect 279068 153036 279069 153100
rect 279003 153035 279069 153036
rect 280843 153100 280909 153101
rect 280843 153036 280844 153100
rect 280908 153036 280909 153100
rect 280843 153035 280909 153036
rect 283787 153100 283853 153101
rect 283787 153036 283788 153100
rect 283852 153036 283853 153100
rect 283787 153035 283853 153036
rect 285995 153100 286061 153101
rect 285995 153036 285996 153100
rect 286060 153036 286061 153100
rect 285995 153035 286061 153036
rect 290963 153100 291029 153101
rect 290963 153036 290964 153100
rect 291028 153036 291029 153100
rect 290963 153035 291029 153036
rect 277166 151950 277410 152010
rect 276979 151947 277045 151948
rect 277350 151877 277410 151950
rect 277347 151876 277413 151877
rect 277347 151812 277348 151876
rect 277412 151812 277413 151876
rect 277347 151811 277413 151812
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 130308 276134 132618
rect 279234 136894 279854 153000
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 130308 279854 136338
rect 282954 140614 283574 153000
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 130308 283574 140058
rect 289794 147454 290414 153000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 130308 290414 146898
rect 293514 151174 294134 153000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 130308 294134 150618
rect 297234 137834 297854 153000
rect 297234 137598 297266 137834
rect 297502 137598 297586 137834
rect 297822 137598 297854 137834
rect 297234 137514 297854 137598
rect 297234 137278 297266 137514
rect 297502 137278 297586 137514
rect 297822 137278 297854 137514
rect 297234 130308 297854 137278
rect 300954 141554 301574 153000
rect 300954 141318 300986 141554
rect 301222 141318 301306 141554
rect 301542 141318 301574 141554
rect 300954 141234 301574 141318
rect 300954 140998 300986 141234
rect 301222 140998 301306 141234
rect 301542 140998 301574 141234
rect 300954 130308 301574 140998
rect 307794 146514 308414 153000
rect 311022 152829 311082 154530
rect 313414 154530 313500 154590
rect 315806 154530 315948 154590
rect 313414 154325 313474 154530
rect 315806 154461 315866 154530
rect 315803 154460 315869 154461
rect 315803 154396 315804 154460
rect 315868 154396 315869 154460
rect 318472 154458 318532 155040
rect 315803 154395 315869 154396
rect 318382 154398 318532 154458
rect 320920 154458 320980 155040
rect 323368 154458 323428 155040
rect 325952 154730 326012 155040
rect 343224 154730 343284 155040
rect 320920 154398 321018 154458
rect 313411 154324 313477 154325
rect 313411 154260 313412 154324
rect 313476 154260 313477 154324
rect 313411 154259 313477 154260
rect 311019 152828 311085 152829
rect 311019 152764 311020 152828
rect 311084 152764 311085 152828
rect 311019 152763 311085 152764
rect 307794 146278 307826 146514
rect 308062 146278 308146 146514
rect 308382 146278 308414 146514
rect 307794 146194 308414 146278
rect 307794 145958 307826 146194
rect 308062 145958 308146 146194
rect 308382 145958 308414 146194
rect 307794 130308 308414 145958
rect 311514 133174 312134 153000
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 130308 312134 132618
rect 315234 136894 315854 153000
rect 318382 152965 318442 154398
rect 320958 153101 321018 154398
rect 322982 154398 323428 154458
rect 325742 154670 326012 154730
rect 343222 154670 343284 154730
rect 343360 154730 343420 155040
rect 343360 154670 343466 154730
rect 320955 153100 321021 153101
rect 320955 153036 320956 153100
rect 321020 153036 321021 153100
rect 320955 153035 321021 153036
rect 318379 152964 318445 152965
rect 318379 152900 318380 152964
rect 318444 152900 318445 152964
rect 318379 152899 318445 152900
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 130308 315854 136338
rect 318954 140614 319574 153000
rect 322982 151741 323042 154398
rect 325742 153370 325802 154670
rect 325558 153310 325802 153370
rect 325558 152149 325618 153310
rect 325555 152148 325621 152149
rect 325555 152084 325556 152148
rect 325620 152084 325621 152148
rect 325555 152083 325621 152084
rect 322979 151740 323045 151741
rect 322979 151676 322980 151740
rect 323044 151676 323045 151740
rect 322979 151675 323045 151676
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 130308 319574 140058
rect 325794 147454 326414 153000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 130308 326414 146898
rect 329514 151174 330134 153000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 130308 330134 150618
rect 333234 137834 333854 153000
rect 333234 137598 333266 137834
rect 333502 137598 333586 137834
rect 333822 137598 333854 137834
rect 333234 137514 333854 137598
rect 333234 137278 333266 137514
rect 333502 137278 333586 137514
rect 333822 137278 333854 137514
rect 333234 130308 333854 137278
rect 336954 141554 337574 153000
rect 343222 152829 343282 154670
rect 343219 152828 343285 152829
rect 343219 152764 343220 152828
rect 343284 152764 343285 152828
rect 343219 152763 343285 152764
rect 343406 152557 343466 154670
rect 343403 152556 343469 152557
rect 343403 152492 343404 152556
rect 343468 152492 343469 152556
rect 343403 152491 343469 152492
rect 336954 141318 336986 141554
rect 337222 141318 337306 141554
rect 337542 141318 337574 141554
rect 336954 141234 337574 141318
rect 336954 140998 336986 141234
rect 337222 140998 337306 141234
rect 337542 140998 337574 141234
rect 336954 130308 337574 140998
rect 343794 146514 344414 153000
rect 343794 146278 343826 146514
rect 344062 146278 344146 146514
rect 344382 146278 344414 146514
rect 343794 146194 344414 146278
rect 343794 145958 343826 146194
rect 344062 145958 344146 146194
rect 344382 145958 344414 146194
rect 343794 130308 344414 145958
rect 347514 133174 348134 153000
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 130308 348134 132618
rect 351234 136894 351854 153000
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 130308 351854 136338
rect 354954 140614 355574 153000
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 130308 355574 140058
rect 338435 129844 338501 129845
rect 338435 129780 338436 129844
rect 338500 129780 338501 129844
rect 338435 129779 338501 129780
rect 339723 129844 339789 129845
rect 339723 129780 339724 129844
rect 339788 129780 339789 129844
rect 339723 129779 339789 129780
rect 350947 129844 351013 129845
rect 350947 129780 350948 129844
rect 351012 129780 351013 129844
rect 350947 129779 351013 129780
rect 338438 128890 338498 129779
rect 339726 128890 339786 129779
rect 350950 128890 351010 129779
rect 338438 128830 338524 128890
rect 338464 128202 338524 128830
rect 339688 128830 339786 128890
rect 350840 128830 351010 128890
rect 339688 128202 339748 128830
rect 350840 128202 350900 128830
rect 220952 111454 221300 111486
rect 220952 111218 221008 111454
rect 221244 111218 221300 111454
rect 220952 111134 221300 111218
rect 220952 110898 221008 111134
rect 221244 110898 221300 111134
rect 220952 110866 221300 110898
rect 355320 111454 355668 111486
rect 355320 111218 355376 111454
rect 355612 111218 355668 111454
rect 355320 111134 355668 111218
rect 355320 110898 355376 111134
rect 355612 110898 355668 111134
rect 355320 110866 355668 110898
rect 220272 93454 220620 93486
rect 220272 93218 220328 93454
rect 220564 93218 220620 93454
rect 220272 93134 220620 93218
rect 220272 92898 220328 93134
rect 220564 92898 220620 93134
rect 220272 92866 220620 92898
rect 356000 93454 356348 93486
rect 356000 93218 356056 93454
rect 356292 93218 356348 93454
rect 356000 93134 356348 93218
rect 356000 92898 356056 93134
rect 356292 92898 356348 93134
rect 356000 92866 356348 92898
rect 220952 75454 221300 75486
rect 220952 75218 221008 75454
rect 221244 75218 221300 75454
rect 220952 75134 221300 75218
rect 220952 74898 221008 75134
rect 221244 74898 221300 75134
rect 220952 74866 221300 74898
rect 355320 75454 355668 75486
rect 355320 75218 355376 75454
rect 355612 75218 355668 75454
rect 355320 75134 355668 75218
rect 355320 74898 355376 75134
rect 355612 74898 355668 75134
rect 355320 74866 355668 74898
rect 220272 57454 220620 57486
rect 220272 57218 220328 57454
rect 220564 57218 220620 57454
rect 220272 57134 220620 57218
rect 220272 56898 220328 57134
rect 220564 56898 220620 57134
rect 220272 56866 220620 56898
rect 356000 57454 356348 57486
rect 356000 57218 356056 57454
rect 356292 57218 356348 57454
rect 356000 57134 356348 57218
rect 356000 56898 356056 57134
rect 356292 56898 356348 57134
rect 356000 56866 356348 56898
rect 236056 44845 236116 45106
rect 237144 44845 237204 45106
rect 236053 44844 236119 44845
rect 236053 44780 236054 44844
rect 236118 44780 236119 44844
rect 236053 44779 236119 44780
rect 237141 44844 237207 44845
rect 237141 44780 237142 44844
rect 237206 44780 237207 44844
rect 237141 44779 237207 44780
rect 238232 44570 238292 45106
rect 239592 44570 239652 45106
rect 238158 44510 238292 44570
rect 239262 44510 239652 44570
rect 240544 44570 240604 45106
rect 241768 44570 241828 45106
rect 243128 44845 243188 45106
rect 244216 44845 244276 45106
rect 243125 44844 243191 44845
rect 243125 44780 243126 44844
rect 243190 44780 243191 44844
rect 243125 44779 243191 44780
rect 244213 44844 244279 44845
rect 244213 44780 244214 44844
rect 244278 44780 244279 44844
rect 244213 44779 244279 44780
rect 245440 44570 245500 45106
rect 246528 44570 246588 45106
rect 240544 44510 240610 44570
rect 219939 41308 220005 41309
rect 219939 41244 219940 41308
rect 220004 41244 220005 41308
rect 219939 41243 220005 41244
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 43000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 43000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 43000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 43000
rect 238158 42805 238218 44510
rect 239262 42805 239322 44510
rect 238155 42804 238221 42805
rect 238155 42740 238156 42804
rect 238220 42740 238221 42804
rect 238155 42739 238221 42740
rect 239259 42804 239325 42805
rect 239259 42740 239260 42804
rect 239324 42740 239325 42804
rect 239259 42739 239325 42740
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 43000
rect 240550 42805 240610 44510
rect 241654 44510 241828 44570
rect 245334 44510 245500 44570
rect 246438 44510 246588 44570
rect 247616 44570 247676 45106
rect 248296 44570 248356 45106
rect 248704 44570 248764 45106
rect 247616 44510 247786 44570
rect 241654 42805 241714 44510
rect 240547 42804 240613 42805
rect 240547 42740 240548 42804
rect 240612 42740 240613 42804
rect 240547 42739 240613 42740
rect 241651 42804 241717 42805
rect 241651 42740 241652 42804
rect 241716 42740 241717 42804
rect 241651 42739 241717 42740
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 43000
rect 245334 42805 245394 44510
rect 246438 42805 246498 44510
rect 245331 42804 245397 42805
rect 245331 42740 245332 42804
rect 245396 42740 245397 42804
rect 245331 42739 245397 42740
rect 246435 42804 246501 42805
rect 246435 42740 246436 42804
rect 246500 42740 246501 42804
rect 246435 42739 246501 42740
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 43000
rect 247726 41853 247786 44510
rect 248278 44510 248356 44570
rect 248646 44510 248764 44570
rect 250064 44570 250124 45106
rect 250744 44709 250804 45106
rect 250741 44708 250807 44709
rect 250741 44644 250742 44708
rect 250806 44644 250807 44708
rect 251288 44706 251348 45106
rect 250741 44643 250807 44644
rect 251222 44646 251348 44706
rect 250064 44510 250178 44570
rect 248278 41989 248338 44510
rect 248646 41989 248706 44510
rect 250118 42805 250178 44510
rect 251222 42805 251282 44646
rect 252376 44570 252436 45106
rect 253464 44570 253524 45106
rect 252326 44510 252436 44570
rect 253430 44510 253524 44570
rect 253600 44570 253660 45106
rect 254552 44570 254612 45106
rect 255912 44709 255972 45106
rect 255909 44708 255975 44709
rect 255909 44644 255910 44708
rect 255974 44644 255975 44708
rect 255909 44643 255975 44644
rect 256048 44570 256108 45106
rect 257000 44709 257060 45106
rect 258088 44709 258148 45106
rect 256997 44708 257063 44709
rect 256997 44644 256998 44708
rect 257062 44644 257063 44708
rect 256997 44643 257063 44644
rect 258085 44708 258151 44709
rect 258085 44644 258086 44708
rect 258150 44644 258151 44708
rect 258085 44643 258151 44644
rect 258496 44573 258556 45106
rect 259448 44573 259508 45106
rect 260672 44573 260732 45106
rect 253600 44510 253674 44570
rect 250115 42804 250181 42805
rect 250115 42740 250116 42804
rect 250180 42740 250181 42804
rect 250115 42739 250181 42740
rect 251219 42804 251285 42805
rect 251219 42740 251220 42804
rect 251284 42740 251285 42804
rect 251219 42739 251285 42740
rect 252326 41989 252386 44510
rect 253430 42805 253490 44510
rect 253427 42804 253493 42805
rect 253427 42740 253428 42804
rect 253492 42740 253493 42804
rect 253427 42739 253493 42740
rect 253614 42125 253674 44510
rect 254534 44510 254612 44570
rect 256006 44510 256108 44570
rect 258493 44572 258559 44573
rect 253611 42124 253677 42125
rect 253611 42060 253612 42124
rect 253676 42060 253677 42124
rect 253611 42059 253677 42060
rect 248275 41988 248341 41989
rect 248275 41924 248276 41988
rect 248340 41924 248341 41988
rect 248275 41923 248341 41924
rect 248643 41988 248709 41989
rect 248643 41924 248644 41988
rect 248708 41924 248709 41988
rect 248643 41923 248709 41924
rect 252323 41988 252389 41989
rect 252323 41924 252324 41988
rect 252388 41924 252389 41988
rect 252323 41923 252389 41924
rect 247723 41852 247789 41853
rect 247723 41788 247724 41852
rect 247788 41788 247789 41852
rect 247723 41787 247789 41788
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 43000
rect 254534 42125 254594 44510
rect 256006 42261 256066 44510
rect 258493 44508 258494 44572
rect 258558 44508 258559 44572
rect 258493 44507 258559 44508
rect 259445 44572 259511 44573
rect 259445 44508 259446 44572
rect 259510 44508 259511 44572
rect 259445 44507 259511 44508
rect 260669 44572 260735 44573
rect 260669 44508 260670 44572
rect 260734 44508 260735 44572
rect 261080 44570 261140 45106
rect 261760 44573 261820 45106
rect 262848 44709 262908 45106
rect 262845 44708 262911 44709
rect 262845 44644 262846 44708
rect 262910 44644 262911 44708
rect 262845 44643 262911 44644
rect 260669 44507 260735 44508
rect 260974 44510 261140 44570
rect 261757 44572 261823 44573
rect 256003 42260 256069 42261
rect 256003 42196 256004 42260
rect 256068 42196 256069 42260
rect 256003 42195 256069 42196
rect 254531 42124 254597 42125
rect 254531 42060 254532 42124
rect 254596 42060 254597 42124
rect 254531 42059 254597 42060
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 43000
rect 260974 42805 261034 44510
rect 261757 44508 261758 44572
rect 261822 44508 261823 44572
rect 263528 44570 263588 45106
rect 263936 44573 263996 45106
rect 263933 44572 263999 44573
rect 263528 44510 263610 44570
rect 261757 44507 261823 44508
rect 260971 42804 261037 42805
rect 260971 42740 260972 42804
rect 261036 42740 261037 42804
rect 260971 42739 261037 42740
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 43000
rect 263550 42397 263610 44510
rect 263933 44508 263934 44572
rect 263998 44508 263999 44572
rect 265296 44570 265356 45106
rect 265976 44570 266036 45106
rect 266384 44570 266444 45106
rect 267608 44570 267668 45106
rect 263933 44507 263999 44508
rect 265206 44510 265356 44570
rect 265942 44510 266036 44570
rect 266310 44510 266444 44570
rect 267598 44510 267668 44570
rect 268288 44570 268348 45106
rect 268696 44570 268756 45106
rect 269784 44570 269844 45106
rect 271008 44570 271068 45106
rect 268288 44510 268394 44570
rect 268696 44510 268762 44570
rect 269784 44510 269866 44570
rect 265206 43213 265266 44510
rect 265942 43349 266002 44510
rect 265939 43348 266005 43349
rect 265939 43284 265940 43348
rect 266004 43284 266005 43348
rect 265939 43283 266005 43284
rect 265203 43212 265269 43213
rect 265203 43148 265204 43212
rect 265268 43148 265269 43212
rect 265203 43147 265269 43148
rect 263547 42396 263613 42397
rect 263547 42332 263548 42396
rect 263612 42332 263613 42396
rect 263547 42331 263613 42332
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 43000
rect 266310 42397 266370 44510
rect 267598 42397 267658 44510
rect 268334 42805 268394 44510
rect 268702 42805 268762 44510
rect 268331 42804 268397 42805
rect 268331 42740 268332 42804
rect 268396 42740 268397 42804
rect 268331 42739 268397 42740
rect 268699 42804 268765 42805
rect 268699 42740 268700 42804
rect 268764 42740 268765 42804
rect 268699 42739 268765 42740
rect 269806 42397 269866 44510
rect 270910 44510 271068 44570
rect 271144 44570 271204 45106
rect 272232 44570 272292 45106
rect 273320 44570 273380 45106
rect 273592 44570 273652 45106
rect 274408 44570 274468 45106
rect 275768 44570 275828 45106
rect 271144 44510 271338 44570
rect 270910 42533 270970 44510
rect 271278 42805 271338 44510
rect 272198 44510 272292 44570
rect 273302 44510 273380 44570
rect 273486 44510 273652 44570
rect 274406 44510 274468 44570
rect 275326 44510 275828 44570
rect 276040 44570 276100 45106
rect 276992 44570 277052 45106
rect 276040 44510 276306 44570
rect 272198 43213 272258 44510
rect 272195 43212 272261 43213
rect 272195 43148 272196 43212
rect 272260 43148 272261 43212
rect 272195 43147 272261 43148
rect 271275 42804 271341 42805
rect 271275 42740 271276 42804
rect 271340 42740 271341 42804
rect 271275 42739 271341 42740
rect 270907 42532 270973 42533
rect 270907 42468 270908 42532
rect 270972 42468 270973 42532
rect 270907 42467 270973 42468
rect 266307 42396 266373 42397
rect 266307 42332 266308 42396
rect 266372 42332 266373 42396
rect 266307 42331 266373 42332
rect 267595 42396 267661 42397
rect 267595 42332 267596 42396
rect 267660 42332 267661 42396
rect 267595 42331 267661 42332
rect 269803 42396 269869 42397
rect 269803 42332 269804 42396
rect 269868 42332 269869 42396
rect 269803 42331 269869 42332
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 43000
rect 273302 42805 273362 44510
rect 273486 43485 273546 44510
rect 273483 43484 273549 43485
rect 273483 43420 273484 43484
rect 273548 43420 273549 43484
rect 273483 43419 273549 43420
rect 273299 42804 273365 42805
rect 273299 42740 273300 42804
rect 273364 42740 273365 42804
rect 273299 42739 273365 42740
rect 274406 42261 274466 44510
rect 275326 42261 275386 44510
rect 274403 42260 274469 42261
rect 274403 42196 274404 42260
rect 274468 42196 274469 42260
rect 274403 42195 274469 42196
rect 275323 42260 275389 42261
rect 275323 42196 275324 42260
rect 275388 42196 275389 42260
rect 275323 42195 275389 42196
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 43000
rect 276246 42805 276306 44510
rect 276982 44510 277052 44570
rect 278080 44570 278140 45106
rect 278488 44570 278548 45106
rect 278080 44510 278146 44570
rect 276982 42805 277042 44510
rect 278086 42805 278146 44510
rect 278454 44510 278548 44570
rect 279168 44570 279228 45106
rect 280936 44570 280996 45106
rect 279168 44510 279250 44570
rect 278454 43757 278514 44510
rect 279190 43893 279250 44510
rect 280846 44510 280996 44570
rect 283520 44570 283580 45106
rect 285968 44570 286028 45106
rect 288280 44570 288340 45106
rect 291000 44570 291060 45106
rect 293448 44570 293508 45106
rect 283520 44510 283850 44570
rect 285968 44510 286058 44570
rect 279187 43892 279253 43893
rect 279187 43828 279188 43892
rect 279252 43828 279253 43892
rect 279187 43827 279253 43828
rect 278451 43756 278517 43757
rect 278451 43692 278452 43756
rect 278516 43692 278517 43756
rect 278451 43691 278517 43692
rect 280846 43621 280906 44510
rect 280843 43620 280909 43621
rect 280843 43556 280844 43620
rect 280908 43556 280909 43620
rect 280843 43555 280909 43556
rect 276243 42804 276309 42805
rect 276243 42740 276244 42804
rect 276308 42740 276309 42804
rect 276243 42739 276309 42740
rect 276979 42804 277045 42805
rect 276979 42740 276980 42804
rect 277044 42740 277045 42804
rect 276979 42739 277045 42740
rect 278083 42804 278149 42805
rect 278083 42740 278084 42804
rect 278148 42740 278149 42804
rect 278083 42739 278149 42740
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 43000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 43000
rect 283790 41717 283850 44510
rect 285998 43757 286058 44510
rect 288206 44510 288340 44570
rect 290966 44510 291060 44570
rect 293358 44510 293508 44570
rect 295896 44570 295956 45106
rect 298480 44570 298540 45106
rect 300928 44570 300988 45106
rect 303512 44570 303572 45106
rect 305960 44573 306020 45106
rect 308544 44573 308604 45106
rect 295896 44510 295994 44570
rect 298480 44510 298570 44570
rect 285995 43756 286061 43757
rect 285995 43692 285996 43756
rect 286060 43692 286061 43756
rect 285995 43691 286061 43692
rect 288206 42669 288266 44510
rect 290966 44029 291026 44510
rect 290963 44028 291029 44029
rect 290963 43964 290964 44028
rect 291028 43964 291029 44028
rect 290963 43963 291029 43964
rect 288203 42668 288269 42669
rect 288203 42604 288204 42668
rect 288268 42604 288269 42668
rect 288203 42603 288269 42604
rect 283787 41716 283853 41717
rect 283787 41652 283788 41716
rect 283852 41652 283853 41716
rect 283787 41651 283853 41652
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 43000
rect 293358 42805 293418 44510
rect 295934 44165 295994 44510
rect 295931 44164 295997 44165
rect 295931 44100 295932 44164
rect 295996 44100 295997 44164
rect 295931 44099 295997 44100
rect 293355 42804 293421 42805
rect 293355 42740 293356 42804
rect 293420 42740 293421 42804
rect 293355 42739 293421 42740
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 43000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 43000
rect 298510 42805 298570 44510
rect 300902 44510 300988 44570
rect 303478 44510 303572 44570
rect 305957 44572 306023 44573
rect 300902 44165 300962 44510
rect 300899 44164 300965 44165
rect 300899 44100 300900 44164
rect 300964 44100 300965 44164
rect 300899 44099 300965 44100
rect 298507 42804 298573 42805
rect 298507 42740 298508 42804
rect 298572 42740 298573 42804
rect 298507 42739 298573 42740
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 43000
rect 303478 42805 303538 44510
rect 305957 44508 305958 44572
rect 306022 44508 306023 44572
rect 305957 44507 306023 44508
rect 308541 44572 308607 44573
rect 308541 44508 308542 44572
rect 308606 44508 308607 44572
rect 310992 44570 311052 45106
rect 313440 44570 313500 45106
rect 315888 44709 315948 45106
rect 315885 44708 315951 44709
rect 315885 44644 315886 44708
rect 315950 44644 315951 44708
rect 318472 44706 318532 45106
rect 315885 44643 315951 44644
rect 318382 44646 318532 44706
rect 310992 44510 311082 44570
rect 308541 44507 308607 44508
rect 303475 42804 303541 42805
rect 303475 42740 303476 42804
rect 303540 42740 303541 42804
rect 303475 42739 303541 42740
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 43000
rect 311022 42805 311082 44510
rect 313414 44510 313500 44570
rect 311019 42804 311085 42805
rect 311019 42740 311020 42804
rect 311084 42740 311085 42804
rect 311019 42739 311085 42740
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 43000
rect 313414 42805 313474 44510
rect 313411 42804 313477 42805
rect 313411 42740 313412 42804
rect 313476 42740 313477 42804
rect 313411 42739 313477 42740
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 43000
rect 318382 42805 318442 44646
rect 320920 44570 320980 45106
rect 323368 44706 323428 45106
rect 323350 44646 323428 44706
rect 320920 44510 321018 44570
rect 318379 42804 318445 42805
rect 318379 42740 318380 42804
rect 318444 42740 318445 42804
rect 318379 42739 318445 42740
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 43000
rect 320958 42805 321018 44510
rect 323350 44301 323410 44646
rect 325952 44570 326012 45106
rect 343224 44570 343284 45106
rect 325926 44510 326012 44570
rect 343222 44510 343284 44570
rect 343360 44570 343420 45106
rect 343360 44510 343466 44570
rect 323347 44300 323413 44301
rect 323347 44236 323348 44300
rect 323412 44236 323413 44300
rect 323347 44235 323413 44236
rect 325926 43213 325986 44510
rect 325923 43212 325989 43213
rect 325923 43148 325924 43212
rect 325988 43148 325989 43212
rect 325923 43147 325989 43148
rect 320955 42804 321021 42805
rect 320955 42740 320956 42804
rect 321020 42740 321021 42804
rect 320955 42739 321021 42740
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 43000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 43000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 43000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 43000
rect 343222 42805 343282 44510
rect 343406 42805 343466 44510
rect 357942 44165 358002 492491
rect 360699 492420 360765 492421
rect 360699 492356 360700 492420
rect 360764 492356 360765 492420
rect 360699 492355 360765 492356
rect 359779 476780 359845 476781
rect 359779 476716 359780 476780
rect 359844 476716 359845 476780
rect 359779 476715 359845 476716
rect 359411 465764 359477 465765
rect 359411 465700 359412 465764
rect 359476 465700 359477 465764
rect 359411 465699 359477 465700
rect 359414 264893 359474 465699
rect 359595 462908 359661 462909
rect 359595 462844 359596 462908
rect 359660 462844 359661 462908
rect 359595 462843 359661 462844
rect 359411 264892 359477 264893
rect 359411 264828 359412 264892
rect 359476 264828 359477 264892
rect 359411 264827 359477 264828
rect 359598 264757 359658 462843
rect 359782 369069 359842 476715
rect 359963 471204 360029 471205
rect 359963 471140 359964 471204
rect 360028 471140 360029 471204
rect 359963 471139 360029 471140
rect 359966 371245 360026 471139
rect 359963 371244 360029 371245
rect 359963 371180 359964 371244
rect 360028 371180 360029 371244
rect 359963 371179 360029 371180
rect 359779 369068 359845 369069
rect 359779 369004 359780 369068
rect 359844 369004 359845 369068
rect 359779 369003 359845 369004
rect 359595 264756 359661 264757
rect 359595 264692 359596 264756
rect 359660 264692 359661 264756
rect 359595 264691 359661 264692
rect 360702 44301 360762 492355
rect 361794 471454 362414 506898
rect 365514 511174 366134 533000
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 364931 492284 364997 492285
rect 364931 492220 364932 492284
rect 364996 492220 364997 492284
rect 364931 492219 364997 492220
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 363459 467260 363525 467261
rect 363459 467196 363460 467260
rect 363524 467196 363525 467260
rect 363459 467195 363525 467196
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 360699 44300 360765 44301
rect 360699 44236 360700 44300
rect 360764 44236 360765 44300
rect 360699 44235 360765 44236
rect 357939 44164 358005 44165
rect 357939 44100 357940 44164
rect 358004 44100 358005 44164
rect 357939 44099 358005 44100
rect 343219 42804 343285 42805
rect 343219 42740 343220 42804
rect 343284 42740 343285 42804
rect 343219 42739 343285 42740
rect 343403 42804 343469 42805
rect 343403 42740 343404 42804
rect 343468 42740 343469 42804
rect 343403 42739 343469 42740
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 43000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 43000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 43000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 43000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 74898
rect 363462 42125 363522 467195
rect 364934 44029 364994 492219
rect 365514 475174 366134 510618
rect 369234 514894 369854 533000
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 367691 492148 367757 492149
rect 367691 492084 367692 492148
rect 367756 492084 367757 492148
rect 367691 492083 367757 492084
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 364931 44028 364997 44029
rect 364931 43964 364932 44028
rect 364996 43964 364997 44028
rect 364931 43963 364997 43964
rect 365514 43174 366134 78618
rect 367694 43893 367754 492083
rect 369234 478894 369854 514338
rect 372954 518614 373574 533000
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 371739 492012 371805 492013
rect 371739 491948 371740 492012
rect 371804 491948 371805 492012
rect 371739 491947 371805 491948
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 370451 478140 370517 478141
rect 370451 478076 370452 478140
rect 370516 478076 370517 478140
rect 370451 478075 370517 478076
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 137834 369854 154338
rect 369234 137598 369266 137834
rect 369502 137598 369586 137834
rect 369822 137598 369854 137834
rect 369234 137514 369854 137598
rect 369234 137278 369266 137514
rect 369502 137278 369586 137514
rect 369822 137278 369854 137514
rect 369234 118894 369854 137278
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 367691 43892 367757 43893
rect 367691 43828 367692 43892
rect 367756 43828 367757 43892
rect 367691 43827 367757 43828
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 363459 42124 363525 42125
rect 363459 42060 363460 42124
rect 363524 42060 363525 42124
rect 363459 42059 363525 42060
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 46338
rect 370454 42669 370514 478075
rect 371742 43621 371802 491947
rect 372954 482614 373574 518058
rect 379794 525454 380414 533000
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 374499 491876 374565 491877
rect 374499 491812 374500 491876
rect 374564 491812 374565 491876
rect 374499 491811 374565 491812
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 357554 373574 374058
rect 372954 357318 372986 357554
rect 373222 357318 373306 357554
rect 373542 357318 373574 357554
rect 372954 357234 373574 357318
rect 372954 356998 372986 357234
rect 373222 356998 373306 357234
rect 373542 356998 373574 357234
rect 372954 338614 373574 356998
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 249554 373574 266058
rect 372954 249318 372986 249554
rect 373222 249318 373306 249554
rect 373542 249318 373574 249554
rect 372954 249234 373574 249318
rect 372954 248998 372986 249234
rect 373222 248998 373306 249234
rect 373542 248998 373574 249234
rect 372954 230614 373574 248998
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 141554 373574 158058
rect 372954 141318 372986 141554
rect 373222 141318 373306 141554
rect 373542 141318 373574 141554
rect 372954 141234 373574 141318
rect 372954 140998 372986 141234
rect 373222 140998 373306 141234
rect 373542 140998 373574 141234
rect 372954 122614 373574 140998
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 371739 43620 371805 43621
rect 371739 43556 371740 43620
rect 371804 43556 371805 43620
rect 371739 43555 371805 43556
rect 370451 42668 370517 42669
rect 370451 42604 370452 42668
rect 370516 42604 370517 42668
rect 370451 42603 370517 42604
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 50058
rect 374502 43757 374562 491811
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 378179 487796 378245 487797
rect 378179 487732 378180 487796
rect 378244 487732 378245 487796
rect 378179 487731 378245 487732
rect 374683 483716 374749 483717
rect 374683 483652 374684 483716
rect 374748 483652 374749 483716
rect 374683 483651 374749 483652
rect 374499 43756 374565 43757
rect 374499 43692 374500 43756
rect 374564 43692 374565 43756
rect 374499 43691 374565 43692
rect 374686 42261 374746 483651
rect 375971 475420 376037 475421
rect 375971 475356 375972 475420
rect 376036 475356 376037 475420
rect 375971 475355 376037 475356
rect 374683 42260 374749 42261
rect 374683 42196 374684 42260
rect 374748 42196 374749 42260
rect 374683 42195 374749 42196
rect 375974 41989 376034 475355
rect 377259 474060 377325 474061
rect 377259 473996 377260 474060
rect 377324 473996 377325 474060
rect 377259 473995 377325 473996
rect 376155 472564 376221 472565
rect 376155 472500 376156 472564
rect 376220 472500 376221 472564
rect 376155 472499 376221 472500
rect 376158 42533 376218 472499
rect 376707 463044 376773 463045
rect 376707 462980 376708 463044
rect 376772 462980 376773 463044
rect 376707 462979 376773 462980
rect 376710 372741 376770 462979
rect 376891 460188 376957 460189
rect 376891 460124 376892 460188
rect 376956 460124 376957 460188
rect 376891 460123 376957 460124
rect 376894 373965 376954 460123
rect 376891 373964 376957 373965
rect 376891 373900 376892 373964
rect 376956 373900 376957 373964
rect 376891 373899 376957 373900
rect 376707 372740 376773 372741
rect 376707 372676 376708 372740
rect 376772 372676 376773 372740
rect 376707 372675 376773 372676
rect 376710 372469 376770 372675
rect 376707 372468 376773 372469
rect 376707 372404 376708 372468
rect 376772 372404 376773 372468
rect 376707 372403 376773 372404
rect 377262 371109 377322 473995
rect 377995 372740 378061 372741
rect 377995 372676 377996 372740
rect 378060 372676 378061 372740
rect 377995 372675 378061 372676
rect 377259 371108 377325 371109
rect 377259 371044 377260 371108
rect 377324 371044 377325 371108
rect 377259 371043 377325 371044
rect 377811 370428 377877 370429
rect 377811 370364 377812 370428
rect 377876 370364 377877 370428
rect 377811 370363 377877 370364
rect 377259 349756 377325 349757
rect 377259 349692 377260 349756
rect 377324 349692 377325 349756
rect 377259 349691 377325 349692
rect 377262 239869 377322 349691
rect 377814 260133 377874 370363
rect 377998 260949 378058 372675
rect 378182 262989 378242 487731
rect 378731 479500 378797 479501
rect 378731 479436 378732 479500
rect 378796 479436 378797 479500
rect 378731 479435 378797 479436
rect 378179 262988 378245 262989
rect 378179 262924 378180 262988
rect 378244 262924 378245 262988
rect 378179 262923 378245 262924
rect 377995 260948 378061 260949
rect 377995 260884 377996 260948
rect 378060 260884 378061 260948
rect 377995 260883 378061 260884
rect 377811 260132 377877 260133
rect 377811 260068 377812 260132
rect 377876 260068 377877 260132
rect 377811 260067 377877 260068
rect 377259 239868 377325 239869
rect 377259 239804 377260 239868
rect 377324 239804 377325 239868
rect 377259 239803 377325 239804
rect 377995 239460 378061 239461
rect 377995 239396 377996 239460
rect 378060 239396 378061 239460
rect 377995 239395 378061 239396
rect 377259 133788 377325 133789
rect 377259 133724 377260 133788
rect 377324 133724 377325 133788
rect 377259 133723 377325 133724
rect 376155 42532 376221 42533
rect 376155 42468 376156 42532
rect 376220 42468 376221 42532
rect 376155 42467 376221 42468
rect 375971 41988 376037 41989
rect 375971 41924 375972 41988
rect 376036 41924 376037 41988
rect 375971 41923 376037 41924
rect 377262 41037 377322 133723
rect 377811 133108 377877 133109
rect 377811 133044 377812 133108
rect 377876 133044 377877 133108
rect 377811 133043 377877 133044
rect 377814 41173 377874 133043
rect 377998 130933 378058 239395
rect 377995 130932 378061 130933
rect 377995 130868 377996 130932
rect 378060 130868 378061 130932
rect 377995 130867 378061 130868
rect 377998 129845 378058 130867
rect 377995 129844 378061 129845
rect 377995 129780 377996 129844
rect 378060 129780 378061 129844
rect 377995 129779 378061 129780
rect 378734 42397 378794 479435
rect 378915 467124 378981 467125
rect 378915 467060 378916 467124
rect 378980 467060 378981 467124
rect 378915 467059 378981 467060
rect 378731 42396 378797 42397
rect 378731 42332 378732 42396
rect 378796 42332 378797 42396
rect 378731 42331 378797 42332
rect 378918 41581 378978 467059
rect 379794 460308 380414 488898
rect 383514 529174 384134 533000
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 460308 384134 492618
rect 387234 532894 387854 533000
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460308 387854 496338
rect 390954 500614 391574 533000
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 460308 391574 464058
rect 397794 507454 398414 533000
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 460308 398414 470898
rect 401514 511174 402134 533000
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 460308 402134 474618
rect 405234 514894 405854 533000
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 460308 405854 478338
rect 408954 518614 409574 533000
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 460308 409574 482058
rect 415794 525454 416414 533000
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 460308 416414 488898
rect 419514 529174 420134 533000
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 460308 420134 492618
rect 423234 532894 423854 533000
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460308 423854 496338
rect 426954 500614 427574 533000
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 460308 427574 464058
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 460308 434414 470898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 460308 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 460308 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 460308 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 460308 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 637000 459854 640338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 637000 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 637000 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 637000 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 637000 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 637000 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 637000 488414 668898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637000 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 637000 495854 640338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 637000 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 637000 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 637000 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 479568 597454 479888 597486
rect 479568 597218 479610 597454
rect 479846 597218 479888 597454
rect 479568 597134 479888 597218
rect 479568 596898 479610 597134
rect 479846 596898 479888 597134
rect 479568 596866 479888 596898
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 460308 456134 492618
rect 459234 568894 459854 583000
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460308 459854 496338
rect 462954 572614 463574 583000
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 460308 463574 464058
rect 469794 579454 470414 583000
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 460308 470414 470898
rect 473514 547174 474134 583000
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 460308 474134 474618
rect 477234 550894 477854 583000
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 460308 477854 478338
rect 480954 554614 481574 583000
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 460308 481574 482058
rect 487794 561454 488414 583000
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 460308 488414 488898
rect 491514 565174 492134 583000
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 460308 492134 492618
rect 495234 568894 495854 583000
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460308 495854 496338
rect 498954 572614 499574 583000
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498515 461004 498581 461005
rect 498515 460940 498516 461004
rect 498580 460940 498581 461004
rect 498515 460939 498581 460940
rect 498518 458690 498578 460939
rect 498954 460308 499574 464058
rect 505794 579454 506414 583000
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 499803 461004 499869 461005
rect 499803 460940 499804 461004
rect 499868 460940 499869 461004
rect 499803 460939 499869 460940
rect 499806 458690 499866 460939
rect 505794 460308 506414 470898
rect 509514 547174 510134 583000
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 460308 510134 474618
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 510843 462228 510909 462229
rect 510843 462164 510844 462228
rect 510908 462164 510909 462228
rect 510843 462163 510909 462164
rect 510846 458690 510906 462163
rect 513234 460308 513854 478338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 460308 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 498464 458630 498578 458690
rect 499688 458630 499866 458690
rect 510840 458630 510906 458690
rect 498464 458202 498524 458630
rect 499688 458202 499748 458630
rect 510840 458202 510900 458630
rect 380272 453454 380620 453486
rect 380272 453218 380328 453454
rect 380564 453218 380620 453454
rect 380272 453134 380620 453218
rect 380272 452898 380328 453134
rect 380564 452898 380620 453134
rect 380272 452866 380620 452898
rect 516000 453454 516348 453486
rect 516000 453218 516056 453454
rect 516292 453218 516348 453454
rect 516000 453134 516348 453218
rect 516000 452898 516056 453134
rect 516292 452898 516348 453134
rect 516000 452866 516348 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 380952 435454 381300 435486
rect 380952 435218 381008 435454
rect 381244 435218 381300 435454
rect 380952 435134 381300 435218
rect 380952 434898 381008 435134
rect 381244 434898 381300 435134
rect 380952 434866 381300 434898
rect 515320 435454 515668 435486
rect 515320 435218 515376 435454
rect 515612 435218 515668 435454
rect 515320 435134 515668 435218
rect 515320 434898 515376 435134
rect 515612 434898 515668 435134
rect 515320 434866 515668 434898
rect 380272 417454 380620 417486
rect 380272 417218 380328 417454
rect 380564 417218 380620 417454
rect 380272 417134 380620 417218
rect 380272 416898 380328 417134
rect 380564 416898 380620 417134
rect 380272 416866 380620 416898
rect 516000 417454 516348 417486
rect 516000 417218 516056 417454
rect 516292 417218 516348 417454
rect 516000 417134 516348 417218
rect 516000 416898 516056 417134
rect 516292 416898 516348 417134
rect 516000 416866 516348 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 380952 399454 381300 399486
rect 380952 399218 381008 399454
rect 381244 399218 381300 399454
rect 380952 399134 381300 399218
rect 380952 398898 381008 399134
rect 381244 398898 381300 399134
rect 380952 398866 381300 398898
rect 515320 399454 515668 399486
rect 515320 399218 515376 399454
rect 515612 399218 515668 399454
rect 515320 399134 515668 399218
rect 515320 398898 515376 399134
rect 515612 398898 515668 399134
rect 515320 398866 515668 398898
rect 380272 381454 380620 381486
rect 380272 381218 380328 381454
rect 380564 381218 380620 381454
rect 380272 381134 380620 381218
rect 380272 380898 380328 381134
rect 380564 380898 380620 381134
rect 380272 380866 380620 380898
rect 516000 381454 516348 381486
rect 516000 381218 516056 381454
rect 516292 381218 516348 381454
rect 516000 381134 516348 381218
rect 516000 380898 516056 381134
rect 516292 380898 516348 381134
rect 516000 380866 516348 380898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 407803 375052 407869 375053
rect 396086 374990 396274 375050
rect 379467 369884 379533 369885
rect 379467 369820 379468 369884
rect 379532 369820 379533 369884
rect 379467 369819 379533 369820
rect 379470 364350 379530 369819
rect 379470 364290 379714 364350
rect 379654 240277 379714 364290
rect 379794 362514 380414 373000
rect 379794 362278 379826 362514
rect 380062 362278 380146 362514
rect 380382 362278 380414 362514
rect 379794 362194 380414 362278
rect 379794 361958 379826 362194
rect 380062 361958 380146 362194
rect 380382 361958 380414 362194
rect 379794 350308 380414 361958
rect 383514 366234 384134 373000
rect 383514 365998 383546 366234
rect 383782 365998 383866 366234
rect 384102 365998 384134 366234
rect 383514 365914 384134 365998
rect 383514 365678 383546 365914
rect 383782 365678 383866 365914
rect 384102 365678 384134 365914
rect 383514 350308 384134 365678
rect 387234 352894 387854 373000
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 350308 387854 352338
rect 390954 356614 391574 373000
rect 396214 372061 396274 374990
rect 396582 374990 397174 375050
rect 397502 374990 398262 375050
rect 398974 374990 399622 375050
rect 400262 374990 400574 375050
rect 401798 374990 402346 375050
rect 396211 372060 396277 372061
rect 396211 371996 396212 372060
rect 396276 371996 396277 372060
rect 396211 371995 396277 371996
rect 396582 371381 396642 374990
rect 397502 371925 397562 374990
rect 397499 371924 397565 371925
rect 397499 371860 397500 371924
rect 397564 371860 397565 371924
rect 397499 371859 397565 371860
rect 396579 371380 396645 371381
rect 396579 371316 396580 371380
rect 396644 371316 396645 371380
rect 396579 371315 396645 371316
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 350308 391574 356058
rect 397794 363454 398414 373000
rect 398974 372061 399034 374990
rect 400262 372197 400322 374990
rect 400259 372196 400325 372197
rect 400259 372132 400260 372196
rect 400324 372132 400325 372196
rect 400259 372131 400325 372132
rect 398971 372060 399037 372061
rect 398971 371996 398972 372060
rect 399036 371996 399037 372060
rect 398971 371995 399037 371996
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 350308 398414 362898
rect 401514 367174 402134 373000
rect 402286 371789 402346 374990
rect 403022 374990 403158 375050
rect 403574 374990 404246 375050
rect 404862 374990 405470 375050
rect 406150 374990 406558 375050
rect 407254 374990 407646 375050
rect 402283 371788 402349 371789
rect 402283 371724 402284 371788
rect 402348 371724 402349 371788
rect 402283 371723 402349 371724
rect 403022 371381 403082 374990
rect 403574 371381 403634 374990
rect 404862 373829 404922 374990
rect 404859 373828 404925 373829
rect 404859 373764 404860 373828
rect 404924 373764 404925 373828
rect 404859 373763 404925 373764
rect 403019 371380 403085 371381
rect 403019 371316 403020 371380
rect 403084 371316 403085 371380
rect 403019 371315 403085 371316
rect 403571 371380 403637 371381
rect 403571 371316 403572 371380
rect 403636 371316 403637 371380
rect 403571 371315 403637 371316
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 350308 402134 366618
rect 405234 370894 405854 373000
rect 406150 372197 406210 374990
rect 406147 372196 406213 372197
rect 406147 372132 406148 372196
rect 406212 372132 406213 372196
rect 406147 372131 406213 372132
rect 407254 371653 407314 374990
rect 407803 374988 407804 375052
rect 407868 375050 407869 375052
rect 418291 375052 418357 375053
rect 407868 374990 408326 375050
rect 408542 374990 408734 375050
rect 410014 374990 410094 375050
rect 407868 374988 407869 374990
rect 407803 374987 407869 374988
rect 407251 371652 407317 371653
rect 407251 371588 407252 371652
rect 407316 371588 407317 371652
rect 407251 371587 407317 371588
rect 408542 371381 408602 374990
rect 408539 371380 408605 371381
rect 408539 371316 408540 371380
rect 408604 371316 408605 371380
rect 408539 371315 408605 371316
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 350308 405854 370338
rect 408954 357554 409574 373000
rect 410014 371789 410074 374990
rect 410744 374645 410804 375020
rect 410741 374644 410807 374645
rect 410741 374580 410742 374644
rect 410806 374580 410807 374644
rect 410741 374579 410807 374580
rect 410011 371788 410077 371789
rect 410011 371724 410012 371788
rect 410076 371724 410077 371788
rect 410011 371723 410077 371724
rect 411302 371517 411362 375050
rect 411854 374990 412406 375050
rect 412774 374990 413494 375050
rect 413630 374990 413754 375050
rect 411854 371789 411914 374990
rect 411851 371788 411917 371789
rect 411851 371724 411852 371788
rect 411916 371724 411917 371788
rect 411851 371723 411917 371724
rect 412774 371653 412834 374990
rect 413694 371925 413754 374990
rect 414062 374990 414582 375050
rect 415718 374990 415942 375050
rect 416078 374990 416146 375050
rect 413691 371924 413757 371925
rect 413691 371860 413692 371924
rect 413756 371860 413757 371924
rect 413691 371859 413757 371860
rect 412771 371652 412837 371653
rect 412771 371588 412772 371652
rect 412836 371588 412837 371652
rect 412771 371587 412837 371588
rect 411299 371516 411365 371517
rect 411299 371452 411300 371516
rect 411364 371452 411365 371516
rect 411299 371451 411365 371452
rect 414062 371381 414122 374990
rect 415718 374237 415778 374990
rect 415715 374236 415781 374237
rect 415715 374172 415716 374236
rect 415780 374172 415781 374236
rect 415715 374171 415781 374172
rect 416086 374010 416146 374990
rect 415534 373950 416146 374010
rect 416822 374990 417030 375050
rect 415534 371381 415594 373950
rect 414059 371380 414125 371381
rect 414059 371316 414060 371380
rect 414124 371316 414125 371380
rect 414059 371315 414125 371316
rect 415531 371380 415597 371381
rect 415531 371316 415532 371380
rect 415596 371316 415597 371380
rect 415531 371315 415597 371316
rect 408954 357318 408986 357554
rect 409222 357318 409306 357554
rect 409542 357318 409574 357554
rect 408954 357234 409574 357318
rect 408954 356998 408986 357234
rect 409222 356998 409306 357234
rect 409542 356998 409574 357234
rect 408954 350308 409574 356998
rect 415794 362514 416414 373000
rect 416822 371381 416882 374990
rect 418110 371381 418170 375050
rect 418291 374988 418292 375052
rect 418356 375050 418357 375052
rect 440371 375052 440437 375053
rect 418356 374990 418526 375050
rect 418846 374990 419478 375050
rect 420318 374990 420702 375050
rect 418356 374988 418357 374990
rect 418291 374987 418357 374988
rect 418846 371517 418906 374990
rect 418843 371516 418909 371517
rect 418843 371452 418844 371516
rect 418908 371452 418909 371516
rect 418843 371451 418909 371452
rect 416819 371380 416885 371381
rect 416819 371316 416820 371380
rect 416884 371316 416885 371380
rect 416819 371315 416885 371316
rect 418107 371380 418173 371381
rect 418107 371316 418108 371380
rect 418172 371316 418173 371380
rect 418107 371315 418173 371316
rect 415794 362278 415826 362514
rect 416062 362278 416146 362514
rect 416382 362278 416414 362514
rect 415794 362194 416414 362278
rect 415794 361958 415826 362194
rect 416062 361958 416146 362194
rect 416382 361958 416414 362194
rect 415794 350308 416414 361958
rect 419514 366234 420134 373000
rect 420318 371381 420378 374990
rect 421054 373829 421114 375050
rect 421238 374990 421790 375050
rect 422342 374990 422878 375050
rect 423078 374990 423558 375050
rect 423966 374990 424058 375050
rect 421051 373828 421117 373829
rect 421051 373764 421052 373828
rect 421116 373764 421117 373828
rect 421051 373763 421117 373764
rect 421238 371381 421298 374990
rect 422342 371517 422402 374990
rect 423078 373829 423138 374990
rect 423075 373828 423141 373829
rect 423075 373764 423076 373828
rect 423140 373764 423141 373828
rect 423075 373763 423141 373764
rect 422339 371516 422405 371517
rect 422339 371452 422340 371516
rect 422404 371452 422405 371516
rect 422339 371451 422405 371452
rect 420315 371380 420381 371381
rect 420315 371316 420316 371380
rect 420380 371316 420381 371380
rect 420315 371315 420381 371316
rect 421235 371380 421301 371381
rect 421235 371316 421236 371380
rect 421300 371316 421301 371380
rect 421235 371315 421301 371316
rect 419514 365998 419546 366234
rect 419782 365998 419866 366234
rect 420102 365998 420134 366234
rect 419514 365914 420134 365998
rect 419514 365678 419546 365914
rect 419782 365678 419866 365914
rect 420102 365678 420134 365914
rect 419514 350308 420134 365678
rect 423234 352894 423854 373000
rect 423998 371381 424058 374990
rect 425286 372605 425346 375050
rect 425470 374990 426006 375050
rect 425470 373829 425530 374990
rect 425467 373828 425533 373829
rect 425467 373764 425468 373828
rect 425532 373764 425533 373828
rect 425467 373763 425533 373764
rect 426390 372605 426450 375050
rect 427638 374990 427738 375050
rect 425283 372604 425349 372605
rect 425283 372540 425284 372604
rect 425348 372540 425349 372604
rect 425283 372539 425349 372540
rect 426387 372604 426453 372605
rect 426387 372540 426388 372604
rect 426452 372540 426453 372604
rect 426387 372539 426453 372540
rect 423995 371380 424061 371381
rect 423995 371316 423996 371380
rect 424060 371316 424061 371380
rect 423995 371315 424061 371316
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 350308 423854 352338
rect 426954 356614 427574 373000
rect 427678 371517 427738 374990
rect 427862 374990 428318 375050
rect 428598 374990 428726 375050
rect 429334 374990 429814 375050
rect 430622 374990 431038 375050
rect 427675 371516 427741 371517
rect 427675 371452 427676 371516
rect 427740 371452 427741 371516
rect 427675 371451 427741 371452
rect 427862 371381 427922 374990
rect 428598 372605 428658 374990
rect 428595 372604 428661 372605
rect 428595 372540 428596 372604
rect 428660 372540 428661 372604
rect 428595 372539 428661 372540
rect 429334 371381 429394 374990
rect 430622 371789 430682 374990
rect 430619 371788 430685 371789
rect 430619 371724 430620 371788
rect 430684 371724 430685 371788
rect 430619 371723 430685 371724
rect 431174 371381 431234 375050
rect 432094 374990 432262 375050
rect 432094 371381 432154 374990
rect 433320 374509 433380 375020
rect 433592 374509 433652 375020
rect 433750 374990 434438 375050
rect 435222 374990 435798 375050
rect 433317 374508 433383 374509
rect 433317 374444 433318 374508
rect 433382 374444 433383 374508
rect 433317 374443 433383 374444
rect 433589 374508 433655 374509
rect 433589 374444 433590 374508
rect 433654 374444 433655 374508
rect 433589 374443 433655 374444
rect 433750 374010 433810 374990
rect 434851 374236 434917 374237
rect 434851 374172 434852 374236
rect 434916 374172 434917 374236
rect 434851 374171 434917 374172
rect 433566 373950 433810 374010
rect 433566 372469 433626 373950
rect 434854 373690 434914 374171
rect 435222 373965 435282 374990
rect 436040 374370 436100 375020
rect 435406 374310 436100 374370
rect 436326 374990 437022 375050
rect 438110 374990 438226 375050
rect 435219 373964 435285 373965
rect 435219 373900 435220 373964
rect 435284 373900 435285 373964
rect 435219 373899 435285 373900
rect 435406 373690 435466 374310
rect 434854 373630 435466 373690
rect 433563 372468 433629 372469
rect 433563 372404 433564 372468
rect 433628 372404 433629 372468
rect 433563 372403 433629 372404
rect 427859 371380 427925 371381
rect 427859 371316 427860 371380
rect 427924 371316 427925 371380
rect 427859 371315 427925 371316
rect 429331 371380 429397 371381
rect 429331 371316 429332 371380
rect 429396 371316 429397 371380
rect 429331 371315 429397 371316
rect 431171 371380 431237 371381
rect 431171 371316 431172 371380
rect 431236 371316 431237 371380
rect 431171 371315 431237 371316
rect 432091 371380 432157 371381
rect 432091 371316 432092 371380
rect 432156 371316 432157 371380
rect 432091 371315 432157 371316
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 350308 427574 356058
rect 433794 363454 434414 373000
rect 436326 371381 436386 374990
rect 438166 373149 438226 374990
rect 438350 374990 438518 375050
rect 439198 374990 439514 375050
rect 438163 373148 438229 373149
rect 438163 373084 438164 373148
rect 438228 373084 438229 373148
rect 438163 373083 438229 373084
rect 436323 371380 436389 371381
rect 436323 371316 436324 371380
rect 436388 371316 436389 371380
rect 436323 371315 436389 371316
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 350308 434414 362898
rect 437514 367174 438134 373000
rect 438350 371381 438410 374990
rect 439454 373829 439514 374990
rect 440371 374988 440372 375052
rect 440436 375050 440437 375052
rect 443131 375052 443197 375053
rect 440436 374990 440966 375050
rect 440436 374988 440437 374990
rect 440371 374987 440437 374988
rect 443131 374988 443132 375052
rect 443196 375050 443197 375052
rect 443196 374990 443550 375050
rect 443196 374988 443197 374990
rect 443131 374987 443197 374988
rect 445968 374509 446028 375020
rect 448280 374509 448340 375020
rect 450310 374990 451030 375050
rect 452886 374990 453478 375050
rect 455462 374990 455926 375050
rect 458222 374990 458510 375050
rect 460958 374990 461042 375050
rect 445965 374508 446031 374509
rect 445965 374444 445966 374508
rect 446030 374444 446031 374508
rect 445965 374443 446031 374444
rect 448277 374508 448343 374509
rect 448277 374444 448278 374508
rect 448342 374444 448343 374508
rect 448277 374443 448343 374444
rect 439451 373828 439517 373829
rect 439451 373764 439452 373828
rect 439516 373764 439517 373828
rect 439451 373763 439517 373764
rect 450310 373693 450370 374990
rect 450307 373692 450373 373693
rect 450307 373628 450308 373692
rect 450372 373628 450373 373692
rect 450307 373627 450373 373628
rect 452886 373557 452946 374990
rect 452883 373556 452949 373557
rect 452883 373492 452884 373556
rect 452948 373492 452949 373556
rect 452883 373491 452949 373492
rect 455462 373421 455522 374990
rect 458222 373557 458282 374990
rect 460982 373829 461042 374990
rect 462822 374990 463542 375050
rect 465398 374990 465990 375050
rect 467974 374990 468574 375050
rect 470734 374990 471022 375050
rect 473310 374990 473470 375050
rect 475334 374990 475918 375050
rect 478094 374990 478502 375050
rect 480302 374990 480950 375050
rect 483246 374990 483398 375050
rect 485822 374990 485982 375050
rect 503118 374990 503254 375050
rect 503390 374990 503546 375050
rect 460979 373828 461045 373829
rect 460979 373764 460980 373828
rect 461044 373764 461045 373828
rect 460979 373763 461045 373764
rect 462822 373557 462882 374990
rect 458219 373556 458285 373557
rect 458219 373492 458220 373556
rect 458284 373492 458285 373556
rect 458219 373491 458285 373492
rect 462819 373556 462885 373557
rect 462819 373492 462820 373556
rect 462884 373492 462885 373556
rect 462819 373491 462885 373492
rect 455459 373420 455525 373421
rect 455459 373356 455460 373420
rect 455524 373356 455525 373420
rect 455459 373355 455525 373356
rect 438347 371380 438413 371381
rect 438347 371316 438348 371380
rect 438412 371316 438413 371380
rect 438347 371315 438413 371316
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 350308 438134 366618
rect 441234 370894 441854 373000
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 350308 441854 370338
rect 444954 357554 445574 373000
rect 444954 357318 444986 357554
rect 445222 357318 445306 357554
rect 445542 357318 445574 357554
rect 444954 357234 445574 357318
rect 444954 356998 444986 357234
rect 445222 356998 445306 357234
rect 445542 356998 445574 357234
rect 444954 350308 445574 356998
rect 451794 362514 452414 373000
rect 451794 362278 451826 362514
rect 452062 362278 452146 362514
rect 452382 362278 452414 362514
rect 451794 362194 452414 362278
rect 451794 361958 451826 362194
rect 452062 361958 452146 362194
rect 452382 361958 452414 362194
rect 451794 350308 452414 361958
rect 455514 366234 456134 373000
rect 455514 365998 455546 366234
rect 455782 365998 455866 366234
rect 456102 365998 456134 366234
rect 455514 365914 456134 365998
rect 455514 365678 455546 365914
rect 455782 365678 455866 365914
rect 456102 365678 456134 365914
rect 455514 350308 456134 365678
rect 459234 352894 459854 373000
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 350308 459854 352338
rect 462954 356614 463574 373000
rect 465398 371653 465458 374990
rect 465395 371652 465461 371653
rect 465395 371588 465396 371652
rect 465460 371588 465461 371652
rect 465395 371587 465461 371588
rect 467974 371381 468034 374990
rect 467971 371380 468037 371381
rect 467971 371316 467972 371380
rect 468036 371316 468037 371380
rect 467971 371315 468037 371316
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 350308 463574 356058
rect 469794 363454 470414 373000
rect 470734 372333 470794 374990
rect 470731 372332 470797 372333
rect 470731 372268 470732 372332
rect 470796 372268 470797 372332
rect 470731 372267 470797 372268
rect 473310 371381 473370 374990
rect 473307 371380 473373 371381
rect 473307 371316 473308 371380
rect 473372 371316 473373 371380
rect 473307 371315 473373 371316
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 350308 470414 362898
rect 473514 367174 474134 373000
rect 475334 371245 475394 374990
rect 475331 371244 475397 371245
rect 475331 371180 475332 371244
rect 475396 371180 475397 371244
rect 475331 371179 475397 371180
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 350308 474134 366618
rect 477234 370894 477854 373000
rect 478094 371109 478154 374990
rect 480302 371381 480362 374990
rect 480299 371380 480365 371381
rect 480299 371316 480300 371380
rect 480364 371316 480365 371380
rect 480299 371315 480365 371316
rect 478091 371108 478157 371109
rect 478091 371044 478092 371108
rect 478156 371044 478157 371108
rect 478091 371043 478157 371044
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 350308 477854 370338
rect 480954 357554 481574 373000
rect 483246 371925 483306 374990
rect 483243 371924 483309 371925
rect 483243 371860 483244 371924
rect 483308 371860 483309 371924
rect 483243 371859 483309 371860
rect 485822 371381 485882 374990
rect 485819 371380 485885 371381
rect 485819 371316 485820 371380
rect 485884 371316 485885 371380
rect 485819 371315 485885 371316
rect 480954 357318 480986 357554
rect 481222 357318 481306 357554
rect 481542 357318 481574 357554
rect 480954 357234 481574 357318
rect 480954 356998 480986 357234
rect 481222 356998 481306 357234
rect 481542 356998 481574 357234
rect 480954 350308 481574 356998
rect 487794 362514 488414 373000
rect 487794 362278 487826 362514
rect 488062 362278 488146 362514
rect 488382 362278 488414 362514
rect 487794 362194 488414 362278
rect 487794 361958 487826 362194
rect 488062 361958 488146 362194
rect 488382 361958 488414 362194
rect 487794 350308 488414 361958
rect 491514 366234 492134 373000
rect 491514 365998 491546 366234
rect 491782 365998 491866 366234
rect 492102 365998 492134 366234
rect 491514 365914 492134 365998
rect 491514 365678 491546 365914
rect 491782 365678 491866 365914
rect 492102 365678 492134 365914
rect 491514 350308 492134 365678
rect 495234 352894 495854 373000
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 350308 495854 352338
rect 498954 356614 499574 373000
rect 503118 372197 503178 374990
rect 503115 372196 503181 372197
rect 503115 372132 503116 372196
rect 503180 372132 503181 372196
rect 503115 372131 503181 372132
rect 503486 371381 503546 374990
rect 503483 371380 503549 371381
rect 503483 371316 503484 371380
rect 503548 371316 503549 371380
rect 503483 371315 503549 371316
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498515 350572 498581 350573
rect 498515 350508 498516 350572
rect 498580 350508 498581 350572
rect 498515 350507 498581 350508
rect 498518 348530 498578 350507
rect 498954 350308 499574 356058
rect 505794 363454 506414 373000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 499803 350572 499869 350573
rect 499803 350508 499804 350572
rect 499868 350508 499869 350572
rect 499803 350507 499869 350508
rect 499806 348530 499866 350507
rect 505794 350308 506414 362898
rect 509514 367174 510134 373000
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 350308 510134 366618
rect 513234 370894 513854 373000
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 510843 350572 510909 350573
rect 510843 350508 510844 350572
rect 510908 350508 510909 350572
rect 510843 350507 510909 350508
rect 510846 348530 510906 350507
rect 513234 350308 513854 370338
rect 516954 357554 517574 373000
rect 516954 357318 516986 357554
rect 517222 357318 517306 357554
rect 517542 357318 517574 357554
rect 516954 357234 517574 357318
rect 516954 356998 516986 357234
rect 517222 356998 517306 357234
rect 517542 356998 517574 357234
rect 516954 350308 517574 356998
rect 498464 348470 498578 348530
rect 499688 348470 499866 348530
rect 510840 348470 510906 348530
rect 498464 348202 498524 348470
rect 499688 348202 499748 348470
rect 510840 348202 510900 348470
rect 380272 345454 380620 345486
rect 380272 345218 380328 345454
rect 380564 345218 380620 345454
rect 380272 345134 380620 345218
rect 380272 344898 380328 345134
rect 380564 344898 380620 345134
rect 380272 344866 380620 344898
rect 516000 345454 516348 345486
rect 516000 345218 516056 345454
rect 516292 345218 516348 345454
rect 516000 345134 516348 345218
rect 516000 344898 516056 345134
rect 516292 344898 516348 345134
rect 516000 344866 516348 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 380952 327454 381300 327486
rect 380952 327218 381008 327454
rect 381244 327218 381300 327454
rect 380952 327134 381300 327218
rect 380952 326898 381008 327134
rect 381244 326898 381300 327134
rect 380952 326866 381300 326898
rect 515320 327454 515668 327486
rect 515320 327218 515376 327454
rect 515612 327218 515668 327454
rect 515320 327134 515668 327218
rect 515320 326898 515376 327134
rect 515612 326898 515668 327134
rect 515320 326866 515668 326898
rect 380272 309454 380620 309486
rect 380272 309218 380328 309454
rect 380564 309218 380620 309454
rect 380272 309134 380620 309218
rect 380272 308898 380328 309134
rect 380564 308898 380620 309134
rect 380272 308866 380620 308898
rect 516000 309454 516348 309486
rect 516000 309218 516056 309454
rect 516292 309218 516348 309454
rect 516000 309134 516348 309218
rect 516000 308898 516056 309134
rect 516292 308898 516348 309134
rect 516000 308866 516348 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 380952 291454 381300 291486
rect 380952 291218 381008 291454
rect 381244 291218 381300 291454
rect 380952 291134 381300 291218
rect 380952 290898 381008 291134
rect 381244 290898 381300 291134
rect 380952 290866 381300 290898
rect 515320 291454 515668 291486
rect 515320 291218 515376 291454
rect 515612 291218 515668 291454
rect 515320 291134 515668 291218
rect 515320 290898 515376 291134
rect 515612 290898 515668 291134
rect 515320 290866 515668 290898
rect 380272 273454 380620 273486
rect 380272 273218 380328 273454
rect 380564 273218 380620 273454
rect 380272 273134 380620 273218
rect 380272 272898 380328 273134
rect 380564 272898 380620 273134
rect 380272 272866 380620 272898
rect 516000 273454 516348 273486
rect 516000 273218 516056 273454
rect 516292 273218 516348 273454
rect 516000 273134 516348 273218
rect 516000 272898 516056 273134
rect 516292 272898 516348 273134
rect 516000 272866 516348 272898
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 396056 264890 396116 265106
rect 397144 264890 397204 265106
rect 396030 264830 396116 264890
rect 397134 264830 397204 264890
rect 398232 264890 398292 265106
rect 399592 264890 399652 265106
rect 400544 264890 400604 265106
rect 401768 264890 401828 265106
rect 403128 264890 403188 265106
rect 404216 264890 404276 265106
rect 405440 264890 405500 265106
rect 406528 264890 406588 265106
rect 398232 264830 398298 264890
rect 379794 254514 380414 263000
rect 379794 254278 379826 254514
rect 380062 254278 380146 254514
rect 380382 254278 380414 254514
rect 379794 254194 380414 254278
rect 379794 253958 379826 254194
rect 380062 253958 380146 254194
rect 380382 253958 380414 254194
rect 379794 240308 380414 253958
rect 383514 241174 384134 263000
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 240308 384134 240618
rect 387234 244894 387854 263000
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 240308 387854 244338
rect 390954 248614 391574 263000
rect 396030 262309 396090 264830
rect 397134 262853 397194 264830
rect 398238 263533 398298 264830
rect 399526 264830 399652 264890
rect 400446 264830 400604 264890
rect 401734 264830 401828 264890
rect 403022 264830 403188 264890
rect 404126 264830 404276 264890
rect 405414 264830 405500 264890
rect 406518 264830 406588 264890
rect 407616 264890 407676 265106
rect 408296 264890 408356 265106
rect 408704 264890 408764 265106
rect 410064 264890 410124 265106
rect 407616 264830 407682 264890
rect 408296 264830 408418 264890
rect 408704 264830 408786 264890
rect 398235 263532 398301 263533
rect 398235 263468 398236 263532
rect 398300 263468 398301 263532
rect 398235 263467 398301 263468
rect 397131 262852 397197 262853
rect 397131 262788 397132 262852
rect 397196 262788 397197 262852
rect 397131 262787 397197 262788
rect 396027 262308 396093 262309
rect 396027 262244 396028 262308
rect 396092 262244 396093 262308
rect 396027 262243 396093 262244
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 240308 391574 248058
rect 397794 255454 398414 263000
rect 399526 262309 399586 264830
rect 400446 262309 400506 264830
rect 401734 263533 401794 264830
rect 401731 263532 401797 263533
rect 401731 263468 401732 263532
rect 401796 263468 401797 263532
rect 401731 263467 401797 263468
rect 399523 262308 399589 262309
rect 399523 262244 399524 262308
rect 399588 262244 399589 262308
rect 399523 262243 399589 262244
rect 400443 262308 400509 262309
rect 400443 262244 400444 262308
rect 400508 262244 400509 262308
rect 400443 262243 400509 262244
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 240308 398414 254898
rect 401514 259174 402134 263000
rect 403022 262309 403082 264830
rect 404126 262445 404186 264830
rect 405414 263533 405474 264830
rect 405411 263532 405477 263533
rect 405411 263468 405412 263532
rect 405476 263468 405477 263532
rect 405411 263467 405477 263468
rect 405234 262894 405854 263000
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 404123 262444 404189 262445
rect 404123 262380 404124 262444
rect 404188 262380 404189 262444
rect 404123 262379 404189 262380
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 403019 262308 403085 262309
rect 403019 262244 403020 262308
rect 403084 262244 403085 262308
rect 403019 262243 403085 262244
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 240308 402134 258618
rect 405234 240308 405854 262338
rect 406518 262309 406578 264830
rect 407622 262309 407682 264830
rect 408358 263533 408418 264830
rect 408355 263532 408421 263533
rect 408355 263468 408356 263532
rect 408420 263468 408421 263532
rect 408355 263467 408421 263468
rect 408726 262309 408786 264830
rect 410014 264830 410124 264890
rect 410744 264890 410804 265106
rect 411288 264890 411348 265106
rect 412376 264890 412436 265106
rect 413464 264890 413524 265106
rect 410744 264830 410810 264890
rect 411288 264830 411362 264890
rect 412376 264830 412466 264890
rect 406515 262308 406581 262309
rect 406515 262244 406516 262308
rect 406580 262244 406581 262308
rect 406515 262243 406581 262244
rect 407619 262308 407685 262309
rect 407619 262244 407620 262308
rect 407684 262244 407685 262308
rect 407619 262243 407685 262244
rect 408723 262308 408789 262309
rect 408723 262244 408724 262308
rect 408788 262244 408789 262308
rect 408723 262243 408789 262244
rect 408954 249554 409574 263000
rect 410014 262309 410074 264830
rect 410750 263533 410810 264830
rect 410747 263532 410813 263533
rect 410747 263468 410748 263532
rect 410812 263468 410813 263532
rect 410747 263467 410813 263468
rect 411302 262309 411362 264830
rect 412406 262445 412466 264830
rect 413326 264830 413524 264890
rect 413600 264890 413660 265106
rect 414552 264890 414612 265106
rect 415912 264890 415972 265106
rect 413600 264830 413754 264890
rect 414552 264830 414674 264890
rect 413326 262853 413386 264830
rect 413694 263533 413754 264830
rect 413691 263532 413757 263533
rect 413691 263468 413692 263532
rect 413756 263468 413757 263532
rect 413691 263467 413757 263468
rect 413323 262852 413389 262853
rect 413323 262788 413324 262852
rect 413388 262788 413389 262852
rect 413323 262787 413389 262788
rect 412403 262444 412469 262445
rect 412403 262380 412404 262444
rect 412468 262380 412469 262444
rect 412403 262379 412469 262380
rect 414614 262309 414674 264830
rect 415902 264830 415972 264890
rect 416048 264890 416108 265106
rect 417000 264890 417060 265106
rect 418088 264890 418148 265106
rect 416048 264830 416146 264890
rect 417000 264830 417066 264890
rect 418088 264830 418170 264890
rect 415902 263669 415962 264830
rect 415899 263668 415965 263669
rect 415899 263604 415900 263668
rect 415964 263604 415965 263668
rect 415899 263603 415965 263604
rect 416086 263533 416146 264830
rect 416083 263532 416149 263533
rect 416083 263468 416084 263532
rect 416148 263468 416149 263532
rect 416083 263467 416149 263468
rect 410011 262308 410077 262309
rect 410011 262244 410012 262308
rect 410076 262244 410077 262308
rect 410011 262243 410077 262244
rect 411299 262308 411365 262309
rect 411299 262244 411300 262308
rect 411364 262244 411365 262308
rect 411299 262243 411365 262244
rect 414611 262308 414677 262309
rect 414611 262244 414612 262308
rect 414676 262244 414677 262308
rect 414611 262243 414677 262244
rect 408954 249318 408986 249554
rect 409222 249318 409306 249554
rect 409542 249318 409574 249554
rect 408954 249234 409574 249318
rect 408954 248998 408986 249234
rect 409222 248998 409306 249234
rect 409542 248998 409574 249234
rect 408954 240308 409574 248998
rect 415794 254514 416414 263000
rect 417006 262309 417066 264830
rect 418110 262853 418170 264830
rect 418496 264621 418556 265106
rect 419448 264890 419508 265106
rect 419398 264830 419508 264890
rect 420672 264890 420732 265106
rect 420672 264830 420746 264890
rect 418493 264620 418559 264621
rect 418493 264556 418494 264620
rect 418558 264556 418559 264620
rect 418493 264555 418559 264556
rect 419398 263533 419458 264830
rect 419395 263532 419461 263533
rect 419395 263468 419396 263532
rect 419460 263468 419461 263532
rect 419395 263467 419461 263468
rect 418107 262852 418173 262853
rect 418107 262788 418108 262852
rect 418172 262788 418173 262852
rect 418107 262787 418173 262788
rect 417003 262308 417069 262309
rect 417003 262244 417004 262308
rect 417068 262244 417069 262308
rect 417003 262243 417069 262244
rect 415794 254278 415826 254514
rect 416062 254278 416146 254514
rect 416382 254278 416414 254514
rect 415794 254194 416414 254278
rect 415794 253958 415826 254194
rect 416062 253958 416146 254194
rect 416382 253958 416414 254194
rect 415794 240308 416414 253958
rect 419514 241174 420134 263000
rect 420686 262989 420746 264830
rect 421080 264621 421140 265106
rect 421760 264890 421820 265106
rect 422848 264890 422908 265106
rect 421760 264830 421850 264890
rect 422848 264830 422954 264890
rect 421077 264620 421143 264621
rect 421077 264556 421078 264620
rect 421142 264556 421143 264620
rect 421077 264555 421143 264556
rect 421790 262989 421850 264830
rect 420683 262988 420749 262989
rect 420683 262924 420684 262988
rect 420748 262924 420749 262988
rect 420683 262923 420749 262924
rect 421787 262988 421853 262989
rect 421787 262924 421788 262988
rect 421852 262924 421853 262988
rect 421787 262923 421853 262924
rect 422894 262309 422954 264830
rect 423528 264621 423588 265106
rect 423936 264890 423996 265106
rect 425296 264890 425356 265106
rect 423936 264830 424058 264890
rect 423525 264620 423591 264621
rect 423525 264556 423526 264620
rect 423590 264556 423591 264620
rect 423525 264555 423591 264556
rect 422891 262308 422957 262309
rect 422891 262244 422892 262308
rect 422956 262244 422957 262308
rect 422891 262243 422957 262244
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 240308 420134 240618
rect 423234 244894 423854 263000
rect 423998 262581 424058 264830
rect 425286 264830 425356 264890
rect 425286 263533 425346 264830
rect 425976 264621 426036 265106
rect 426384 264890 426444 265106
rect 427608 264890 427668 265106
rect 428288 264890 428348 265106
rect 428696 264890 428756 265106
rect 426384 264830 426450 264890
rect 425973 264620 426039 264621
rect 425973 264556 425974 264620
rect 426038 264556 426039 264620
rect 425973 264555 426039 264556
rect 426390 263533 426450 264830
rect 427494 264830 427668 264890
rect 428230 264830 428348 264890
rect 428598 264830 428756 264890
rect 427494 263533 427554 264830
rect 428230 263533 428290 264830
rect 425283 263532 425349 263533
rect 425283 263468 425284 263532
rect 425348 263468 425349 263532
rect 425283 263467 425349 263468
rect 426387 263532 426453 263533
rect 426387 263468 426388 263532
rect 426452 263468 426453 263532
rect 426387 263467 426453 263468
rect 427491 263532 427557 263533
rect 427491 263468 427492 263532
rect 427556 263468 427557 263532
rect 427491 263467 427557 263468
rect 428227 263532 428293 263533
rect 428227 263468 428228 263532
rect 428292 263468 428293 263532
rect 428227 263467 428293 263468
rect 423995 262580 424061 262581
rect 423995 262516 423996 262580
rect 424060 262516 424061 262580
rect 423995 262515 424061 262516
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 240308 423854 244338
rect 426954 248614 427574 263000
rect 428598 262309 428658 264830
rect 429784 264621 429844 265106
rect 431008 264890 431068 265106
rect 430990 264830 431068 264890
rect 431144 264890 431204 265106
rect 432232 264890 432292 265106
rect 433320 264890 433380 265106
rect 433592 264890 433652 265106
rect 431144 264830 431234 264890
rect 432232 264830 432338 264890
rect 433320 264830 433442 264890
rect 429781 264620 429847 264621
rect 429781 264556 429782 264620
rect 429846 264556 429847 264620
rect 429781 264555 429847 264556
rect 430990 263533 431050 264830
rect 430987 263532 431053 263533
rect 430987 263468 430988 263532
rect 431052 263468 431053 263532
rect 430987 263467 431053 263468
rect 431174 262309 431234 264830
rect 432278 263533 432338 264830
rect 433382 263533 433442 264830
rect 433566 264830 433652 264890
rect 434408 264890 434468 265106
rect 435768 264890 435828 265106
rect 436040 264890 436100 265106
rect 436992 264890 437052 265106
rect 434408 264830 434546 264890
rect 435768 264830 435834 264890
rect 432275 263532 432341 263533
rect 432275 263468 432276 263532
rect 432340 263468 432341 263532
rect 432275 263467 432341 263468
rect 433379 263532 433445 263533
rect 433379 263468 433380 263532
rect 433444 263468 433445 263532
rect 433379 263467 433445 263468
rect 433566 262989 433626 264830
rect 434486 263533 434546 264830
rect 434483 263532 434549 263533
rect 434483 263468 434484 263532
rect 434548 263468 434549 263532
rect 434483 263467 434549 263468
rect 433563 262988 433629 262989
rect 433563 262924 433564 262988
rect 433628 262924 433629 262988
rect 433563 262923 433629 262924
rect 428595 262308 428661 262309
rect 428595 262244 428596 262308
rect 428660 262244 428661 262308
rect 428595 262243 428661 262244
rect 431171 262308 431237 262309
rect 431171 262244 431172 262308
rect 431236 262244 431237 262308
rect 431171 262243 431237 262244
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 240308 427574 248058
rect 433794 255454 434414 263000
rect 435774 262989 435834 264830
rect 435958 264830 436100 264890
rect 436878 264830 437052 264890
rect 438080 264890 438140 265106
rect 438488 264890 438548 265106
rect 439168 264890 439228 265106
rect 440936 264890 440996 265106
rect 443520 264890 443580 265106
rect 438080 264830 438226 264890
rect 438488 264830 438594 264890
rect 439168 264830 439330 264890
rect 435958 263533 436018 264830
rect 435955 263532 436021 263533
rect 435955 263468 435956 263532
rect 436020 263468 436021 263532
rect 435955 263467 436021 263468
rect 435771 262988 435837 262989
rect 435771 262924 435772 262988
rect 435836 262924 435837 262988
rect 435771 262923 435837 262924
rect 436878 262309 436938 264830
rect 438166 263533 438226 264830
rect 438163 263532 438229 263533
rect 438163 263468 438164 263532
rect 438228 263468 438229 263532
rect 438163 263467 438229 263468
rect 436875 262308 436941 262309
rect 436875 262244 436876 262308
rect 436940 262244 436941 262308
rect 436875 262243 436941 262244
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 240308 434414 254898
rect 437514 259174 438134 263000
rect 438534 262989 438594 264830
rect 438531 262988 438597 262989
rect 438531 262924 438532 262988
rect 438596 262924 438597 262988
rect 438531 262923 438597 262924
rect 439270 262309 439330 264830
rect 440926 264830 440996 264890
rect 443502 264830 443580 264890
rect 440926 263533 440986 264830
rect 443502 263533 443562 264830
rect 445968 264757 446028 265106
rect 448280 264890 448340 265106
rect 451000 264890 451060 265106
rect 453448 264890 453508 265106
rect 455896 264890 455956 265106
rect 458480 264890 458540 265106
rect 448280 264830 448346 264890
rect 451000 264830 451106 264890
rect 445965 264756 446031 264757
rect 445965 264692 445966 264756
rect 446030 264692 446031 264756
rect 445965 264691 446031 264692
rect 448286 263533 448346 264830
rect 451046 263533 451106 264830
rect 453438 264830 453508 264890
rect 455830 264830 455956 264890
rect 458406 264830 458540 264890
rect 460928 264890 460988 265106
rect 463512 264890 463572 265106
rect 465960 264890 466020 265106
rect 460928 264830 461042 264890
rect 463512 264830 463618 264890
rect 453438 263533 453498 264830
rect 455830 263533 455890 264830
rect 440923 263532 440989 263533
rect 440923 263468 440924 263532
rect 440988 263468 440989 263532
rect 440923 263467 440989 263468
rect 443499 263532 443565 263533
rect 443499 263468 443500 263532
rect 443564 263468 443565 263532
rect 443499 263467 443565 263468
rect 448283 263532 448349 263533
rect 448283 263468 448284 263532
rect 448348 263468 448349 263532
rect 448283 263467 448349 263468
rect 451043 263532 451109 263533
rect 451043 263468 451044 263532
rect 451108 263468 451109 263532
rect 451043 263467 451109 263468
rect 453435 263532 453501 263533
rect 453435 263468 453436 263532
rect 453500 263468 453501 263532
rect 453435 263467 453501 263468
rect 455827 263532 455893 263533
rect 455827 263468 455828 263532
rect 455892 263468 455893 263532
rect 455827 263467 455893 263468
rect 441234 262894 441854 263000
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 439267 262308 439333 262309
rect 439267 262244 439268 262308
rect 439332 262244 439333 262308
rect 439267 262243 439333 262244
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 240308 438134 258618
rect 441234 240308 441854 262338
rect 444954 249554 445574 263000
rect 444954 249318 444986 249554
rect 445222 249318 445306 249554
rect 445542 249318 445574 249554
rect 444954 249234 445574 249318
rect 444954 248998 444986 249234
rect 445222 248998 445306 249234
rect 445542 248998 445574 249234
rect 444954 240308 445574 248998
rect 451794 254514 452414 263000
rect 451794 254278 451826 254514
rect 452062 254278 452146 254514
rect 452382 254278 452414 254514
rect 451794 254194 452414 254278
rect 451794 253958 451826 254194
rect 452062 253958 452146 254194
rect 452382 253958 452414 254194
rect 451794 240308 452414 253958
rect 455514 241174 456134 263000
rect 458406 262717 458466 264830
rect 460982 263125 461042 264830
rect 463558 263397 463618 264830
rect 465950 264830 466020 264890
rect 463555 263396 463621 263397
rect 463555 263332 463556 263396
rect 463620 263332 463621 263396
rect 463555 263331 463621 263332
rect 465950 263261 466010 264830
rect 468544 264757 468604 265106
rect 470992 264757 471052 265106
rect 473440 264893 473500 265106
rect 473437 264892 473503 264893
rect 473437 264828 473438 264892
rect 473502 264828 473503 264892
rect 473437 264827 473503 264828
rect 468541 264756 468607 264757
rect 468541 264692 468542 264756
rect 468606 264692 468607 264756
rect 468541 264691 468607 264692
rect 470989 264756 471055 264757
rect 470989 264692 470990 264756
rect 471054 264692 471055 264756
rect 470989 264691 471055 264692
rect 475888 264621 475948 265106
rect 478472 264757 478532 265106
rect 480920 264893 480980 265106
rect 480917 264892 480983 264893
rect 480917 264828 480918 264892
rect 480982 264828 480983 264892
rect 480917 264827 480983 264828
rect 483368 264757 483428 265106
rect 485952 264757 486012 265106
rect 503224 264890 503284 265106
rect 503118 264830 503284 264890
rect 503360 264890 503420 265106
rect 503360 264830 503546 264890
rect 478469 264756 478535 264757
rect 478469 264692 478470 264756
rect 478534 264692 478535 264756
rect 478469 264691 478535 264692
rect 483365 264756 483431 264757
rect 483365 264692 483366 264756
rect 483430 264692 483431 264756
rect 483365 264691 483431 264692
rect 485949 264756 486015 264757
rect 485949 264692 485950 264756
rect 486014 264692 486015 264756
rect 485949 264691 486015 264692
rect 475885 264620 475951 264621
rect 475885 264556 475886 264620
rect 475950 264556 475951 264620
rect 475885 264555 475951 264556
rect 465947 263260 466013 263261
rect 465947 263196 465948 263260
rect 466012 263196 466013 263260
rect 465947 263195 466013 263196
rect 460979 263124 461045 263125
rect 460979 263060 460980 263124
rect 461044 263060 461045 263124
rect 460979 263059 461045 263060
rect 458403 262716 458469 262717
rect 458403 262652 458404 262716
rect 458468 262652 458469 262716
rect 458403 262651 458469 262652
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 240308 456134 240618
rect 459234 244894 459854 263000
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 240308 459854 244338
rect 462954 248614 463574 263000
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 240308 463574 248058
rect 469794 255454 470414 263000
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 240308 470414 254898
rect 473514 259174 474134 263000
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 240308 474134 258618
rect 477234 262894 477854 263000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 240308 477854 262338
rect 480954 249554 481574 263000
rect 480954 249318 480986 249554
rect 481222 249318 481306 249554
rect 481542 249318 481574 249554
rect 480954 249234 481574 249318
rect 480954 248998 480986 249234
rect 481222 248998 481306 249234
rect 481542 248998 481574 249234
rect 480954 240308 481574 248998
rect 487794 254514 488414 263000
rect 487794 254278 487826 254514
rect 488062 254278 488146 254514
rect 488382 254278 488414 254514
rect 487794 254194 488414 254278
rect 487794 253958 487826 254194
rect 488062 253958 488146 254194
rect 488382 253958 488414 254194
rect 487794 240308 488414 253958
rect 491514 241174 492134 263000
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 240308 492134 240618
rect 495234 244894 495854 263000
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 240308 495854 244338
rect 498954 248614 499574 263000
rect 503118 262309 503178 264830
rect 503486 263533 503546 264830
rect 503483 263532 503549 263533
rect 503483 263468 503484 263532
rect 503548 263468 503549 263532
rect 503483 263467 503549 263468
rect 503115 262308 503181 262309
rect 503115 262244 503116 262308
rect 503180 262244 503181 262308
rect 503115 262243 503181 262244
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 240308 499574 248058
rect 505794 255454 506414 263000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 240308 506414 254898
rect 509514 259174 510134 263000
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 240308 510134 258618
rect 513234 262894 513854 263000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 510843 241500 510909 241501
rect 510843 241436 510844 241500
rect 510908 241436 510909 241500
rect 510843 241435 510909 241436
rect 379651 240276 379717 240277
rect 379651 240212 379652 240276
rect 379716 240212 379717 240276
rect 379651 240211 379717 240212
rect 498515 240276 498581 240277
rect 498515 240212 498516 240276
rect 498580 240212 498581 240276
rect 498515 240211 498581 240212
rect 499803 240276 499869 240277
rect 499803 240212 499804 240276
rect 499868 240212 499869 240276
rect 499803 240211 499869 240212
rect 379651 239596 379717 239597
rect 379651 239532 379652 239596
rect 379716 239532 379717 239596
rect 379651 239531 379717 239532
rect 379467 151332 379533 151333
rect 379467 151268 379468 151332
rect 379532 151330 379533 151332
rect 379654 151330 379714 239531
rect 498518 238770 498578 240211
rect 499806 238770 499866 240211
rect 510846 238770 510906 241435
rect 513234 240308 513854 262338
rect 516954 249554 517574 263000
rect 516954 249318 516986 249554
rect 517222 249318 517306 249554
rect 517542 249318 517574 249554
rect 516954 249234 517574 249318
rect 516954 248998 516986 249234
rect 517222 248998 517306 249234
rect 517542 248998 517574 249234
rect 516954 240308 517574 248998
rect 498464 238710 498578 238770
rect 499688 238710 499866 238770
rect 510840 238710 510906 238770
rect 498464 238202 498524 238710
rect 499688 238202 499748 238710
rect 510840 238202 510900 238710
rect 380272 237454 380620 237486
rect 380272 237218 380328 237454
rect 380564 237218 380620 237454
rect 380272 237134 380620 237218
rect 380272 236898 380328 237134
rect 380564 236898 380620 237134
rect 380272 236866 380620 236898
rect 516000 237454 516348 237486
rect 516000 237218 516056 237454
rect 516292 237218 516348 237454
rect 516000 237134 516348 237218
rect 516000 236898 516056 237134
rect 516292 236898 516348 237134
rect 516000 236866 516348 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 380952 219454 381300 219486
rect 380952 219218 381008 219454
rect 381244 219218 381300 219454
rect 380952 219134 381300 219218
rect 380952 218898 381008 219134
rect 381244 218898 381300 219134
rect 380952 218866 381300 218898
rect 515320 219454 515668 219486
rect 515320 219218 515376 219454
rect 515612 219218 515668 219454
rect 515320 219134 515668 219218
rect 515320 218898 515376 219134
rect 515612 218898 515668 219134
rect 515320 218866 515668 218898
rect 380272 201454 380620 201486
rect 380272 201218 380328 201454
rect 380564 201218 380620 201454
rect 380272 201134 380620 201218
rect 380272 200898 380328 201134
rect 380564 200898 380620 201134
rect 380272 200866 380620 200898
rect 516000 201454 516348 201486
rect 516000 201218 516056 201454
rect 516292 201218 516348 201454
rect 516000 201134 516348 201218
rect 516000 200898 516056 201134
rect 516292 200898 516348 201134
rect 516000 200866 516348 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 380952 183454 381300 183486
rect 380952 183218 381008 183454
rect 381244 183218 381300 183454
rect 380952 183134 381300 183218
rect 380952 182898 381008 183134
rect 381244 182898 381300 183134
rect 380952 182866 381300 182898
rect 515320 183454 515668 183486
rect 515320 183218 515376 183454
rect 515612 183218 515668 183454
rect 515320 183134 515668 183218
rect 515320 182898 515376 183134
rect 515612 182898 515668 183134
rect 515320 182866 515668 182898
rect 380272 165454 380620 165486
rect 380272 165218 380328 165454
rect 380564 165218 380620 165454
rect 380272 165134 380620 165218
rect 380272 164898 380328 165134
rect 380564 164898 380620 165134
rect 380272 164866 380620 164898
rect 516000 165454 516348 165486
rect 516000 165218 516056 165454
rect 516292 165218 516348 165454
rect 516000 165134 516348 165218
rect 516000 164898 516056 165134
rect 516292 164898 516348 165134
rect 516000 164866 516348 164898
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 396056 154590 396116 155040
rect 397144 154590 397204 155040
rect 396030 154530 396116 154590
rect 397134 154530 397204 154590
rect 398232 154590 398292 155040
rect 399592 154590 399652 155040
rect 400544 154590 400604 155040
rect 401768 154590 401828 155040
rect 403128 154590 403188 155040
rect 404216 154590 404276 155040
rect 405440 154590 405500 155040
rect 406528 154590 406588 155040
rect 398232 154530 398298 154590
rect 396030 153101 396090 154530
rect 396027 153100 396093 153101
rect 396027 153036 396028 153100
rect 396092 153036 396093 153100
rect 396027 153035 396093 153036
rect 379532 151270 379714 151330
rect 379532 151268 379533 151270
rect 379467 151267 379533 151268
rect 379654 45570 379714 151270
rect 379794 146514 380414 153000
rect 379794 146278 379826 146514
rect 380062 146278 380146 146514
rect 380382 146278 380414 146514
rect 379794 146194 380414 146278
rect 379794 145958 379826 146194
rect 380062 145958 380146 146194
rect 380382 145958 380414 146194
rect 379794 130308 380414 145958
rect 383514 133174 384134 153000
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 130308 384134 132618
rect 387234 136894 387854 153000
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 130308 387854 136338
rect 390954 140614 391574 153000
rect 397134 152557 397194 154530
rect 398238 153237 398298 154530
rect 399526 154530 399652 154590
rect 400446 154530 400604 154590
rect 401734 154530 401828 154590
rect 403022 154530 403188 154590
rect 404126 154530 404276 154590
rect 405046 154530 405500 154590
rect 406518 154530 406588 154590
rect 407616 154590 407676 155040
rect 408296 154590 408356 155040
rect 407616 154530 407682 154590
rect 398235 153236 398301 153237
rect 398235 153172 398236 153236
rect 398300 153172 398301 153236
rect 398235 153171 398301 153172
rect 399526 153101 399586 154530
rect 400446 153101 400506 154530
rect 401734 153237 401794 154530
rect 401731 153236 401797 153237
rect 401731 153172 401732 153236
rect 401796 153172 401797 153236
rect 401731 153171 401797 153172
rect 403022 153101 403082 154530
rect 399523 153100 399589 153101
rect 399523 153036 399524 153100
rect 399588 153036 399589 153100
rect 399523 153035 399589 153036
rect 400443 153100 400509 153101
rect 400443 153036 400444 153100
rect 400508 153036 400509 153100
rect 400443 153035 400509 153036
rect 403019 153100 403085 153101
rect 403019 153036 403020 153100
rect 403084 153036 403085 153100
rect 403019 153035 403085 153036
rect 397131 152556 397197 152557
rect 397131 152492 397132 152556
rect 397196 152492 397197 152556
rect 397131 152491 397197 152492
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 130308 391574 140058
rect 397794 147454 398414 153000
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 130308 398414 146898
rect 401514 151174 402134 153000
rect 404126 152557 404186 154530
rect 405046 153101 405106 154530
rect 406518 153101 406578 154530
rect 407622 153101 407682 154530
rect 408174 154530 408356 154590
rect 408704 154590 408764 155040
rect 410064 154590 410124 155040
rect 408704 154530 408786 154590
rect 405043 153100 405109 153101
rect 405043 153036 405044 153100
rect 405108 153036 405109 153100
rect 405043 153035 405109 153036
rect 406515 153100 406581 153101
rect 406515 153036 406516 153100
rect 406580 153036 406581 153100
rect 406515 153035 406581 153036
rect 407619 153100 407685 153101
rect 407619 153036 407620 153100
rect 407684 153036 407685 153100
rect 407619 153035 407685 153036
rect 404123 152556 404189 152557
rect 404123 152492 404124 152556
rect 404188 152492 404189 152556
rect 404123 152491 404189 152492
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 130308 402134 150618
rect 405234 137834 405854 153000
rect 408174 152421 408234 154530
rect 408726 153101 408786 154530
rect 410014 154530 410124 154590
rect 410744 154590 410804 155040
rect 411288 154590 411348 155040
rect 412376 154590 412436 155040
rect 413464 154590 413524 155040
rect 413600 154730 413660 155040
rect 413600 154670 413754 154730
rect 410744 154530 410810 154590
rect 411288 154530 411362 154590
rect 412376 154530 412466 154590
rect 413464 154530 413570 154590
rect 410014 153101 410074 154530
rect 408723 153100 408789 153101
rect 408723 153036 408724 153100
rect 408788 153036 408789 153100
rect 408723 153035 408789 153036
rect 410011 153100 410077 153101
rect 410011 153036 410012 153100
rect 410076 153036 410077 153100
rect 410011 153035 410077 153036
rect 408171 152420 408237 152421
rect 408171 152356 408172 152420
rect 408236 152356 408237 152420
rect 408171 152355 408237 152356
rect 405234 137598 405266 137834
rect 405502 137598 405586 137834
rect 405822 137598 405854 137834
rect 405234 137514 405854 137598
rect 405234 137278 405266 137514
rect 405502 137278 405586 137514
rect 405822 137278 405854 137514
rect 405234 130308 405854 137278
rect 408954 141554 409574 153000
rect 410750 152557 410810 154530
rect 411302 153101 411362 154530
rect 411299 153100 411365 153101
rect 411299 153036 411300 153100
rect 411364 153036 411365 153100
rect 411299 153035 411365 153036
rect 412406 152557 412466 154530
rect 413510 153101 413570 154530
rect 413507 153100 413573 153101
rect 413507 153036 413508 153100
rect 413572 153036 413573 153100
rect 413507 153035 413573 153036
rect 413694 152557 413754 154670
rect 414552 154590 414612 155040
rect 415912 154590 415972 155040
rect 414430 154530 414612 154590
rect 415534 154530 415972 154590
rect 416048 154590 416108 155040
rect 417000 154590 417060 155040
rect 418088 154730 418148 155040
rect 418088 154670 418170 154730
rect 416048 154530 416146 154590
rect 417000 154530 417066 154590
rect 414430 153101 414490 154530
rect 415534 153101 415594 154530
rect 416086 153237 416146 154530
rect 416083 153236 416149 153237
rect 416083 153172 416084 153236
rect 416148 153172 416149 153236
rect 416083 153171 416149 153172
rect 417006 153101 417066 154530
rect 418110 153101 418170 154670
rect 418496 154590 418556 155040
rect 419448 154590 419508 155040
rect 418478 154530 418556 154590
rect 419214 154530 419508 154590
rect 420672 154590 420732 155040
rect 421080 154590 421140 155040
rect 420672 154530 420746 154590
rect 418478 154461 418538 154530
rect 418475 154460 418541 154461
rect 418475 154396 418476 154460
rect 418540 154396 418541 154460
rect 418475 154395 418541 154396
rect 414427 153100 414493 153101
rect 414427 153036 414428 153100
rect 414492 153036 414493 153100
rect 414427 153035 414493 153036
rect 415531 153100 415597 153101
rect 415531 153036 415532 153100
rect 415596 153036 415597 153100
rect 415531 153035 415597 153036
rect 417003 153100 417069 153101
rect 417003 153036 417004 153100
rect 417068 153036 417069 153100
rect 417003 153035 417069 153036
rect 418107 153100 418173 153101
rect 418107 153036 418108 153100
rect 418172 153036 418173 153100
rect 418107 153035 418173 153036
rect 410747 152556 410813 152557
rect 410747 152492 410748 152556
rect 410812 152492 410813 152556
rect 410747 152491 410813 152492
rect 412403 152556 412469 152557
rect 412403 152492 412404 152556
rect 412468 152492 412469 152556
rect 412403 152491 412469 152492
rect 413691 152556 413757 152557
rect 413691 152492 413692 152556
rect 413756 152492 413757 152556
rect 413691 152491 413757 152492
rect 408954 141318 408986 141554
rect 409222 141318 409306 141554
rect 409542 141318 409574 141554
rect 408954 141234 409574 141318
rect 408954 140998 408986 141234
rect 409222 140998 409306 141234
rect 409542 140998 409574 141234
rect 408954 130308 409574 140998
rect 415794 146514 416414 153000
rect 419214 152557 419274 154530
rect 420686 153101 420746 154530
rect 421054 154530 421140 154590
rect 421760 154590 421820 155040
rect 422848 154590 422908 155040
rect 423528 154590 423588 155040
rect 421760 154530 421850 154590
rect 422848 154530 422954 154590
rect 421054 154461 421114 154530
rect 421051 154460 421117 154461
rect 421051 154396 421052 154460
rect 421116 154396 421117 154460
rect 421051 154395 421117 154396
rect 421790 153101 421850 154530
rect 422894 153101 422954 154530
rect 423446 154530 423588 154590
rect 423936 154590 423996 155040
rect 425296 154590 425356 155040
rect 423936 154530 424058 154590
rect 423446 153917 423506 154530
rect 423443 153916 423509 153917
rect 423443 153852 423444 153916
rect 423508 153852 423509 153916
rect 423443 153851 423509 153852
rect 423998 153101 424058 154530
rect 425286 154530 425356 154590
rect 425976 154590 426036 155040
rect 426384 154730 426444 155040
rect 426384 154670 426450 154730
rect 425976 154530 426082 154590
rect 425286 153101 425346 154530
rect 426022 154461 426082 154530
rect 426019 154460 426085 154461
rect 426019 154396 426020 154460
rect 426084 154396 426085 154460
rect 426019 154395 426085 154396
rect 426390 153101 426450 154670
rect 427608 154590 427668 155040
rect 428288 154590 428348 155040
rect 428696 154590 428756 155040
rect 429784 154590 429844 155040
rect 431008 154590 431068 155040
rect 427608 154530 427738 154590
rect 420683 153100 420749 153101
rect 420683 153036 420684 153100
rect 420748 153036 420749 153100
rect 420683 153035 420749 153036
rect 421787 153100 421853 153101
rect 421787 153036 421788 153100
rect 421852 153036 421853 153100
rect 421787 153035 421853 153036
rect 422891 153100 422957 153101
rect 422891 153036 422892 153100
rect 422956 153036 422957 153100
rect 422891 153035 422957 153036
rect 423995 153100 424061 153101
rect 423995 153036 423996 153100
rect 424060 153036 424061 153100
rect 423995 153035 424061 153036
rect 425283 153100 425349 153101
rect 425283 153036 425284 153100
rect 425348 153036 425349 153100
rect 425283 153035 425349 153036
rect 426387 153100 426453 153101
rect 426387 153036 426388 153100
rect 426452 153036 426453 153100
rect 426387 153035 426453 153036
rect 419211 152556 419277 152557
rect 419211 152492 419212 152556
rect 419276 152492 419277 152556
rect 419211 152491 419277 152492
rect 415794 146278 415826 146514
rect 416062 146278 416146 146514
rect 416382 146278 416414 146514
rect 415794 146194 416414 146278
rect 415794 145958 415826 146194
rect 416062 145958 416146 146194
rect 416382 145958 416414 146194
rect 415794 130308 416414 145958
rect 419514 133174 420134 153000
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 130308 420134 132618
rect 423234 136894 423854 153000
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 130308 423854 136338
rect 426954 140614 427574 153000
rect 427678 152557 427738 154530
rect 427862 154530 428348 154590
rect 428598 154530 428756 154590
rect 429702 154530 429844 154590
rect 430622 154530 431068 154590
rect 431144 154590 431204 155040
rect 432232 154590 432292 155040
rect 431144 154530 431234 154590
rect 427675 152556 427741 152557
rect 427675 152492 427676 152556
rect 427740 152492 427741 152556
rect 427675 152491 427741 152492
rect 427862 151605 427922 154530
rect 428598 153101 428658 154530
rect 429702 153101 429762 154530
rect 428595 153100 428661 153101
rect 428595 153036 428596 153100
rect 428660 153036 428661 153100
rect 428595 153035 428661 153036
rect 429699 153100 429765 153101
rect 429699 153036 429700 153100
rect 429764 153036 429765 153100
rect 429699 153035 429765 153036
rect 430622 151741 430682 154530
rect 431174 153101 431234 154530
rect 431726 154530 432292 154590
rect 433320 154590 433380 155040
rect 433592 154590 433652 155040
rect 433320 154530 433442 154590
rect 431726 153101 431786 154530
rect 431171 153100 431237 153101
rect 431171 153036 431172 153100
rect 431236 153036 431237 153100
rect 431171 153035 431237 153036
rect 431723 153100 431789 153101
rect 431723 153036 431724 153100
rect 431788 153036 431789 153100
rect 431723 153035 431789 153036
rect 433382 152557 433442 154530
rect 433566 154530 433652 154590
rect 434408 154590 434468 155040
rect 435768 154590 435828 155040
rect 436040 154590 436100 155040
rect 436992 154590 437052 155040
rect 434408 154530 434730 154590
rect 435768 154530 435834 154590
rect 433566 153101 433626 154530
rect 434670 153101 434730 154530
rect 433563 153100 433629 153101
rect 433563 153036 433564 153100
rect 433628 153036 433629 153100
rect 433563 153035 433629 153036
rect 434667 153100 434733 153101
rect 434667 153036 434668 153100
rect 434732 153036 434733 153100
rect 434667 153035 434733 153036
rect 433379 152556 433445 152557
rect 433379 152492 433380 152556
rect 433444 152492 433445 152556
rect 433379 152491 433445 152492
rect 430619 151740 430685 151741
rect 430619 151676 430620 151740
rect 430684 151676 430685 151740
rect 430619 151675 430685 151676
rect 427859 151604 427925 151605
rect 427859 151540 427860 151604
rect 427924 151540 427925 151604
rect 427859 151539 427925 151540
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 130308 427574 140058
rect 433794 147454 434414 153000
rect 435774 152557 435834 154530
rect 435958 154530 436100 154590
rect 436878 154530 437052 154590
rect 438080 154590 438140 155040
rect 438488 154590 438548 155040
rect 439168 154590 439228 155040
rect 440936 154590 440996 155040
rect 443520 154730 443580 155040
rect 445968 154730 446028 155040
rect 438080 154530 438410 154590
rect 438488 154530 438594 154590
rect 439168 154530 439330 154590
rect 435958 153101 436018 154530
rect 436878 153101 436938 154530
rect 438350 153101 438410 154530
rect 435955 153100 436021 153101
rect 435955 153036 435956 153100
rect 436020 153036 436021 153100
rect 435955 153035 436021 153036
rect 436875 153100 436941 153101
rect 436875 153036 436876 153100
rect 436940 153036 436941 153100
rect 436875 153035 436941 153036
rect 438347 153100 438413 153101
rect 438347 153036 438348 153100
rect 438412 153036 438413 153100
rect 438347 153035 438413 153036
rect 435771 152556 435837 152557
rect 435771 152492 435772 152556
rect 435836 152492 435837 152556
rect 435771 152491 435837 152492
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 130308 434414 146898
rect 437514 151174 438134 153000
rect 438534 152557 438594 154530
rect 439270 153101 439330 154530
rect 440926 154530 440996 154590
rect 443502 154670 443580 154730
rect 445894 154670 446028 154730
rect 448280 154730 448340 155040
rect 451000 154730 451060 155040
rect 448280 154670 448346 154730
rect 451000 154670 451106 154730
rect 440926 153101 440986 154530
rect 443502 154461 443562 154670
rect 443499 154460 443565 154461
rect 443499 154396 443500 154460
rect 443564 154396 443565 154460
rect 443499 154395 443565 154396
rect 445894 153101 445954 154670
rect 448286 153101 448346 154670
rect 451046 153101 451106 154670
rect 453448 154590 453508 155040
rect 455896 154590 455956 155040
rect 458480 154590 458540 155040
rect 453438 154530 453508 154590
rect 455830 154530 455956 154590
rect 458406 154530 458540 154590
rect 460928 154590 460988 155040
rect 463512 154590 463572 155040
rect 465960 154590 466020 155040
rect 468544 154590 468604 155040
rect 470992 154730 471052 155040
rect 460928 154530 461042 154590
rect 463512 154530 463618 154590
rect 453438 153101 453498 154530
rect 455830 153237 455890 154530
rect 455827 153236 455893 153237
rect 455827 153172 455828 153236
rect 455892 153172 455893 153236
rect 455827 153171 455893 153172
rect 458406 153101 458466 154530
rect 439267 153100 439333 153101
rect 439267 153036 439268 153100
rect 439332 153036 439333 153100
rect 439267 153035 439333 153036
rect 440923 153100 440989 153101
rect 440923 153036 440924 153100
rect 440988 153036 440989 153100
rect 440923 153035 440989 153036
rect 445891 153100 445957 153101
rect 445891 153036 445892 153100
rect 445956 153036 445957 153100
rect 445891 153035 445957 153036
rect 448283 153100 448349 153101
rect 448283 153036 448284 153100
rect 448348 153036 448349 153100
rect 448283 153035 448349 153036
rect 451043 153100 451109 153101
rect 451043 153036 451044 153100
rect 451108 153036 451109 153100
rect 451043 153035 451109 153036
rect 453435 153100 453501 153101
rect 453435 153036 453436 153100
rect 453500 153036 453501 153100
rect 453435 153035 453501 153036
rect 458403 153100 458469 153101
rect 458403 153036 458404 153100
rect 458468 153036 458469 153100
rect 458403 153035 458469 153036
rect 438531 152556 438597 152557
rect 438531 152492 438532 152556
rect 438596 152492 438597 152556
rect 438531 152491 438597 152492
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 130308 438134 150618
rect 441234 137834 441854 153000
rect 441234 137598 441266 137834
rect 441502 137598 441586 137834
rect 441822 137598 441854 137834
rect 441234 137514 441854 137598
rect 441234 137278 441266 137514
rect 441502 137278 441586 137514
rect 441822 137278 441854 137514
rect 441234 130308 441854 137278
rect 444954 141554 445574 153000
rect 444954 141318 444986 141554
rect 445222 141318 445306 141554
rect 445542 141318 445574 141554
rect 444954 141234 445574 141318
rect 444954 140998 444986 141234
rect 445222 140998 445306 141234
rect 445542 140998 445574 141234
rect 444954 130308 445574 140998
rect 451794 146514 452414 153000
rect 451794 146278 451826 146514
rect 452062 146278 452146 146514
rect 452382 146278 452414 146514
rect 451794 146194 452414 146278
rect 451794 145958 451826 146194
rect 452062 145958 452146 146194
rect 452382 145958 452414 146194
rect 451794 130308 452414 145958
rect 455514 133174 456134 153000
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 130308 456134 132618
rect 459234 136894 459854 153000
rect 460982 152693 461042 154530
rect 463558 153237 463618 154530
rect 465950 154530 466020 154590
rect 468526 154530 468604 154590
rect 470918 154670 471052 154730
rect 473440 154730 473500 155040
rect 475888 154730 475948 155040
rect 478472 154730 478532 155040
rect 480920 154730 480980 155040
rect 483368 154730 483428 155040
rect 473440 154670 473554 154730
rect 463555 153236 463621 153237
rect 463555 153172 463556 153236
rect 463620 153172 463621 153236
rect 463555 153171 463621 153172
rect 460979 152692 461045 152693
rect 460979 152628 460980 152692
rect 461044 152628 461045 152692
rect 460979 152627 461045 152628
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 130308 459854 136338
rect 462954 140614 463574 153000
rect 465950 152285 466010 154530
rect 468526 152829 468586 154530
rect 470918 154053 470978 154670
rect 473494 154189 473554 154670
rect 475886 154670 475948 154730
rect 478462 154670 478532 154730
rect 480854 154670 480980 154730
rect 483246 154670 483428 154730
rect 485952 154730 486012 155040
rect 503224 154730 503284 155040
rect 485952 154670 486066 154730
rect 475886 154325 475946 154670
rect 478462 154325 478522 154670
rect 475883 154324 475949 154325
rect 475883 154260 475884 154324
rect 475948 154260 475949 154324
rect 475883 154259 475949 154260
rect 478459 154324 478525 154325
rect 478459 154260 478460 154324
rect 478524 154260 478525 154324
rect 478459 154259 478525 154260
rect 480854 154189 480914 154670
rect 473491 154188 473557 154189
rect 473491 154124 473492 154188
rect 473556 154124 473557 154188
rect 473491 154123 473557 154124
rect 480851 154188 480917 154189
rect 480851 154124 480852 154188
rect 480916 154124 480917 154188
rect 480851 154123 480917 154124
rect 483246 154053 483306 154670
rect 470915 154052 470981 154053
rect 470915 153988 470916 154052
rect 470980 153988 470981 154052
rect 470915 153987 470981 153988
rect 483243 154052 483309 154053
rect 483243 153988 483244 154052
rect 483308 153988 483309 154052
rect 483243 153987 483309 153988
rect 486006 153917 486066 154670
rect 503118 154670 503284 154730
rect 503360 154730 503420 155040
rect 503360 154670 503546 154730
rect 486003 153916 486069 153917
rect 486003 153852 486004 153916
rect 486068 153852 486069 153916
rect 486003 153851 486069 153852
rect 468523 152828 468589 152829
rect 468523 152764 468524 152828
rect 468588 152764 468589 152828
rect 468523 152763 468589 152764
rect 465947 152284 466013 152285
rect 465947 152220 465948 152284
rect 466012 152220 466013 152284
rect 465947 152219 466013 152220
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 130308 463574 140058
rect 469794 147454 470414 153000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 130308 470414 146898
rect 473514 151174 474134 153000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 130308 474134 150618
rect 477234 137834 477854 153000
rect 477234 137598 477266 137834
rect 477502 137598 477586 137834
rect 477822 137598 477854 137834
rect 477234 137514 477854 137598
rect 477234 137278 477266 137514
rect 477502 137278 477586 137514
rect 477822 137278 477854 137514
rect 477234 130308 477854 137278
rect 480954 141554 481574 153000
rect 480954 141318 480986 141554
rect 481222 141318 481306 141554
rect 481542 141318 481574 141554
rect 480954 141234 481574 141318
rect 480954 140998 480986 141234
rect 481222 140998 481306 141234
rect 481542 140998 481574 141234
rect 480954 130308 481574 140998
rect 487794 146514 488414 153000
rect 487794 146278 487826 146514
rect 488062 146278 488146 146514
rect 488382 146278 488414 146514
rect 487794 146194 488414 146278
rect 487794 145958 487826 146194
rect 488062 145958 488146 146194
rect 488382 145958 488414 146194
rect 487794 130308 488414 145958
rect 491514 133174 492134 153000
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 130308 492134 132618
rect 495234 136894 495854 153000
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 130308 495854 136338
rect 498954 140614 499574 153000
rect 503118 152557 503178 154670
rect 503486 152693 503546 154670
rect 503483 152692 503549 152693
rect 503483 152628 503484 152692
rect 503548 152628 503549 152692
rect 503483 152627 503549 152628
rect 503115 152556 503181 152557
rect 503115 152492 503116 152556
rect 503180 152492 503181 152556
rect 503115 152491 503181 152492
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 130308 499574 140058
rect 505794 147454 506414 153000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 130308 506414 146898
rect 509514 151174 510134 153000
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 130308 510134 150618
rect 513234 137834 513854 153000
rect 513234 137598 513266 137834
rect 513502 137598 513586 137834
rect 513822 137598 513854 137834
rect 513234 137514 513854 137598
rect 513234 137278 513266 137514
rect 513502 137278 513586 137514
rect 513822 137278 513854 137514
rect 510843 130388 510909 130389
rect 510843 130324 510844 130388
rect 510908 130324 510909 130388
rect 510843 130323 510909 130324
rect 498515 129844 498581 129845
rect 498515 129780 498516 129844
rect 498580 129780 498581 129844
rect 498515 129779 498581 129780
rect 499803 129844 499869 129845
rect 499803 129780 499804 129844
rect 499868 129780 499869 129844
rect 499803 129779 499869 129780
rect 498518 128890 498578 129779
rect 499806 128890 499866 129779
rect 510846 128890 510906 130323
rect 513234 130308 513854 137278
rect 516954 141554 517574 153000
rect 516954 141318 516986 141554
rect 517222 141318 517306 141554
rect 517542 141318 517574 141554
rect 516954 141234 517574 141318
rect 516954 140998 516986 141234
rect 517222 140998 517306 141234
rect 517542 140998 517574 141234
rect 516954 130308 517574 140998
rect 498464 128830 498578 128890
rect 499688 128830 499866 128890
rect 510840 128830 510906 128890
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 498464 128202 498524 128830
rect 499688 128202 499748 128830
rect 510840 128202 510900 128830
rect 380952 111454 381300 111486
rect 380952 111218 381008 111454
rect 381244 111218 381300 111454
rect 380952 111134 381300 111218
rect 380952 110898 381008 111134
rect 381244 110898 381300 111134
rect 380952 110866 381300 110898
rect 515320 111454 515668 111486
rect 515320 111218 515376 111454
rect 515612 111218 515668 111454
rect 515320 111134 515668 111218
rect 515320 110898 515376 111134
rect 515612 110898 515668 111134
rect 515320 110866 515668 110898
rect 380272 93454 380620 93486
rect 380272 93218 380328 93454
rect 380564 93218 380620 93454
rect 380272 93134 380620 93218
rect 380272 92898 380328 93134
rect 380564 92898 380620 93134
rect 380272 92866 380620 92898
rect 516000 93454 516348 93486
rect 516000 93218 516056 93454
rect 516292 93218 516348 93454
rect 516000 93134 516348 93218
rect 516000 92898 516056 93134
rect 516292 92898 516348 93134
rect 516000 92866 516348 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 380952 75454 381300 75486
rect 380952 75218 381008 75454
rect 381244 75218 381300 75454
rect 380952 75134 381300 75218
rect 380952 74898 381008 75134
rect 381244 74898 381300 75134
rect 380952 74866 381300 74898
rect 515320 75454 515668 75486
rect 515320 75218 515376 75454
rect 515612 75218 515668 75454
rect 515320 75134 515668 75218
rect 515320 74898 515376 75134
rect 515612 74898 515668 75134
rect 515320 74866 515668 74898
rect 380272 57454 380620 57486
rect 380272 57218 380328 57454
rect 380564 57218 380620 57454
rect 380272 57134 380620 57218
rect 380272 56898 380328 57134
rect 380564 56898 380620 57134
rect 380272 56866 380620 56898
rect 516000 57454 516348 57486
rect 516000 57218 516056 57454
rect 516292 57218 516348 57454
rect 516000 57134 516348 57218
rect 516000 56898 516056 57134
rect 516292 56898 516348 57134
rect 516000 56866 516348 56898
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 379470 45510 379714 45570
rect 378915 41580 378981 41581
rect 378915 41516 378916 41580
rect 378980 41516 378981 41580
rect 378915 41515 378981 41516
rect 377811 41172 377877 41173
rect 377811 41108 377812 41172
rect 377876 41108 377877 41172
rect 377811 41107 377877 41108
rect 377259 41036 377325 41037
rect 377259 40972 377260 41036
rect 377324 40972 377325 41036
rect 377259 40971 377325 40972
rect 379470 40901 379530 45510
rect 396056 44845 396116 45106
rect 397144 44845 397204 45106
rect 396053 44844 396119 44845
rect 396053 44780 396054 44844
rect 396118 44780 396119 44844
rect 396053 44779 396119 44780
rect 397141 44844 397207 44845
rect 397141 44780 397142 44844
rect 397206 44780 397207 44844
rect 397141 44779 397207 44780
rect 398232 44570 398292 45106
rect 399592 44842 399652 45106
rect 400544 44842 400604 45106
rect 399526 44782 399652 44842
rect 400446 44782 400604 44842
rect 398232 44510 398298 44570
rect 398238 43213 398298 44510
rect 398235 43212 398301 43213
rect 398235 43148 398236 43212
rect 398300 43148 398301 43212
rect 398235 43147 398301 43148
rect 379467 40900 379533 40901
rect 379467 40836 379468 40900
rect 379532 40836 379533 40900
rect 379467 40835 379533 40836
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 43000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 43000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 43000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 43000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 43000
rect 399526 42805 399586 44782
rect 399523 42804 399589 42805
rect 399523 42740 399524 42804
rect 399588 42740 399589 42804
rect 399523 42739 399589 42740
rect 400446 41853 400506 44782
rect 401768 44570 401828 45106
rect 403128 44845 403188 45106
rect 403125 44844 403191 44845
rect 403125 44780 403126 44844
rect 403190 44780 403191 44844
rect 403125 44779 403191 44780
rect 404216 44573 404276 45106
rect 405440 44573 405500 45106
rect 406528 44573 406588 45106
rect 401734 44510 401828 44570
rect 404213 44572 404279 44573
rect 401734 43213 401794 44510
rect 404213 44508 404214 44572
rect 404278 44508 404279 44572
rect 404213 44507 404279 44508
rect 405437 44572 405503 44573
rect 405437 44508 405438 44572
rect 405502 44508 405503 44572
rect 405437 44507 405503 44508
rect 406525 44572 406591 44573
rect 406525 44508 406526 44572
rect 406590 44508 406591 44572
rect 407616 44570 407676 45106
rect 408296 44570 408356 45106
rect 408704 44570 408764 45106
rect 410064 44570 410124 45106
rect 410744 44709 410804 45106
rect 410741 44708 410807 44709
rect 410741 44644 410742 44708
rect 410806 44644 410807 44708
rect 410741 44643 410807 44644
rect 407616 44510 407682 44570
rect 408296 44510 408418 44570
rect 408704 44510 408786 44570
rect 406525 44507 406591 44508
rect 407622 43485 407682 44510
rect 407619 43484 407685 43485
rect 407619 43420 407620 43484
rect 407684 43420 407685 43484
rect 407619 43419 407685 43420
rect 401731 43212 401797 43213
rect 401731 43148 401732 43212
rect 401796 43148 401797 43212
rect 401731 43147 401797 43148
rect 400443 41852 400509 41853
rect 400443 41788 400444 41852
rect 400508 41788 400509 41852
rect 400443 41787 400509 41788
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 43000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 43000
rect 408358 42805 408418 44510
rect 408726 42805 408786 44510
rect 410014 44510 410124 44570
rect 411288 44570 411348 45106
rect 412376 44570 412436 45106
rect 413464 44570 413524 45106
rect 411288 44510 411362 44570
rect 412376 44510 412466 44570
rect 408355 42804 408421 42805
rect 408355 42740 408356 42804
rect 408420 42740 408421 42804
rect 408355 42739 408421 42740
rect 408723 42804 408789 42805
rect 408723 42740 408724 42804
rect 408788 42740 408789 42804
rect 408723 42739 408789 42740
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 43000
rect 410014 42805 410074 44510
rect 411302 42805 411362 44510
rect 412406 42805 412466 44510
rect 413326 44510 413524 44570
rect 413600 44570 413660 45106
rect 414552 44845 414612 45106
rect 414549 44844 414615 44845
rect 414549 44780 414550 44844
rect 414614 44780 414615 44844
rect 414549 44779 414615 44780
rect 415912 44570 415972 45106
rect 413600 44510 413754 44570
rect 413326 42805 413386 44510
rect 413694 42805 413754 44510
rect 415534 44510 415972 44570
rect 416048 44570 416108 45106
rect 417000 44845 417060 45106
rect 416997 44844 417063 44845
rect 416997 44780 416998 44844
rect 417062 44780 417063 44844
rect 416997 44779 417063 44780
rect 418088 44573 418148 45106
rect 418088 44572 418173 44573
rect 416048 44510 416698 44570
rect 418088 44510 418108 44572
rect 415534 42805 415594 44510
rect 410011 42804 410077 42805
rect 410011 42740 410012 42804
rect 410076 42740 410077 42804
rect 410011 42739 410077 42740
rect 411299 42804 411365 42805
rect 411299 42740 411300 42804
rect 411364 42740 411365 42804
rect 411299 42739 411365 42740
rect 412403 42804 412469 42805
rect 412403 42740 412404 42804
rect 412468 42740 412469 42804
rect 412403 42739 412469 42740
rect 413323 42804 413389 42805
rect 413323 42740 413324 42804
rect 413388 42740 413389 42804
rect 413323 42739 413389 42740
rect 413691 42804 413757 42805
rect 413691 42740 413692 42804
rect 413756 42740 413757 42804
rect 413691 42739 413757 42740
rect 415531 42804 415597 42805
rect 415531 42740 415532 42804
rect 415596 42740 415597 42804
rect 415531 42739 415597 42740
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 43000
rect 416638 41989 416698 44510
rect 418107 44508 418108 44510
rect 418172 44508 418173 44572
rect 418496 44570 418556 45106
rect 419448 44709 419508 45106
rect 419445 44708 419511 44709
rect 419445 44644 419446 44708
rect 419510 44644 419511 44708
rect 419445 44643 419511 44644
rect 420672 44573 420732 45106
rect 418107 44507 418173 44508
rect 418478 44510 418556 44570
rect 420669 44572 420735 44573
rect 416635 41988 416701 41989
rect 416635 41924 416636 41988
rect 416700 41924 416701 41988
rect 416635 41923 416701 41924
rect 418478 41445 418538 44510
rect 420669 44508 420670 44572
rect 420734 44508 420735 44572
rect 421080 44570 421140 45106
rect 421760 44573 421820 45106
rect 422848 44573 422908 45106
rect 423528 44573 423588 45106
rect 423936 44709 423996 45106
rect 423933 44708 423999 44709
rect 423933 44644 423934 44708
rect 423998 44644 423999 44708
rect 423933 44643 423999 44644
rect 420669 44507 420735 44508
rect 421054 44510 421140 44570
rect 421757 44572 421823 44573
rect 421054 43485 421114 44510
rect 421757 44508 421758 44572
rect 421822 44508 421823 44572
rect 421757 44507 421823 44508
rect 422845 44572 422911 44573
rect 422845 44508 422846 44572
rect 422910 44508 422911 44572
rect 422845 44507 422911 44508
rect 423525 44572 423591 44573
rect 423525 44508 423526 44572
rect 423590 44508 423591 44572
rect 425296 44570 425356 45106
rect 425976 44573 426036 45106
rect 423525 44507 423591 44508
rect 425286 44510 425356 44570
rect 425973 44572 426039 44573
rect 425286 44437 425346 44510
rect 425973 44508 425974 44572
rect 426038 44508 426039 44572
rect 426384 44570 426444 45106
rect 427608 44570 427668 45106
rect 428288 44570 428348 45106
rect 428696 44570 428756 45106
rect 429784 44570 429844 45106
rect 431008 44570 431068 45106
rect 426384 44510 426450 44570
rect 427608 44510 427738 44570
rect 425973 44507 426039 44508
rect 425283 44436 425349 44437
rect 425283 44372 425284 44436
rect 425348 44372 425349 44436
rect 425283 44371 425349 44372
rect 421051 43484 421117 43485
rect 421051 43420 421052 43484
rect 421116 43420 421117 43484
rect 421051 43419 421117 43420
rect 418475 41444 418541 41445
rect 418475 41380 418476 41444
rect 418540 41380 418541 41444
rect 418475 41379 418541 41380
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 43000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 43000
rect 426390 42805 426450 44510
rect 426387 42804 426453 42805
rect 426387 42740 426388 42804
rect 426452 42740 426453 42804
rect 426387 42739 426453 42740
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 43000
rect 427678 42805 427738 44510
rect 428230 44510 428348 44570
rect 428598 44510 428756 44570
rect 429702 44510 429844 44570
rect 430990 44510 431068 44570
rect 431144 44570 431204 45106
rect 432232 44570 432292 45106
rect 433320 44570 433380 45106
rect 433592 44570 433652 45106
rect 431144 44510 431234 44570
rect 432232 44510 432338 44570
rect 433320 44510 433442 44570
rect 428230 43485 428290 44510
rect 428227 43484 428293 43485
rect 428227 43420 428228 43484
rect 428292 43420 428293 43484
rect 428227 43419 428293 43420
rect 428598 42805 428658 44510
rect 429702 42805 429762 44510
rect 430990 42805 431050 44510
rect 427675 42804 427741 42805
rect 427675 42740 427676 42804
rect 427740 42740 427741 42804
rect 427675 42739 427741 42740
rect 428595 42804 428661 42805
rect 428595 42740 428596 42804
rect 428660 42740 428661 42804
rect 428595 42739 428661 42740
rect 429699 42804 429765 42805
rect 429699 42740 429700 42804
rect 429764 42740 429765 42804
rect 429699 42739 429765 42740
rect 430987 42804 431053 42805
rect 430987 42740 430988 42804
rect 431052 42740 431053 42804
rect 430987 42739 431053 42740
rect 431174 41989 431234 44510
rect 432278 42805 432338 44510
rect 433382 42805 433442 44510
rect 433566 44510 433652 44570
rect 434408 44570 434468 45106
rect 435768 44570 435828 45106
rect 436040 44570 436100 45106
rect 436992 44570 437052 45106
rect 434408 44510 434730 44570
rect 435768 44510 435834 44570
rect 432275 42804 432341 42805
rect 432275 42740 432276 42804
rect 432340 42740 432341 42804
rect 432275 42739 432341 42740
rect 433379 42804 433445 42805
rect 433379 42740 433380 42804
rect 433444 42740 433445 42804
rect 433379 42739 433445 42740
rect 433566 42125 433626 44510
rect 433563 42124 433629 42125
rect 433563 42060 433564 42124
rect 433628 42060 433629 42124
rect 433563 42059 433629 42060
rect 431171 41988 431237 41989
rect 431171 41924 431172 41988
rect 431236 41924 431237 41988
rect 431171 41923 431237 41924
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 43000
rect 434670 42805 434730 44510
rect 434667 42804 434733 42805
rect 434667 42740 434668 42804
rect 434732 42740 434733 42804
rect 434667 42739 434733 42740
rect 435774 42125 435834 44510
rect 435958 44510 436100 44570
rect 436878 44510 437052 44570
rect 438080 44570 438140 45106
rect 438488 44570 438548 45106
rect 439168 44573 439228 45106
rect 439165 44572 439231 44573
rect 438080 44510 438410 44570
rect 438488 44510 438594 44570
rect 435958 42805 436018 44510
rect 436878 42805 436938 44510
rect 435955 42804 436021 42805
rect 435955 42740 435956 42804
rect 436020 42740 436021 42804
rect 435955 42739 436021 42740
rect 436875 42804 436941 42805
rect 436875 42740 436876 42804
rect 436940 42740 436941 42804
rect 436875 42739 436941 42740
rect 435771 42124 435837 42125
rect 435771 42060 435772 42124
rect 435836 42060 435837 42124
rect 435771 42059 435837 42060
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 43000
rect 438350 41445 438410 44510
rect 438534 42805 438594 44510
rect 439165 44508 439166 44572
rect 439230 44508 439231 44572
rect 440936 44570 440996 45106
rect 443520 44570 443580 45106
rect 445968 44570 446028 45106
rect 439165 44507 439231 44508
rect 440926 44510 440996 44570
rect 443502 44510 443580 44570
rect 445894 44510 446028 44570
rect 448280 44570 448340 45106
rect 451000 44570 451060 45106
rect 453448 44570 453508 45106
rect 455896 44573 455956 45106
rect 458480 44573 458540 45106
rect 448280 44510 448346 44570
rect 451000 44510 451106 44570
rect 440926 42805 440986 44510
rect 438531 42804 438597 42805
rect 438531 42740 438532 42804
rect 438596 42740 438597 42804
rect 438531 42739 438597 42740
rect 440923 42804 440989 42805
rect 440923 42740 440924 42804
rect 440988 42740 440989 42804
rect 440923 42739 440989 42740
rect 438347 41444 438413 41445
rect 438347 41380 438348 41444
rect 438412 41380 438413 41444
rect 438347 41379 438413 41380
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 43000
rect 443502 42805 443562 44510
rect 443499 42804 443565 42805
rect 443499 42740 443500 42804
rect 443564 42740 443565 42804
rect 443499 42739 443565 42740
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 43000
rect 445894 42805 445954 44510
rect 448286 42805 448346 44510
rect 445891 42804 445957 42805
rect 445891 42740 445892 42804
rect 445956 42740 445957 42804
rect 445891 42739 445957 42740
rect 448283 42804 448349 42805
rect 448283 42740 448284 42804
rect 448348 42740 448349 42804
rect 448283 42739 448349 42740
rect 451046 42261 451106 44510
rect 453438 44510 453508 44570
rect 455893 44572 455959 44573
rect 451043 42260 451109 42261
rect 451043 42196 451044 42260
rect 451108 42196 451109 42260
rect 451043 42195 451109 42196
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 43000
rect 453438 42805 453498 44510
rect 455893 44508 455894 44572
rect 455958 44508 455959 44572
rect 455893 44507 455959 44508
rect 458477 44572 458543 44573
rect 458477 44508 458478 44572
rect 458542 44508 458543 44572
rect 460928 44570 460988 45106
rect 463512 44570 463572 45106
rect 465960 44570 466020 45106
rect 468544 44570 468604 45106
rect 470992 44570 471052 45106
rect 460928 44510 461042 44570
rect 463512 44510 463618 44570
rect 458477 44507 458543 44508
rect 453435 42804 453501 42805
rect 453435 42740 453436 42804
rect 453500 42740 453501 42804
rect 453435 42739 453501 42740
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 43000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 43000
rect 460982 42397 461042 44510
rect 463558 43485 463618 44510
rect 465950 44510 466020 44570
rect 468526 44510 468604 44570
rect 470918 44510 471052 44570
rect 473440 44570 473500 45106
rect 475888 44570 475948 45106
rect 478472 44570 478532 45106
rect 480920 44573 480980 45106
rect 473440 44510 473554 44570
rect 463555 43484 463621 43485
rect 463555 43420 463556 43484
rect 463620 43420 463621 43484
rect 463555 43419 463621 43420
rect 460979 42396 461045 42397
rect 460979 42332 460980 42396
rect 461044 42332 461045 42396
rect 460979 42331 461045 42332
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 43000
rect 465950 42669 466010 44510
rect 468526 43893 468586 44510
rect 468523 43892 468589 43893
rect 468523 43828 468524 43892
rect 468588 43828 468589 43892
rect 468523 43827 468589 43828
rect 465947 42668 466013 42669
rect 465947 42604 465948 42668
rect 466012 42604 466013 42668
rect 465947 42603 466013 42604
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 43000
rect 470918 42533 470978 44510
rect 473494 43757 473554 44510
rect 475886 44510 475948 44570
rect 478462 44510 478532 44570
rect 480917 44572 480983 44573
rect 473491 43756 473557 43757
rect 473491 43692 473492 43756
rect 473556 43692 473557 43756
rect 473491 43691 473557 43692
rect 470915 42532 470981 42533
rect 470915 42468 470916 42532
rect 470980 42468 470981 42532
rect 470915 42467 470981 42468
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 43000
rect 475886 41581 475946 44510
rect 478462 44029 478522 44510
rect 480917 44508 480918 44572
rect 480982 44508 480983 44572
rect 483368 44570 483428 45106
rect 485952 44570 486012 45106
rect 503224 44570 503284 45106
rect 483368 44510 483490 44570
rect 485952 44510 486066 44570
rect 480917 44507 480983 44508
rect 483430 44165 483490 44510
rect 483427 44164 483493 44165
rect 483427 44100 483428 44164
rect 483492 44100 483493 44164
rect 483427 44099 483493 44100
rect 478459 44028 478525 44029
rect 478459 43964 478460 44028
rect 478524 43964 478525 44028
rect 478459 43963 478525 43964
rect 475883 41580 475949 41581
rect 475883 41516 475884 41580
rect 475948 41516 475949 41580
rect 475883 41515 475949 41516
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 43000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 43000
rect 486006 42805 486066 44510
rect 503118 44510 503284 44570
rect 503360 44570 503420 45106
rect 503360 44510 503546 44570
rect 486003 42804 486069 42805
rect 486003 42740 486004 42804
rect 486068 42740 486069 42804
rect 486003 42739 486069 42740
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 43000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 43000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 43000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 43000
rect 503118 42805 503178 44510
rect 503486 42805 503546 44510
rect 503115 42804 503181 42805
rect 503115 42740 503116 42804
rect 503180 42740 503181 42804
rect 503115 42739 503181 42740
rect 503483 42804 503549 42805
rect 503483 42740 503484 42804
rect 503548 42740 503549 42804
rect 503483 42739 503549 42740
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 43000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 43000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 43000
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 43000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 79610 633218 79846 633454
rect 79610 632898 79846 633134
rect 110330 633218 110566 633454
rect 110330 632898 110566 633134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 79610 597218 79846 597454
rect 79610 596898 79846 597134
rect 110330 597218 110566 597454
rect 110330 596898 110566 597134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 64250 579218 64486 579454
rect 64250 578898 64486 579134
rect 94970 579218 95206 579454
rect 94970 578898 95206 579134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 73826 562158 74062 562394
rect 74146 562158 74382 562394
rect 73826 561838 74062 562074
rect 74146 561838 74382 562074
rect 77546 565878 77782 566114
rect 77866 565878 78102 566114
rect 77546 565558 77782 565794
rect 77866 565558 78102 565794
rect 81266 567718 81502 567954
rect 81586 567718 81822 567954
rect 81266 567398 81502 567634
rect 81586 567398 81822 567634
rect 84986 571438 85222 571674
rect 85306 571438 85542 571674
rect 84986 571118 85222 571354
rect 85306 571118 85542 571354
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 562158 110062 562394
rect 110146 562158 110382 562394
rect 109826 561838 110062 562074
rect 110146 561838 110382 562074
rect 113546 565878 113782 566114
rect 113866 565878 114102 566114
rect 113546 565558 113782 565794
rect 113866 565558 114102 565794
rect 117266 567718 117502 567954
rect 117586 567718 117822 567954
rect 117266 567398 117502 567634
rect 117586 567398 117822 567634
rect 120986 571438 121222 571674
rect 121306 571438 121542 571674
rect 120986 571118 121222 571354
rect 121306 571118 121542 571354
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 159610 633218 159846 633454
rect 159610 632898 159846 633134
rect 190330 633218 190566 633454
rect 190330 632898 190566 633134
rect 144250 615218 144486 615454
rect 144250 614898 144486 615134
rect 174970 615218 175206 615454
rect 174970 614898 175206 615134
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 159610 597218 159846 597454
rect 159610 596898 159846 597134
rect 190330 597218 190566 597454
rect 190330 596898 190566 597134
rect 144250 579218 144486 579454
rect 144250 578898 144486 579134
rect 174970 579218 175206 579454
rect 174970 578898 175206 579134
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 562158 146062 562394
rect 146146 562158 146382 562394
rect 145826 561838 146062 562074
rect 146146 561838 146382 562074
rect 149546 565878 149782 566114
rect 149866 565878 150102 566114
rect 149546 565558 149782 565794
rect 149866 565558 150102 565794
rect 153266 567718 153502 567954
rect 153586 567718 153822 567954
rect 153266 567398 153502 567634
rect 153586 567398 153822 567634
rect 156986 571438 157222 571674
rect 157306 571438 157542 571674
rect 156986 571118 157222 571354
rect 157306 571118 157542 571354
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 562158 182062 562394
rect 182146 562158 182382 562394
rect 181826 561838 182062 562074
rect 182146 561838 182382 562074
rect 185546 565878 185782 566114
rect 185866 565878 186102 566114
rect 185546 565558 185782 565794
rect 185866 565558 186102 565794
rect 189266 567718 189502 567954
rect 189586 567718 189822 567954
rect 189266 567398 189502 567634
rect 189586 567398 189822 567634
rect 192986 571438 193222 571674
rect 193306 571438 193542 571674
rect 192986 571118 193222 571354
rect 193306 571118 193542 571354
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 239610 633218 239846 633454
rect 239610 632898 239846 633134
rect 270330 633218 270566 633454
rect 270330 632898 270566 633134
rect 224250 615218 224486 615454
rect 224250 614898 224486 615134
rect 254970 615218 255206 615454
rect 254970 614898 255206 615134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 239610 597218 239846 597454
rect 239610 596898 239846 597134
rect 270330 597218 270566 597454
rect 270330 596898 270566 597134
rect 224250 579218 224486 579454
rect 224250 578898 224486 579134
rect 254970 579218 255206 579454
rect 254970 578898 255206 579134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 562158 218062 562394
rect 218146 562158 218382 562394
rect 217826 561838 218062 562074
rect 218146 561838 218382 562074
rect 221546 565878 221782 566114
rect 221866 565878 222102 566114
rect 221546 565558 221782 565794
rect 221866 565558 222102 565794
rect 225266 567718 225502 567954
rect 225586 567718 225822 567954
rect 225266 567398 225502 567634
rect 225586 567398 225822 567634
rect 228986 571438 229222 571674
rect 229306 571438 229542 571674
rect 228986 571118 229222 571354
rect 229306 571118 229542 571354
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 562158 254062 562394
rect 254146 562158 254382 562394
rect 253826 561838 254062 562074
rect 254146 561838 254382 562074
rect 257546 565878 257782 566114
rect 257866 565878 258102 566114
rect 257546 565558 257782 565794
rect 257866 565558 258102 565794
rect 261266 567718 261502 567954
rect 261586 567718 261822 567954
rect 261266 567398 261502 567634
rect 261586 567398 261822 567634
rect 264986 571438 265222 571674
rect 265306 571438 265542 571674
rect 264986 571118 265222 571354
rect 265306 571118 265542 571354
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 64250 543218 64486 543454
rect 64250 542898 64486 543134
rect 94970 543218 95206 543454
rect 94970 542898 95206 543134
rect 125690 543218 125926 543454
rect 125690 542898 125926 543134
rect 156410 543218 156646 543454
rect 156410 542898 156646 543134
rect 187130 543218 187366 543454
rect 187130 542898 187366 543134
rect 217850 543218 218086 543454
rect 217850 542898 218086 543134
rect 248570 543218 248806 543454
rect 248570 542898 248806 543134
rect 279290 543218 279526 543454
rect 279290 542898 279526 543134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 79610 525218 79846 525454
rect 79610 524898 79846 525134
rect 110330 525218 110566 525454
rect 110330 524898 110566 525134
rect 141050 525218 141286 525454
rect 141050 524898 141286 525134
rect 171770 525218 172006 525454
rect 171770 524898 172006 525134
rect 202490 525218 202726 525454
rect 202490 524898 202726 525134
rect 233210 525218 233446 525454
rect 233210 524898 233446 525134
rect 263930 525218 264166 525454
rect 263930 524898 264166 525134
rect 294650 525218 294886 525454
rect 294650 524898 294886 525134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 475878 59782 476114
rect 59866 475878 60102 476114
rect 59546 475558 59782 475794
rect 59866 475558 60102 475794
rect 63266 477718 63502 477954
rect 63586 477718 63822 477954
rect 63266 477398 63502 477634
rect 63586 477398 63822 477634
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 475878 95782 476114
rect 95866 475878 96102 476114
rect 95546 475558 95782 475794
rect 95866 475558 96102 475794
rect 99266 477718 99502 477954
rect 99586 477718 99822 477954
rect 99266 477398 99502 477634
rect 99586 477398 99822 477634
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 475878 131782 476114
rect 131866 475878 132102 476114
rect 131546 475558 131782 475794
rect 131866 475558 132102 475794
rect 135266 477718 135502 477954
rect 135586 477718 135822 477954
rect 135266 477398 135502 477634
rect 135586 477398 135822 477634
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 475878 167782 476114
rect 167866 475878 168102 476114
rect 167546 475558 167782 475794
rect 167866 475558 168102 475794
rect 171266 477718 171502 477954
rect 171586 477718 171822 477954
rect 171266 477398 171502 477634
rect 171586 477398 171822 477634
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 61008 399218 61244 399454
rect 61008 398898 61244 399134
rect 195376 399218 195612 399454
rect 195376 398898 195612 399134
rect 60328 381218 60564 381454
rect 60328 380898 60564 381134
rect 196056 381218 196292 381454
rect 196056 380898 196292 381134
rect 59546 365998 59782 366234
rect 59866 365998 60102 366234
rect 59546 365678 59782 365914
rect 59866 365678 60102 365914
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 84986 357318 85222 357554
rect 85306 357318 85542 357554
rect 84986 356998 85222 357234
rect 85306 356998 85542 357234
rect 91826 362278 92062 362514
rect 92146 362278 92382 362514
rect 91826 361958 92062 362194
rect 92146 361958 92382 362194
rect 95546 365998 95782 366234
rect 95866 365998 96102 366234
rect 95546 365678 95782 365914
rect 95866 365678 96102 365914
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 357318 121222 357554
rect 121306 357318 121542 357554
rect 120986 356998 121222 357234
rect 121306 356998 121542 357234
rect 127826 362278 128062 362514
rect 128146 362278 128382 362514
rect 127826 361958 128062 362194
rect 128146 361958 128382 362194
rect 131546 365998 131782 366234
rect 131866 365998 132102 366234
rect 131546 365678 131782 365914
rect 131866 365678 132102 365914
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 156986 357318 157222 357554
rect 157306 357318 157542 357554
rect 156986 356998 157222 357234
rect 157306 356998 157542 357234
rect 163826 362278 164062 362514
rect 164146 362278 164382 362514
rect 163826 361958 164062 362194
rect 164146 361958 164382 362194
rect 167546 365998 167782 366234
rect 167866 365998 168102 366234
rect 167546 365678 167782 365914
rect 167866 365678 168102 365914
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 192986 357318 193222 357554
rect 193306 357318 193542 357554
rect 192986 356998 193222 357234
rect 193306 356998 193542 357234
rect 60328 345218 60564 345454
rect 60328 344898 60564 345134
rect 196056 345218 196292 345454
rect 196056 344898 196292 345134
rect 61008 327218 61244 327454
rect 61008 326898 61244 327134
rect 195376 327218 195612 327454
rect 195376 326898 195612 327134
rect 60328 309218 60564 309454
rect 60328 308898 60564 309134
rect 196056 309218 196292 309454
rect 196056 308898 196292 309134
rect 61008 291218 61244 291454
rect 61008 290898 61244 291134
rect 195376 291218 195612 291454
rect 195376 290898 195612 291134
rect 60328 273218 60564 273454
rect 60328 272898 60564 273134
rect 196056 273218 196292 273454
rect 196056 272898 196292 273134
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 84986 249318 85222 249554
rect 85306 249318 85542 249554
rect 84986 248998 85222 249234
rect 85306 248998 85542 249234
rect 91826 254278 92062 254514
rect 92146 254278 92382 254514
rect 91826 253958 92062 254194
rect 92146 253958 92382 254194
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 120986 249318 121222 249554
rect 121306 249318 121542 249554
rect 120986 248998 121222 249234
rect 121306 248998 121542 249234
rect 127826 254278 128062 254514
rect 128146 254278 128382 254514
rect 127826 253958 128062 254194
rect 128146 253958 128382 254194
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 249318 157222 249554
rect 157306 249318 157542 249554
rect 156986 248998 157222 249234
rect 157306 248998 157542 249234
rect 163826 254278 164062 254514
rect 164146 254278 164382 254514
rect 163826 253958 164062 254194
rect 164146 253958 164382 254194
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 249318 193222 249554
rect 193306 249318 193542 249554
rect 192986 248998 193222 249234
rect 193306 248998 193542 249234
rect 60328 237218 60564 237454
rect 60328 236898 60564 237134
rect 196056 237218 196292 237454
rect 196056 236898 196292 237134
rect 61008 219218 61244 219454
rect 61008 218898 61244 219134
rect 195376 219218 195612 219454
rect 195376 218898 195612 219134
rect 60328 201218 60564 201454
rect 60328 200898 60564 201134
rect 196056 201218 196292 201454
rect 196056 200898 196292 201134
rect 61008 183218 61244 183454
rect 61008 182898 61244 183134
rect 195376 183218 195612 183454
rect 195376 182898 195612 183134
rect 60328 165218 60564 165454
rect 60328 164898 60564 165134
rect 196056 165218 196292 165454
rect 196056 164898 196292 165134
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 137598 81502 137834
rect 81586 137598 81822 137834
rect 81266 137278 81502 137514
rect 81586 137278 81822 137514
rect 84986 141318 85222 141554
rect 85306 141318 85542 141554
rect 84986 140998 85222 141234
rect 85306 140998 85542 141234
rect 91826 146278 92062 146514
rect 92146 146278 92382 146514
rect 91826 145958 92062 146194
rect 92146 145958 92382 146194
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 137598 117502 137834
rect 117586 137598 117822 137834
rect 117266 137278 117502 137514
rect 117586 137278 117822 137514
rect 120986 141318 121222 141554
rect 121306 141318 121542 141554
rect 120986 140998 121222 141234
rect 121306 140998 121542 141234
rect 127826 146278 128062 146514
rect 128146 146278 128382 146514
rect 127826 145958 128062 146194
rect 128146 145958 128382 146194
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 153266 137598 153502 137834
rect 153586 137598 153822 137834
rect 153266 137278 153502 137514
rect 153586 137278 153822 137514
rect 156986 141318 157222 141554
rect 157306 141318 157542 141554
rect 156986 140998 157222 141234
rect 157306 140998 157542 141234
rect 163826 146278 164062 146514
rect 164146 146278 164382 146514
rect 163826 145958 164062 146194
rect 164146 145958 164382 146194
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 137598 189502 137834
rect 189586 137598 189822 137834
rect 189266 137278 189502 137514
rect 189586 137278 189822 137514
rect 192986 141318 193222 141554
rect 193306 141318 193542 141554
rect 192986 140998 193222 141234
rect 193306 140998 193542 141234
rect 61008 111218 61244 111454
rect 61008 110898 61244 111134
rect 195376 111218 195612 111454
rect 195376 110898 195612 111134
rect 60328 93218 60564 93454
rect 60328 92898 60564 93134
rect 196056 93218 196292 93454
rect 196056 92898 196292 93134
rect 61008 75218 61244 75454
rect 61008 74898 61244 75134
rect 195376 75218 195612 75454
rect 195376 74898 195612 75134
rect 60328 57218 60564 57454
rect 60328 56898 60564 57134
rect 196056 57218 196292 57454
rect 196056 56898 196292 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 362278 200062 362514
rect 200146 362278 200382 362514
rect 199826 361958 200062 362194
rect 200146 361958 200382 362194
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 254278 200062 254514
rect 200146 254278 200382 254514
rect 199826 253958 200062 254194
rect 200146 253958 200382 254194
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 146278 200062 146514
rect 200146 146278 200382 146514
rect 199826 145958 200062 146194
rect 200146 145958 200382 146194
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 203546 475878 203782 476114
rect 203866 475878 204102 476114
rect 203546 475558 203782 475794
rect 203866 475558 204102 475794
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 365998 203782 366234
rect 203866 365998 204102 366234
rect 203546 365678 203782 365914
rect 203866 365678 204102 365914
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 207266 477718 207502 477954
rect 207586 477718 207822 477954
rect 207266 477398 207502 477634
rect 207586 477398 207822 477634
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 475878 239782 476114
rect 239866 475878 240102 476114
rect 239546 475558 239782 475794
rect 239866 475558 240102 475794
rect 243266 477718 243502 477954
rect 243586 477718 243822 477954
rect 243266 477398 243502 477634
rect 243586 477398 243822 477634
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 275546 475878 275782 476114
rect 275866 475878 276102 476114
rect 275546 475558 275782 475794
rect 275866 475558 276102 475794
rect 279266 477718 279502 477954
rect 279586 477718 279822 477954
rect 279266 477398 279502 477634
rect 279586 477398 279822 477634
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 339610 633218 339846 633454
rect 339610 632898 339846 633134
rect 370330 633218 370566 633454
rect 370330 632898 370566 633134
rect 401050 633218 401286 633454
rect 401050 632898 401286 633134
rect 324250 615218 324486 615454
rect 324250 614898 324486 615134
rect 354970 615218 355206 615454
rect 354970 614898 355206 615134
rect 385690 615218 385926 615454
rect 385690 614898 385926 615134
rect 416410 615218 416646 615454
rect 416410 614898 416646 615134
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 339610 597218 339846 597454
rect 339610 596898 339846 597134
rect 370330 597218 370566 597454
rect 370330 596898 370566 597134
rect 401050 597218 401286 597454
rect 401050 596898 401286 597134
rect 324250 579218 324486 579454
rect 324250 578898 324486 579134
rect 354970 579218 355206 579454
rect 354970 578898 355206 579134
rect 385690 579218 385926 579454
rect 385690 578898 385926 579134
rect 416410 579218 416646 579454
rect 416410 578898 416646 579134
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 339610 561218 339846 561454
rect 339610 560898 339846 561134
rect 370330 561218 370566 561454
rect 370330 560898 370566 561134
rect 401050 561218 401286 561454
rect 401050 560898 401286 561134
rect 324250 543218 324486 543454
rect 324250 542898 324486 543134
rect 354970 543218 355206 543454
rect 354970 542898 355206 543134
rect 385690 543218 385926 543454
rect 385690 542898 385926 543134
rect 416410 543218 416646 543454
rect 416410 542898 416646 543134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221008 399218 221244 399454
rect 221008 398898 221244 399134
rect 355376 399218 355612 399454
rect 355376 398898 355612 399134
rect 220328 381218 220564 381454
rect 220328 380898 220564 381134
rect 356056 381218 356292 381454
rect 356056 380898 356292 381134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 228986 357318 229222 357554
rect 229306 357318 229542 357554
rect 228986 356998 229222 357234
rect 229306 356998 229542 357234
rect 235826 362278 236062 362514
rect 236146 362278 236382 362514
rect 235826 361958 236062 362194
rect 236146 361958 236382 362194
rect 239546 365998 239782 366234
rect 239866 365998 240102 366234
rect 239546 365678 239782 365914
rect 239866 365678 240102 365914
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 264986 357318 265222 357554
rect 265306 357318 265542 357554
rect 264986 356998 265222 357234
rect 265306 356998 265542 357234
rect 271826 362278 272062 362514
rect 272146 362278 272382 362514
rect 271826 361958 272062 362194
rect 272146 361958 272382 362194
rect 275546 365998 275782 366234
rect 275866 365998 276102 366234
rect 275546 365678 275782 365914
rect 275866 365678 276102 365914
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 300986 357318 301222 357554
rect 301306 357318 301542 357554
rect 300986 356998 301222 357234
rect 301306 356998 301542 357234
rect 307826 362278 308062 362514
rect 308146 362278 308382 362514
rect 307826 361958 308062 362194
rect 308146 361958 308382 362194
rect 311546 365998 311782 366234
rect 311866 365998 312102 366234
rect 311546 365678 311782 365914
rect 311866 365678 312102 365914
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 336986 357318 337222 357554
rect 337306 357318 337542 357554
rect 336986 356998 337222 357234
rect 337306 356998 337542 357234
rect 343826 362278 344062 362514
rect 344146 362278 344382 362514
rect 343826 361958 344062 362194
rect 344146 361958 344382 362194
rect 347546 365998 347782 366234
rect 347866 365998 348102 366234
rect 347546 365678 347782 365914
rect 347866 365678 348102 365914
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 220328 345218 220564 345454
rect 220328 344898 220564 345134
rect 356056 345218 356292 345454
rect 356056 344898 356292 345134
rect 221008 327218 221244 327454
rect 221008 326898 221244 327134
rect 355376 327218 355612 327454
rect 355376 326898 355612 327134
rect 220328 309218 220564 309454
rect 220328 308898 220564 309134
rect 356056 309218 356292 309454
rect 356056 308898 356292 309134
rect 221008 291218 221244 291454
rect 221008 290898 221244 291134
rect 355376 291218 355612 291454
rect 355376 290898 355612 291134
rect 220328 273218 220564 273454
rect 220328 272898 220564 273134
rect 356056 273218 356292 273454
rect 356056 272898 356292 273134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 249318 229222 249554
rect 229306 249318 229542 249554
rect 228986 248998 229222 249234
rect 229306 248998 229542 249234
rect 235826 254278 236062 254514
rect 236146 254278 236382 254514
rect 235826 253958 236062 254194
rect 236146 253958 236382 254194
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 264986 249318 265222 249554
rect 265306 249318 265542 249554
rect 264986 248998 265222 249234
rect 265306 248998 265542 249234
rect 271826 254278 272062 254514
rect 272146 254278 272382 254514
rect 271826 253958 272062 254194
rect 272146 253958 272382 254194
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 249318 301222 249554
rect 301306 249318 301542 249554
rect 300986 248998 301222 249234
rect 301306 248998 301542 249234
rect 307826 254278 308062 254514
rect 308146 254278 308382 254514
rect 307826 253958 308062 254194
rect 308146 253958 308382 254194
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 336986 249318 337222 249554
rect 337306 249318 337542 249554
rect 336986 248998 337222 249234
rect 337306 248998 337542 249234
rect 343826 254278 344062 254514
rect 344146 254278 344382 254514
rect 343826 253958 344062 254194
rect 344146 253958 344382 254194
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 220328 237218 220564 237454
rect 220328 236898 220564 237134
rect 356056 237218 356292 237454
rect 356056 236898 356292 237134
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 201218 220564 201454
rect 220328 200898 220564 201134
rect 356056 201218 356292 201454
rect 356056 200898 356292 201134
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 220328 165218 220564 165454
rect 220328 164898 220564 165134
rect 356056 165218 356292 165454
rect 356056 164898 356292 165134
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 137598 225502 137834
rect 225586 137598 225822 137834
rect 225266 137278 225502 137514
rect 225586 137278 225822 137514
rect 228986 141318 229222 141554
rect 229306 141318 229542 141554
rect 228986 140998 229222 141234
rect 229306 140998 229542 141234
rect 235826 146278 236062 146514
rect 236146 146278 236382 146514
rect 235826 145958 236062 146194
rect 236146 145958 236382 146194
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 137598 261502 137834
rect 261586 137598 261822 137834
rect 261266 137278 261502 137514
rect 261586 137278 261822 137514
rect 264986 141318 265222 141554
rect 265306 141318 265542 141554
rect 264986 140998 265222 141234
rect 265306 140998 265542 141234
rect 271826 146278 272062 146514
rect 272146 146278 272382 146514
rect 271826 145958 272062 146194
rect 272146 145958 272382 146194
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 137598 297502 137834
rect 297586 137598 297822 137834
rect 297266 137278 297502 137514
rect 297586 137278 297822 137514
rect 300986 141318 301222 141554
rect 301306 141318 301542 141554
rect 300986 140998 301222 141234
rect 301306 140998 301542 141234
rect 307826 146278 308062 146514
rect 308146 146278 308382 146514
rect 307826 145958 308062 146194
rect 308146 145958 308382 146194
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 137598 333502 137834
rect 333586 137598 333822 137834
rect 333266 137278 333502 137514
rect 333586 137278 333822 137514
rect 336986 141318 337222 141554
rect 337306 141318 337542 141554
rect 336986 140998 337222 141234
rect 337306 140998 337542 141234
rect 343826 146278 344062 146514
rect 344146 146278 344382 146514
rect 343826 145958 344062 146194
rect 344146 145958 344382 146194
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 221008 111218 221244 111454
rect 221008 110898 221244 111134
rect 355376 111218 355612 111454
rect 355376 110898 355612 111134
rect 220328 93218 220564 93454
rect 220328 92898 220564 93134
rect 356056 93218 356292 93454
rect 356056 92898 356292 93134
rect 221008 75218 221244 75454
rect 221008 74898 221244 75134
rect 355376 75218 355612 75454
rect 355376 74898 355612 75134
rect 220328 57218 220564 57454
rect 220328 56898 220564 57134
rect 356056 57218 356292 57454
rect 356056 56898 356292 57134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 137598 369502 137834
rect 369586 137598 369822 137834
rect 369266 137278 369502 137514
rect 369586 137278 369822 137514
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 357318 373222 357554
rect 373306 357318 373542 357554
rect 372986 356998 373222 357234
rect 373306 356998 373542 357234
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 249318 373222 249554
rect 373306 249318 373542 249554
rect 372986 248998 373222 249234
rect 373306 248998 373542 249234
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 141318 373222 141554
rect 373306 141318 373542 141554
rect 372986 140998 373222 141234
rect 373306 140998 373542 141234
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 479610 597218 479846 597454
rect 479610 596898 479846 597134
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 380328 453218 380564 453454
rect 380328 452898 380564 453134
rect 516056 453218 516292 453454
rect 516056 452898 516292 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 381008 435218 381244 435454
rect 381008 434898 381244 435134
rect 515376 435218 515612 435454
rect 515376 434898 515612 435134
rect 380328 417218 380564 417454
rect 380328 416898 380564 417134
rect 516056 417218 516292 417454
rect 516056 416898 516292 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 381008 399218 381244 399454
rect 381008 398898 381244 399134
rect 515376 399218 515612 399454
rect 515376 398898 515612 399134
rect 380328 381218 380564 381454
rect 380328 380898 380564 381134
rect 516056 381218 516292 381454
rect 516056 380898 516292 381134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 379826 362278 380062 362514
rect 380146 362278 380382 362514
rect 379826 361958 380062 362194
rect 380146 361958 380382 362194
rect 383546 365998 383782 366234
rect 383866 365998 384102 366234
rect 383546 365678 383782 365914
rect 383866 365678 384102 365914
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 408986 357318 409222 357554
rect 409306 357318 409542 357554
rect 408986 356998 409222 357234
rect 409306 356998 409542 357234
rect 415826 362278 416062 362514
rect 416146 362278 416382 362514
rect 415826 361958 416062 362194
rect 416146 361958 416382 362194
rect 419546 365998 419782 366234
rect 419866 365998 420102 366234
rect 419546 365678 419782 365914
rect 419866 365678 420102 365914
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 444986 357318 445222 357554
rect 445306 357318 445542 357554
rect 444986 356998 445222 357234
rect 445306 356998 445542 357234
rect 451826 362278 452062 362514
rect 452146 362278 452382 362514
rect 451826 361958 452062 362194
rect 452146 361958 452382 362194
rect 455546 365998 455782 366234
rect 455866 365998 456102 366234
rect 455546 365678 455782 365914
rect 455866 365678 456102 365914
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 480986 357318 481222 357554
rect 481306 357318 481542 357554
rect 480986 356998 481222 357234
rect 481306 356998 481542 357234
rect 487826 362278 488062 362514
rect 488146 362278 488382 362514
rect 487826 361958 488062 362194
rect 488146 361958 488382 362194
rect 491546 365998 491782 366234
rect 491866 365998 492102 366234
rect 491546 365678 491782 365914
rect 491866 365678 492102 365914
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 516986 357318 517222 357554
rect 517306 357318 517542 357554
rect 516986 356998 517222 357234
rect 517306 356998 517542 357234
rect 380328 345218 380564 345454
rect 380328 344898 380564 345134
rect 516056 345218 516292 345454
rect 516056 344898 516292 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 381008 327218 381244 327454
rect 381008 326898 381244 327134
rect 515376 327218 515612 327454
rect 515376 326898 515612 327134
rect 380328 309218 380564 309454
rect 380328 308898 380564 309134
rect 516056 309218 516292 309454
rect 516056 308898 516292 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 381008 291218 381244 291454
rect 381008 290898 381244 291134
rect 515376 291218 515612 291454
rect 515376 290898 515612 291134
rect 380328 273218 380564 273454
rect 380328 272898 380564 273134
rect 516056 273218 516292 273454
rect 516056 272898 516292 273134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 379826 254278 380062 254514
rect 380146 254278 380382 254514
rect 379826 253958 380062 254194
rect 380146 253958 380382 254194
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 408986 249318 409222 249554
rect 409306 249318 409542 249554
rect 408986 248998 409222 249234
rect 409306 248998 409542 249234
rect 415826 254278 416062 254514
rect 416146 254278 416382 254514
rect 415826 253958 416062 254194
rect 416146 253958 416382 254194
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 444986 249318 445222 249554
rect 445306 249318 445542 249554
rect 444986 248998 445222 249234
rect 445306 248998 445542 249234
rect 451826 254278 452062 254514
rect 452146 254278 452382 254514
rect 451826 253958 452062 254194
rect 452146 253958 452382 254194
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 249318 481222 249554
rect 481306 249318 481542 249554
rect 480986 248998 481222 249234
rect 481306 248998 481542 249234
rect 487826 254278 488062 254514
rect 488146 254278 488382 254514
rect 487826 253958 488062 254194
rect 488146 253958 488382 254194
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 249318 517222 249554
rect 517306 249318 517542 249554
rect 516986 248998 517222 249234
rect 517306 248998 517542 249234
rect 380328 237218 380564 237454
rect 380328 236898 380564 237134
rect 516056 237218 516292 237454
rect 516056 236898 516292 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 381008 219218 381244 219454
rect 381008 218898 381244 219134
rect 515376 219218 515612 219454
rect 515376 218898 515612 219134
rect 380328 201218 380564 201454
rect 380328 200898 380564 201134
rect 516056 201218 516292 201454
rect 516056 200898 516292 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 381008 183218 381244 183454
rect 381008 182898 381244 183134
rect 515376 183218 515612 183454
rect 515376 182898 515612 183134
rect 380328 165218 380564 165454
rect 380328 164898 380564 165134
rect 516056 165218 516292 165454
rect 516056 164898 516292 165134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 379826 146278 380062 146514
rect 380146 146278 380382 146514
rect 379826 145958 380062 146194
rect 380146 145958 380382 146194
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 137598 405502 137834
rect 405586 137598 405822 137834
rect 405266 137278 405502 137514
rect 405586 137278 405822 137514
rect 408986 141318 409222 141554
rect 409306 141318 409542 141554
rect 408986 140998 409222 141234
rect 409306 140998 409542 141234
rect 415826 146278 416062 146514
rect 416146 146278 416382 146514
rect 415826 145958 416062 146194
rect 416146 145958 416382 146194
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 137598 441502 137834
rect 441586 137598 441822 137834
rect 441266 137278 441502 137514
rect 441586 137278 441822 137514
rect 444986 141318 445222 141554
rect 445306 141318 445542 141554
rect 444986 140998 445222 141234
rect 445306 140998 445542 141234
rect 451826 146278 452062 146514
rect 452146 146278 452382 146514
rect 451826 145958 452062 146194
rect 452146 145958 452382 146194
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 137598 477502 137834
rect 477586 137598 477822 137834
rect 477266 137278 477502 137514
rect 477586 137278 477822 137514
rect 480986 141318 481222 141554
rect 481306 141318 481542 141554
rect 480986 140998 481222 141234
rect 481306 140998 481542 141234
rect 487826 146278 488062 146514
rect 488146 146278 488382 146514
rect 487826 145958 488062 146194
rect 488146 145958 488382 146194
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 137598 513502 137834
rect 513586 137598 513822 137834
rect 513266 137278 513502 137514
rect 513586 137278 513822 137514
rect 516986 141318 517222 141554
rect 517306 141318 517542 141554
rect 516986 140998 517222 141234
rect 517306 140998 517542 141234
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 381008 111218 381244 111454
rect 381008 110898 381244 111134
rect 515376 111218 515612 111454
rect 515376 110898 515612 111134
rect 380328 93218 380564 93454
rect 380328 92898 380564 93134
rect 516056 93218 516292 93454
rect 516056 92898 516292 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 381008 75218 381244 75454
rect 381008 74898 381244 75134
rect 515376 75218 515612 75454
rect 515376 74898 515612 75134
rect 380328 57218 380564 57454
rect 380328 56898 380564 57134
rect 516056 57218 516292 57454
rect 516056 56898 516292 57134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 79610 633454
rect 79846 633218 110330 633454
rect 110566 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 159610 633454
rect 159846 633218 190330 633454
rect 190566 633218 239610 633454
rect 239846 633218 270330 633454
rect 270566 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 339610 633454
rect 339846 633218 370330 633454
rect 370566 633218 401050 633454
rect 401286 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 79610 633134
rect 79846 632898 110330 633134
rect 110566 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 159610 633134
rect 159846 632898 190330 633134
rect 190566 632898 239610 633134
rect 239846 632898 270330 633134
rect 270566 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 339610 633134
rect 339846 632898 370330 633134
rect 370566 632898 401050 633134
rect 401286 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 144250 615454
rect 144486 615218 174970 615454
rect 175206 615218 224250 615454
rect 224486 615218 254970 615454
rect 255206 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 324250 615454
rect 324486 615218 354970 615454
rect 355206 615218 385690 615454
rect 385926 615218 416410 615454
rect 416646 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 144250 615134
rect 144486 614898 174970 615134
rect 175206 614898 224250 615134
rect 224486 614898 254970 615134
rect 255206 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 324250 615134
rect 324486 614898 354970 615134
rect 355206 614898 385690 615134
rect 385926 614898 416410 615134
rect 416646 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 79610 597454
rect 79846 597218 110330 597454
rect 110566 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 159610 597454
rect 159846 597218 190330 597454
rect 190566 597218 239610 597454
rect 239846 597218 270330 597454
rect 270566 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 339610 597454
rect 339846 597218 370330 597454
rect 370566 597218 401050 597454
rect 401286 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 479610 597454
rect 479846 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 79610 597134
rect 79846 596898 110330 597134
rect 110566 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 159610 597134
rect 159846 596898 190330 597134
rect 190566 596898 239610 597134
rect 239846 596898 270330 597134
rect 270566 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 339610 597134
rect 339846 596898 370330 597134
rect 370566 596898 401050 597134
rect 401286 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 479610 597134
rect 479846 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64250 579454
rect 64486 579218 94970 579454
rect 95206 579218 144250 579454
rect 144486 579218 174970 579454
rect 175206 579218 224250 579454
rect 224486 579218 254970 579454
rect 255206 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 324250 579454
rect 324486 579218 354970 579454
rect 355206 579218 385690 579454
rect 385926 579218 416410 579454
rect 416646 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64250 579134
rect 64486 578898 94970 579134
rect 95206 578898 144250 579134
rect 144486 578898 174970 579134
rect 175206 578898 224250 579134
rect 224486 578898 254970 579134
rect 255206 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 324250 579134
rect 324486 578898 354970 579134
rect 355206 578898 385690 579134
rect 385926 578898 416410 579134
rect 416646 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect 84954 571674 265574 571706
rect 84954 571438 84986 571674
rect 85222 571438 85306 571674
rect 85542 571438 120986 571674
rect 121222 571438 121306 571674
rect 121542 571438 156986 571674
rect 157222 571438 157306 571674
rect 157542 571438 192986 571674
rect 193222 571438 193306 571674
rect 193542 571438 228986 571674
rect 229222 571438 229306 571674
rect 229542 571438 264986 571674
rect 265222 571438 265306 571674
rect 265542 571438 265574 571674
rect 84954 571354 265574 571438
rect 84954 571118 84986 571354
rect 85222 571118 85306 571354
rect 85542 571118 120986 571354
rect 121222 571118 121306 571354
rect 121542 571118 156986 571354
rect 157222 571118 157306 571354
rect 157542 571118 192986 571354
rect 193222 571118 193306 571354
rect 193542 571118 228986 571354
rect 229222 571118 229306 571354
rect 229542 571118 264986 571354
rect 265222 571118 265306 571354
rect 265542 571118 265574 571354
rect 84954 571086 265574 571118
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect 81234 567954 261854 567986
rect 81234 567718 81266 567954
rect 81502 567718 81586 567954
rect 81822 567718 117266 567954
rect 117502 567718 117586 567954
rect 117822 567718 153266 567954
rect 153502 567718 153586 567954
rect 153822 567718 189266 567954
rect 189502 567718 189586 567954
rect 189822 567718 225266 567954
rect 225502 567718 225586 567954
rect 225822 567718 261266 567954
rect 261502 567718 261586 567954
rect 261822 567718 261854 567954
rect 81234 567634 261854 567718
rect 81234 567398 81266 567634
rect 81502 567398 81586 567634
rect 81822 567398 117266 567634
rect 117502 567398 117586 567634
rect 117822 567398 153266 567634
rect 153502 567398 153586 567634
rect 153822 567398 189266 567634
rect 189502 567398 189586 567634
rect 189822 567398 225266 567634
rect 225502 567398 225586 567634
rect 225822 567398 261266 567634
rect 261502 567398 261586 567634
rect 261822 567398 261854 567634
rect 81234 567366 261854 567398
rect 77514 566114 258134 566146
rect 77514 565878 77546 566114
rect 77782 565878 77866 566114
rect 78102 565878 113546 566114
rect 113782 565878 113866 566114
rect 114102 565878 149546 566114
rect 149782 565878 149866 566114
rect 150102 565878 185546 566114
rect 185782 565878 185866 566114
rect 186102 565878 221546 566114
rect 221782 565878 221866 566114
rect 222102 565878 257546 566114
rect 257782 565878 257866 566114
rect 258102 565878 258134 566114
rect 77514 565794 258134 565878
rect 77514 565558 77546 565794
rect 77782 565558 77866 565794
rect 78102 565558 113546 565794
rect 113782 565558 113866 565794
rect 114102 565558 149546 565794
rect 149782 565558 149866 565794
rect 150102 565558 185546 565794
rect 185782 565558 185866 565794
rect 186102 565558 221546 565794
rect 221782 565558 221866 565794
rect 222102 565558 257546 565794
rect 257782 565558 257866 565794
rect 258102 565558 258134 565794
rect 77514 565526 258134 565558
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect 73794 562394 254414 562426
rect 73794 562158 73826 562394
rect 74062 562158 74146 562394
rect 74382 562158 109826 562394
rect 110062 562158 110146 562394
rect 110382 562158 145826 562394
rect 146062 562158 146146 562394
rect 146382 562158 181826 562394
rect 182062 562158 182146 562394
rect 182382 562158 217826 562394
rect 218062 562158 218146 562394
rect 218382 562158 253826 562394
rect 254062 562158 254146 562394
rect 254382 562158 254414 562394
rect 73794 562074 254414 562158
rect 73794 561838 73826 562074
rect 74062 561838 74146 562074
rect 74382 561838 109826 562074
rect 110062 561838 110146 562074
rect 110382 561838 145826 562074
rect 146062 561838 146146 562074
rect 146382 561838 181826 562074
rect 182062 561838 182146 562074
rect 182382 561838 217826 562074
rect 218062 561838 218146 562074
rect 218382 561838 253826 562074
rect 254062 561838 254146 562074
rect 254382 561838 254414 562074
rect 73794 561806 254414 561838
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 339610 561454
rect 339846 561218 370330 561454
rect 370566 561218 401050 561454
rect 401286 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 339610 561134
rect 339846 560898 370330 561134
rect 370566 560898 401050 561134
rect 401286 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 64250 543454
rect 64486 543218 94970 543454
rect 95206 543218 125690 543454
rect 125926 543218 156410 543454
rect 156646 543218 187130 543454
rect 187366 543218 217850 543454
rect 218086 543218 248570 543454
rect 248806 543218 279290 543454
rect 279526 543218 324250 543454
rect 324486 543218 354970 543454
rect 355206 543218 385690 543454
rect 385926 543218 416410 543454
rect 416646 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 64250 543134
rect 64486 542898 94970 543134
rect 95206 542898 125690 543134
rect 125926 542898 156410 543134
rect 156646 542898 187130 543134
rect 187366 542898 217850 543134
rect 218086 542898 248570 543134
rect 248806 542898 279290 543134
rect 279526 542898 324250 543134
rect 324486 542898 354970 543134
rect 355206 542898 385690 543134
rect 385926 542898 416410 543134
rect 416646 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 79610 525454
rect 79846 525218 110330 525454
rect 110566 525218 141050 525454
rect 141286 525218 171770 525454
rect 172006 525218 202490 525454
rect 202726 525218 233210 525454
rect 233446 525218 263930 525454
rect 264166 525218 294650 525454
rect 294886 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 79610 525134
rect 79846 524898 110330 525134
rect 110566 524898 141050 525134
rect 141286 524898 171770 525134
rect 172006 524898 202490 525134
rect 202726 524898 233210 525134
rect 233446 524898 263930 525134
rect 264166 524898 294650 525134
rect 294886 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect 63234 477954 279854 477986
rect 63234 477718 63266 477954
rect 63502 477718 63586 477954
rect 63822 477718 99266 477954
rect 99502 477718 99586 477954
rect 99822 477718 135266 477954
rect 135502 477718 135586 477954
rect 135822 477718 171266 477954
rect 171502 477718 171586 477954
rect 171822 477718 207266 477954
rect 207502 477718 207586 477954
rect 207822 477718 243266 477954
rect 243502 477718 243586 477954
rect 243822 477718 279266 477954
rect 279502 477718 279586 477954
rect 279822 477718 279854 477954
rect 63234 477634 279854 477718
rect 63234 477398 63266 477634
rect 63502 477398 63586 477634
rect 63822 477398 99266 477634
rect 99502 477398 99586 477634
rect 99822 477398 135266 477634
rect 135502 477398 135586 477634
rect 135822 477398 171266 477634
rect 171502 477398 171586 477634
rect 171822 477398 207266 477634
rect 207502 477398 207586 477634
rect 207822 477398 243266 477634
rect 243502 477398 243586 477634
rect 243822 477398 279266 477634
rect 279502 477398 279586 477634
rect 279822 477398 279854 477634
rect 63234 477366 279854 477398
rect 59514 476114 276134 476146
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 59514 475794 276134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 59514 475526 276134 475558
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 380328 453454
rect 380564 453218 516056 453454
rect 516292 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 380328 453134
rect 380564 452898 516056 453134
rect 516292 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 381008 435454
rect 381244 435218 515376 435454
rect 515612 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 381008 435134
rect 381244 434898 515376 435134
rect 515612 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 380328 417454
rect 380564 417218 516056 417454
rect 516292 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 380328 417134
rect 380564 416898 516056 417134
rect 516292 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 61008 399454
rect 61244 399218 195376 399454
rect 195612 399218 221008 399454
rect 221244 399218 355376 399454
rect 355612 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 381008 399454
rect 381244 399218 515376 399454
rect 515612 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 61008 399134
rect 61244 398898 195376 399134
rect 195612 398898 221008 399134
rect 221244 398898 355376 399134
rect 355612 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 381008 399134
rect 381244 398898 515376 399134
rect 515612 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 60328 381454
rect 60564 381218 196056 381454
rect 196292 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 220328 381454
rect 220564 381218 356056 381454
rect 356292 381218 380328 381454
rect 380564 381218 516056 381454
rect 516292 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 60328 381134
rect 60564 380898 196056 381134
rect 196292 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 220328 381134
rect 220564 380898 356056 381134
rect 356292 380898 380328 381134
rect 380564 380898 516056 381134
rect 516292 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect 59514 366234 492134 366266
rect 59514 365998 59546 366234
rect 59782 365998 59866 366234
rect 60102 365998 95546 366234
rect 95782 365998 95866 366234
rect 96102 365998 131546 366234
rect 131782 365998 131866 366234
rect 132102 365998 167546 366234
rect 167782 365998 167866 366234
rect 168102 365998 203546 366234
rect 203782 365998 203866 366234
rect 204102 365998 239546 366234
rect 239782 365998 239866 366234
rect 240102 365998 275546 366234
rect 275782 365998 275866 366234
rect 276102 365998 311546 366234
rect 311782 365998 311866 366234
rect 312102 365998 347546 366234
rect 347782 365998 347866 366234
rect 348102 365998 383546 366234
rect 383782 365998 383866 366234
rect 384102 365998 419546 366234
rect 419782 365998 419866 366234
rect 420102 365998 455546 366234
rect 455782 365998 455866 366234
rect 456102 365998 491546 366234
rect 491782 365998 491866 366234
rect 492102 365998 492134 366234
rect 59514 365914 492134 365998
rect 59514 365678 59546 365914
rect 59782 365678 59866 365914
rect 60102 365678 95546 365914
rect 95782 365678 95866 365914
rect 96102 365678 131546 365914
rect 131782 365678 131866 365914
rect 132102 365678 167546 365914
rect 167782 365678 167866 365914
rect 168102 365678 203546 365914
rect 203782 365678 203866 365914
rect 204102 365678 239546 365914
rect 239782 365678 239866 365914
rect 240102 365678 275546 365914
rect 275782 365678 275866 365914
rect 276102 365678 311546 365914
rect 311782 365678 311866 365914
rect 312102 365678 347546 365914
rect 347782 365678 347866 365914
rect 348102 365678 383546 365914
rect 383782 365678 383866 365914
rect 384102 365678 419546 365914
rect 419782 365678 419866 365914
rect 420102 365678 455546 365914
rect 455782 365678 455866 365914
rect 456102 365678 491546 365914
rect 491782 365678 491866 365914
rect 492102 365678 492134 365914
rect 59514 365646 492134 365678
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect 91794 362514 488414 362546
rect 91794 362278 91826 362514
rect 92062 362278 92146 362514
rect 92382 362278 127826 362514
rect 128062 362278 128146 362514
rect 128382 362278 163826 362514
rect 164062 362278 164146 362514
rect 164382 362278 199826 362514
rect 200062 362278 200146 362514
rect 200382 362278 235826 362514
rect 236062 362278 236146 362514
rect 236382 362278 271826 362514
rect 272062 362278 272146 362514
rect 272382 362278 307826 362514
rect 308062 362278 308146 362514
rect 308382 362278 343826 362514
rect 344062 362278 344146 362514
rect 344382 362278 379826 362514
rect 380062 362278 380146 362514
rect 380382 362278 415826 362514
rect 416062 362278 416146 362514
rect 416382 362278 451826 362514
rect 452062 362278 452146 362514
rect 452382 362278 487826 362514
rect 488062 362278 488146 362514
rect 488382 362278 488414 362514
rect 91794 362194 488414 362278
rect 91794 361958 91826 362194
rect 92062 361958 92146 362194
rect 92382 361958 127826 362194
rect 128062 361958 128146 362194
rect 128382 361958 163826 362194
rect 164062 361958 164146 362194
rect 164382 361958 199826 362194
rect 200062 361958 200146 362194
rect 200382 361958 235826 362194
rect 236062 361958 236146 362194
rect 236382 361958 271826 362194
rect 272062 361958 272146 362194
rect 272382 361958 307826 362194
rect 308062 361958 308146 362194
rect 308382 361958 343826 362194
rect 344062 361958 344146 362194
rect 344382 361958 379826 362194
rect 380062 361958 380146 362194
rect 380382 361958 415826 362194
rect 416062 361958 416146 362194
rect 416382 361958 451826 362194
rect 452062 361958 452146 362194
rect 452382 361958 487826 362194
rect 488062 361958 488146 362194
rect 488382 361958 488414 362194
rect 91794 361926 488414 361958
rect 84954 357554 517574 357586
rect 84954 357318 84986 357554
rect 85222 357318 85306 357554
rect 85542 357318 120986 357554
rect 121222 357318 121306 357554
rect 121542 357318 156986 357554
rect 157222 357318 157306 357554
rect 157542 357318 192986 357554
rect 193222 357318 193306 357554
rect 193542 357318 228986 357554
rect 229222 357318 229306 357554
rect 229542 357318 264986 357554
rect 265222 357318 265306 357554
rect 265542 357318 300986 357554
rect 301222 357318 301306 357554
rect 301542 357318 336986 357554
rect 337222 357318 337306 357554
rect 337542 357318 372986 357554
rect 373222 357318 373306 357554
rect 373542 357318 408986 357554
rect 409222 357318 409306 357554
rect 409542 357318 444986 357554
rect 445222 357318 445306 357554
rect 445542 357318 480986 357554
rect 481222 357318 481306 357554
rect 481542 357318 516986 357554
rect 517222 357318 517306 357554
rect 517542 357318 517574 357554
rect 84954 357234 517574 357318
rect 84954 356998 84986 357234
rect 85222 356998 85306 357234
rect 85542 356998 120986 357234
rect 121222 356998 121306 357234
rect 121542 356998 156986 357234
rect 157222 356998 157306 357234
rect 157542 356998 192986 357234
rect 193222 356998 193306 357234
rect 193542 356998 228986 357234
rect 229222 356998 229306 357234
rect 229542 356998 264986 357234
rect 265222 356998 265306 357234
rect 265542 356998 300986 357234
rect 301222 356998 301306 357234
rect 301542 356998 336986 357234
rect 337222 356998 337306 357234
rect 337542 356998 372986 357234
rect 373222 356998 373306 357234
rect 373542 356998 408986 357234
rect 409222 356998 409306 357234
rect 409542 356998 444986 357234
rect 445222 356998 445306 357234
rect 445542 356998 480986 357234
rect 481222 356998 481306 357234
rect 481542 356998 516986 357234
rect 517222 356998 517306 357234
rect 517542 356998 517574 357234
rect 84954 356966 517574 356998
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 60328 345454
rect 60564 345218 196056 345454
rect 196292 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 220328 345454
rect 220564 345218 356056 345454
rect 356292 345218 380328 345454
rect 380564 345218 516056 345454
rect 516292 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 60328 345134
rect 60564 344898 196056 345134
rect 196292 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 220328 345134
rect 220564 344898 356056 345134
rect 356292 344898 380328 345134
rect 380564 344898 516056 345134
rect 516292 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 61008 327454
rect 61244 327218 195376 327454
rect 195612 327218 221008 327454
rect 221244 327218 355376 327454
rect 355612 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 381008 327454
rect 381244 327218 515376 327454
rect 515612 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 61008 327134
rect 61244 326898 195376 327134
rect 195612 326898 221008 327134
rect 221244 326898 355376 327134
rect 355612 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 381008 327134
rect 381244 326898 515376 327134
rect 515612 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 60328 309454
rect 60564 309218 196056 309454
rect 196292 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 220328 309454
rect 220564 309218 356056 309454
rect 356292 309218 380328 309454
rect 380564 309218 516056 309454
rect 516292 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 60328 309134
rect 60564 308898 196056 309134
rect 196292 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 220328 309134
rect 220564 308898 356056 309134
rect 356292 308898 380328 309134
rect 380564 308898 516056 309134
rect 516292 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 61008 291454
rect 61244 291218 195376 291454
rect 195612 291218 221008 291454
rect 221244 291218 355376 291454
rect 355612 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 381008 291454
rect 381244 291218 515376 291454
rect 515612 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 61008 291134
rect 61244 290898 195376 291134
rect 195612 290898 221008 291134
rect 221244 290898 355376 291134
rect 355612 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 381008 291134
rect 381244 290898 515376 291134
rect 515612 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 60328 273454
rect 60564 273218 196056 273454
rect 196292 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 220328 273454
rect 220564 273218 356056 273454
rect 356292 273218 380328 273454
rect 380564 273218 516056 273454
rect 516292 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 60328 273134
rect 60564 272898 196056 273134
rect 196292 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 220328 273134
rect 220564 272898 356056 273134
rect 356292 272898 380328 273134
rect 380564 272898 516056 273134
rect 516292 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect 91794 254514 488414 254546
rect 91794 254278 91826 254514
rect 92062 254278 92146 254514
rect 92382 254278 127826 254514
rect 128062 254278 128146 254514
rect 128382 254278 163826 254514
rect 164062 254278 164146 254514
rect 164382 254278 199826 254514
rect 200062 254278 200146 254514
rect 200382 254278 235826 254514
rect 236062 254278 236146 254514
rect 236382 254278 271826 254514
rect 272062 254278 272146 254514
rect 272382 254278 307826 254514
rect 308062 254278 308146 254514
rect 308382 254278 343826 254514
rect 344062 254278 344146 254514
rect 344382 254278 379826 254514
rect 380062 254278 380146 254514
rect 380382 254278 415826 254514
rect 416062 254278 416146 254514
rect 416382 254278 451826 254514
rect 452062 254278 452146 254514
rect 452382 254278 487826 254514
rect 488062 254278 488146 254514
rect 488382 254278 488414 254514
rect 91794 254194 488414 254278
rect 91794 253958 91826 254194
rect 92062 253958 92146 254194
rect 92382 253958 127826 254194
rect 128062 253958 128146 254194
rect 128382 253958 163826 254194
rect 164062 253958 164146 254194
rect 164382 253958 199826 254194
rect 200062 253958 200146 254194
rect 200382 253958 235826 254194
rect 236062 253958 236146 254194
rect 236382 253958 271826 254194
rect 272062 253958 272146 254194
rect 272382 253958 307826 254194
rect 308062 253958 308146 254194
rect 308382 253958 343826 254194
rect 344062 253958 344146 254194
rect 344382 253958 379826 254194
rect 380062 253958 380146 254194
rect 380382 253958 415826 254194
rect 416062 253958 416146 254194
rect 416382 253958 451826 254194
rect 452062 253958 452146 254194
rect 452382 253958 487826 254194
rect 488062 253958 488146 254194
rect 488382 253958 488414 254194
rect 91794 253926 488414 253958
rect 84954 249554 517574 249586
rect 84954 249318 84986 249554
rect 85222 249318 85306 249554
rect 85542 249318 120986 249554
rect 121222 249318 121306 249554
rect 121542 249318 156986 249554
rect 157222 249318 157306 249554
rect 157542 249318 192986 249554
rect 193222 249318 193306 249554
rect 193542 249318 228986 249554
rect 229222 249318 229306 249554
rect 229542 249318 264986 249554
rect 265222 249318 265306 249554
rect 265542 249318 300986 249554
rect 301222 249318 301306 249554
rect 301542 249318 336986 249554
rect 337222 249318 337306 249554
rect 337542 249318 372986 249554
rect 373222 249318 373306 249554
rect 373542 249318 408986 249554
rect 409222 249318 409306 249554
rect 409542 249318 444986 249554
rect 445222 249318 445306 249554
rect 445542 249318 480986 249554
rect 481222 249318 481306 249554
rect 481542 249318 516986 249554
rect 517222 249318 517306 249554
rect 517542 249318 517574 249554
rect 84954 249234 517574 249318
rect 84954 248998 84986 249234
rect 85222 248998 85306 249234
rect 85542 248998 120986 249234
rect 121222 248998 121306 249234
rect 121542 248998 156986 249234
rect 157222 248998 157306 249234
rect 157542 248998 192986 249234
rect 193222 248998 193306 249234
rect 193542 248998 228986 249234
rect 229222 248998 229306 249234
rect 229542 248998 264986 249234
rect 265222 248998 265306 249234
rect 265542 248998 300986 249234
rect 301222 248998 301306 249234
rect 301542 248998 336986 249234
rect 337222 248998 337306 249234
rect 337542 248998 372986 249234
rect 373222 248998 373306 249234
rect 373542 248998 408986 249234
rect 409222 248998 409306 249234
rect 409542 248998 444986 249234
rect 445222 248998 445306 249234
rect 445542 248998 480986 249234
rect 481222 248998 481306 249234
rect 481542 248998 516986 249234
rect 517222 248998 517306 249234
rect 517542 248998 517574 249234
rect 84954 248966 517574 248998
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 60328 237454
rect 60564 237218 196056 237454
rect 196292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 220328 237454
rect 220564 237218 356056 237454
rect 356292 237218 380328 237454
rect 380564 237218 516056 237454
rect 516292 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 60328 237134
rect 60564 236898 196056 237134
rect 196292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 220328 237134
rect 220564 236898 356056 237134
rect 356292 236898 380328 237134
rect 380564 236898 516056 237134
rect 516292 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 61008 219454
rect 61244 219218 195376 219454
rect 195612 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 381008 219454
rect 381244 219218 515376 219454
rect 515612 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 61008 219134
rect 61244 218898 195376 219134
rect 195612 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 381008 219134
rect 381244 218898 515376 219134
rect 515612 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 60328 201454
rect 60564 201218 196056 201454
rect 196292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 220328 201454
rect 220564 201218 356056 201454
rect 356292 201218 380328 201454
rect 380564 201218 516056 201454
rect 516292 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 60328 201134
rect 60564 200898 196056 201134
rect 196292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 220328 201134
rect 220564 200898 356056 201134
rect 356292 200898 380328 201134
rect 380564 200898 516056 201134
rect 516292 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 61008 183454
rect 61244 183218 195376 183454
rect 195612 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 381008 183454
rect 381244 183218 515376 183454
rect 515612 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 61008 183134
rect 61244 182898 195376 183134
rect 195612 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 381008 183134
rect 381244 182898 515376 183134
rect 515612 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 60328 165454
rect 60564 165218 196056 165454
rect 196292 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 220328 165454
rect 220564 165218 356056 165454
rect 356292 165218 380328 165454
rect 380564 165218 516056 165454
rect 516292 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 60328 165134
rect 60564 164898 196056 165134
rect 196292 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 220328 165134
rect 220564 164898 356056 165134
rect 356292 164898 380328 165134
rect 380564 164898 516056 165134
rect 516292 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect 91794 146514 488414 146546
rect 91794 146278 91826 146514
rect 92062 146278 92146 146514
rect 92382 146278 127826 146514
rect 128062 146278 128146 146514
rect 128382 146278 163826 146514
rect 164062 146278 164146 146514
rect 164382 146278 199826 146514
rect 200062 146278 200146 146514
rect 200382 146278 235826 146514
rect 236062 146278 236146 146514
rect 236382 146278 271826 146514
rect 272062 146278 272146 146514
rect 272382 146278 307826 146514
rect 308062 146278 308146 146514
rect 308382 146278 343826 146514
rect 344062 146278 344146 146514
rect 344382 146278 379826 146514
rect 380062 146278 380146 146514
rect 380382 146278 415826 146514
rect 416062 146278 416146 146514
rect 416382 146278 451826 146514
rect 452062 146278 452146 146514
rect 452382 146278 487826 146514
rect 488062 146278 488146 146514
rect 488382 146278 488414 146514
rect 91794 146194 488414 146278
rect 91794 145958 91826 146194
rect 92062 145958 92146 146194
rect 92382 145958 127826 146194
rect 128062 145958 128146 146194
rect 128382 145958 163826 146194
rect 164062 145958 164146 146194
rect 164382 145958 199826 146194
rect 200062 145958 200146 146194
rect 200382 145958 235826 146194
rect 236062 145958 236146 146194
rect 236382 145958 271826 146194
rect 272062 145958 272146 146194
rect 272382 145958 307826 146194
rect 308062 145958 308146 146194
rect 308382 145958 343826 146194
rect 344062 145958 344146 146194
rect 344382 145958 379826 146194
rect 380062 145958 380146 146194
rect 380382 145958 415826 146194
rect 416062 145958 416146 146194
rect 416382 145958 451826 146194
rect 452062 145958 452146 146194
rect 452382 145958 487826 146194
rect 488062 145958 488146 146194
rect 488382 145958 488414 146194
rect 91794 145926 488414 145958
rect 84954 141554 517574 141586
rect 84954 141318 84986 141554
rect 85222 141318 85306 141554
rect 85542 141318 120986 141554
rect 121222 141318 121306 141554
rect 121542 141318 156986 141554
rect 157222 141318 157306 141554
rect 157542 141318 192986 141554
rect 193222 141318 193306 141554
rect 193542 141318 228986 141554
rect 229222 141318 229306 141554
rect 229542 141318 264986 141554
rect 265222 141318 265306 141554
rect 265542 141318 300986 141554
rect 301222 141318 301306 141554
rect 301542 141318 336986 141554
rect 337222 141318 337306 141554
rect 337542 141318 372986 141554
rect 373222 141318 373306 141554
rect 373542 141318 408986 141554
rect 409222 141318 409306 141554
rect 409542 141318 444986 141554
rect 445222 141318 445306 141554
rect 445542 141318 480986 141554
rect 481222 141318 481306 141554
rect 481542 141318 516986 141554
rect 517222 141318 517306 141554
rect 517542 141318 517574 141554
rect 84954 141234 517574 141318
rect 84954 140998 84986 141234
rect 85222 140998 85306 141234
rect 85542 140998 120986 141234
rect 121222 140998 121306 141234
rect 121542 140998 156986 141234
rect 157222 140998 157306 141234
rect 157542 140998 192986 141234
rect 193222 140998 193306 141234
rect 193542 140998 228986 141234
rect 229222 140998 229306 141234
rect 229542 140998 264986 141234
rect 265222 140998 265306 141234
rect 265542 140998 300986 141234
rect 301222 140998 301306 141234
rect 301542 140998 336986 141234
rect 337222 140998 337306 141234
rect 337542 140998 372986 141234
rect 373222 140998 373306 141234
rect 373542 140998 408986 141234
rect 409222 140998 409306 141234
rect 409542 140998 444986 141234
rect 445222 140998 445306 141234
rect 445542 140998 480986 141234
rect 481222 140998 481306 141234
rect 481542 140998 516986 141234
rect 517222 140998 517306 141234
rect 517542 140998 517574 141234
rect 84954 140966 517574 140998
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect 81234 137834 513854 137866
rect 81234 137598 81266 137834
rect 81502 137598 81586 137834
rect 81822 137598 117266 137834
rect 117502 137598 117586 137834
rect 117822 137598 153266 137834
rect 153502 137598 153586 137834
rect 153822 137598 189266 137834
rect 189502 137598 189586 137834
rect 189822 137598 225266 137834
rect 225502 137598 225586 137834
rect 225822 137598 261266 137834
rect 261502 137598 261586 137834
rect 261822 137598 297266 137834
rect 297502 137598 297586 137834
rect 297822 137598 333266 137834
rect 333502 137598 333586 137834
rect 333822 137598 369266 137834
rect 369502 137598 369586 137834
rect 369822 137598 405266 137834
rect 405502 137598 405586 137834
rect 405822 137598 441266 137834
rect 441502 137598 441586 137834
rect 441822 137598 477266 137834
rect 477502 137598 477586 137834
rect 477822 137598 513266 137834
rect 513502 137598 513586 137834
rect 513822 137598 513854 137834
rect 81234 137514 513854 137598
rect 81234 137278 81266 137514
rect 81502 137278 81586 137514
rect 81822 137278 117266 137514
rect 117502 137278 117586 137514
rect 117822 137278 153266 137514
rect 153502 137278 153586 137514
rect 153822 137278 189266 137514
rect 189502 137278 189586 137514
rect 189822 137278 225266 137514
rect 225502 137278 225586 137514
rect 225822 137278 261266 137514
rect 261502 137278 261586 137514
rect 261822 137278 297266 137514
rect 297502 137278 297586 137514
rect 297822 137278 333266 137514
rect 333502 137278 333586 137514
rect 333822 137278 369266 137514
rect 369502 137278 369586 137514
rect 369822 137278 405266 137514
rect 405502 137278 405586 137514
rect 405822 137278 441266 137514
rect 441502 137278 441586 137514
rect 441822 137278 477266 137514
rect 477502 137278 477586 137514
rect 477822 137278 513266 137514
rect 513502 137278 513586 137514
rect 513822 137278 513854 137514
rect 81234 137246 513854 137278
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 61008 111454
rect 61244 111218 195376 111454
rect 195612 111218 221008 111454
rect 221244 111218 355376 111454
rect 355612 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 381008 111454
rect 381244 111218 515376 111454
rect 515612 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 61008 111134
rect 61244 110898 195376 111134
rect 195612 110898 221008 111134
rect 221244 110898 355376 111134
rect 355612 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 381008 111134
rect 381244 110898 515376 111134
rect 515612 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 60328 93454
rect 60564 93218 196056 93454
rect 196292 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 220328 93454
rect 220564 93218 356056 93454
rect 356292 93218 380328 93454
rect 380564 93218 516056 93454
rect 516292 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 60328 93134
rect 60564 92898 196056 93134
rect 196292 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 220328 93134
rect 220564 92898 356056 93134
rect 356292 92898 380328 93134
rect 380564 92898 516056 93134
rect 516292 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 61008 75454
rect 61244 75218 195376 75454
rect 195612 75218 221008 75454
rect 221244 75218 355376 75454
rect 355612 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 381008 75454
rect 381244 75218 515376 75454
rect 515612 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 61008 75134
rect 61244 74898 195376 75134
rect 195612 74898 221008 75134
rect 221244 74898 355376 75134
rect 355612 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 381008 75134
rect 381244 74898 515376 75134
rect 515612 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 60328 57454
rect 60564 57218 196056 57454
rect 196292 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 220328 57454
rect 220564 57218 356056 57454
rect 356292 57218 380328 57454
rect 380564 57218 516056 57454
rect 516292 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 60328 57134
rect 60564 56898 196056 57134
rect 196292 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 220328 57134
rect 220564 56898 356056 57134
rect 356292 56898 380328 57134
rect 380564 56898 516056 57134
rect 516292 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 45000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst1
timestamp 0
transform 1 0 60000 0 1 155000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst2
timestamp 0
transform 1 0 60000 0 1 265000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst0
timestamp 0
transform 1 0 380000 0 1 45000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst1
timestamp 0
transform 1 0 380000 0 1 155000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst2
timestamp 0
transform 1 0 380000 0 1 265000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst3
timestamp 0
transform 1 0 380000 0 1 375000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 375000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst1
timestamp 0
transform 1 0 220000 0 1 45000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst2
timestamp 0
transform 1 0 220000 0 1 155000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst3
timestamp 0
transform 1 0 220000 0 1 265000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst4
timestamp 0
transform 1 0 220000 0 1 375000
box 0 0 136620 83308
use VerySimpleCPU_core  inst_agent_1
timestamp 0
transform 1 0 60000 0 1 575000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_codemaker
timestamp 0
transform 1 0 220000 0 1 575000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_control_tower
timestamp 0
transform 1 0 140000 0 1 575000
box 0 0 60955 63099
use main_controller  inst_main_controller
timestamp 0
transform 1 0 60000 0 1 495000
box 0 0 240000 60000
use main_memory  inst_main_memory
timestamp 0
transform 1 0 320000 0 1 535000
box 0 0 108889 111033
use uart  inst_uart
timestamp 0
transform 1 0 460000 0 1 585000
box 0 0 50000 50000
<< labels >>
rlabel metal3 s 583520 275076 584960 275316 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 453274 703520 453386 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 391818 703520 391930 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 330362 703520 330474 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 268814 703520 268926 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 207358 703520 207470 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 145902 703520 146014 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 84446 703520 84558 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697492 480 697732 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 647172 480 647412 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 596988 480 597228 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 326212 584960 326452 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 546668 480 546908 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 496348 480 496588 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 446164 480 446404 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 395844 480 396084 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 345524 480 345764 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 295204 480 295444 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 245020 480 245260 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 194700 480 194940 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 144380 480 144620 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 377484 584960 377724 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 428620 584960 428860 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 479892 584960 480132 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 531028 584960 531268 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 582164 584960 582404 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 633436 584960 633676 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 576186 703520 576298 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 514730 703520 514842 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6340 584960 6580 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 441404 584960 441644 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 492676 584960 492916 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 543812 584960 544052 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 595084 584960 595324 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 646220 584960 646460 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 560822 703520 560934 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 499366 703520 499478 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 437910 703520 438022 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 376454 703520 376566 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 314998 703520 315110 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 44692 584960 44932 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 253450 703520 253562 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 191994 703520 192106 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 130538 703520 130650 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 69082 703520 69194 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684980 480 685220 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 634660 480 634900 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 584340 480 584580 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 534156 480 534396 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 483836 480 484076 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 433516 480 433756 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 83044 584960 83284 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 383196 480 383436 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 333012 480 333252 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 282692 480 282932 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 232372 480 232612 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 182188 480 182428 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 131868 480 132108 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 94196 480 94436 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 56388 480 56628 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 121396 584960 121636 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 159884 584960 160124 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 198236 584960 198476 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 236588 584960 236828 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 287860 584960 288100 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 338996 584960 339236 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 390268 584960 390508 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 31908 584960 32148 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 466972 584960 467212 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 518244 584960 518484 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 569380 584960 569620 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 620652 584960 620892 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 671788 584960 672028 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 530094 703520 530206 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 468638 703520 468750 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 407182 703520 407294 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 345726 703520 345838 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 284178 703520 284290 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 70260 584960 70500 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 222722 703520 222834 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 161266 703520 161378 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 99810 703520 99922 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 38354 703520 38466 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 659820 480 660060 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 609500 480 609740 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 559180 480 559420 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 508996 480 509236 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 458676 480 458916 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 408356 480 408596 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 108612 584960 108852 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 358172 480 358412 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 307852 480 308092 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 257532 480 257772 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 207212 480 207452 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 157028 480 157268 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 106708 480 106948 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 69036 480 69276 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 31228 480 31468 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 147100 584960 147340 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 185452 584960 185692 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 223804 584960 224044 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 262292 584960 262532 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 313428 584960 313668 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 364700 584960 364940 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 415836 584960 416076 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19124 584960 19364 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 454188 584960 454428 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 505460 584960 505700 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 556596 584960 556836 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 607868 584960 608108 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 659004 584960 659244 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 545458 703520 545570 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 484002 703520 484114 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 422546 703520 422658 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 361090 703520 361202 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 299634 703520 299746 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 57476 584960 57716 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 238086 703520 238198 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 176630 703520 176742 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 115174 703520 115286 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 53718 703520 53830 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 672332 480 672572 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 622148 480 622388 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 571828 480 572068 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 521508 480 521748 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 471188 480 471428 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 421004 480 421244 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 95828 584960 96068 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 370684 480 370924 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 320364 480 320604 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 270180 480 270420 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 219860 480 220100 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 169540 480 169780 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 119220 480 119460 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 81548 480 81788 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 43876 480 44116 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 134316 584960 134556 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 172668 584960 172908 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 211020 584960 211260 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 249508 584960 249748 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 300644 584960 300884 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 351780 584960 352020 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 403052 584960 403292 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125294 -960 125406 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 478574 -960 478686 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 482070 -960 482182 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 485566 -960 485678 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 489154 -960 489266 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 492650 -960 492762 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 496238 -960 496350 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 499734 -960 499846 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 503230 -960 503342 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 506818 -960 506930 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 510314 -960 510426 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 160622 -960 160734 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 513902 -960 514014 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 517398 -960 517510 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 520894 -960 521006 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 524482 -960 524594 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 527978 -960 528090 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 531566 -960 531678 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 535062 -960 535174 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 538558 -960 538670 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 542146 -960 542258 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 545642 -960 545754 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164118 -960 164230 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 549230 -960 549342 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 552726 -960 552838 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 556222 -960 556334 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 559810 -960 559922 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 563306 -960 563418 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 566894 -960 567006 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 570390 -960 570502 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 573886 -960 573998 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 167706 -960 167818 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171202 -960 171314 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 174790 -960 174902 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 178286 -960 178398 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 181782 -960 181894 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 185370 -960 185482 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 188866 -960 188978 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 192454 -960 192566 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 128882 -960 128994 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 195950 -960 196062 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 199446 -960 199558 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203034 -960 203146 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 206530 -960 206642 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210118 -960 210230 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 213614 -960 213726 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 217110 -960 217222 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 220698 -960 220810 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 224194 -960 224306 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 227782 -960 227894 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132378 -960 132490 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 231278 -960 231390 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 234774 -960 234886 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 238362 -960 238474 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 241858 -960 241970 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 245446 -960 245558 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 248942 -960 249054 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 252438 -960 252550 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 256026 -960 256138 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 259522 -960 259634 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 263110 -960 263222 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 135874 -960 135986 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 266606 -960 266718 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 270102 -960 270214 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 273690 -960 273802 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 277186 -960 277298 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 280774 -960 280886 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 298346 -960 298458 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 139462 -960 139574 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 305430 -960 305542 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 312514 -960 312626 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 316010 -960 316122 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 319598 -960 319710 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 323094 -960 323206 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 326682 -960 326794 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 330178 -960 330290 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 333674 -960 333786 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 142958 -960 143070 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 337262 -960 337374 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 340758 -960 340870 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 344346 -960 344458 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 358422 -960 358534 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 362010 -960 362122 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 365506 -960 365618 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 369002 -960 369114 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 146546 -960 146658 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 372590 -960 372702 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 376086 -960 376198 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 379674 -960 379786 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 383170 -960 383282 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 386666 -960 386778 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 390254 -960 390366 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 393750 -960 393862 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 397338 -960 397450 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 400834 -960 400946 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 404330 -960 404442 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150042 -960 150154 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 407918 -960 408030 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 411414 -960 411526 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 415002 -960 415114 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 418498 -960 418610 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 421994 -960 422106 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 425582 -960 425694 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 429078 -960 429190 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 432666 -960 432778 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 436162 -960 436274 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 439658 -960 439770 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 153538 -960 153650 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 443246 -960 443358 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 446742 -960 446854 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 450238 -960 450350 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 453826 -960 453938 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 457322 -960 457434 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 460910 -960 461022 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 474986 -960 475098 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157126 -960 157238 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126490 -960 126602 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 479678 -960 479790 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 483266 -960 483378 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 486762 -960 486874 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 490350 -960 490462 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 493846 -960 493958 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 497342 -960 497454 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 500930 -960 501042 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 504426 -960 504538 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 508014 -960 508126 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 511510 -960 511622 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 161818 -960 161930 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 515006 -960 515118 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 518594 -960 518706 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 522090 -960 522202 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 525678 -960 525790 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 529174 -960 529286 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 532670 -960 532782 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 536258 -960 536370 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 539754 -960 539866 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 543342 -960 543454 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 546838 -960 546950 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 165314 -960 165426 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 550334 -960 550446 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 553922 -960 554034 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 557418 -960 557530 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 561006 -960 561118 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 564502 -960 564614 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 567998 -960 568110 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 571586 -960 571698 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 575082 -960 575194 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 168902 -960 169014 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 172398 -960 172510 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 175894 -960 176006 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 179482 -960 179594 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 182978 -960 183090 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 186566 -960 186678 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190062 -960 190174 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 193558 -960 193670 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 129986 -960 130098 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197146 -960 197258 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 200642 -960 200754 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 204230 -960 204342 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 207726 -960 207838 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 211222 -960 211334 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 214810 -960 214922 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 218306 -960 218418 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 221894 -960 222006 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 225390 -960 225502 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 228886 -960 228998 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 133574 -960 133686 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 232474 -960 232586 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 235970 -960 236082 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 239558 -960 239670 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 243054 -960 243166 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 246550 -960 246662 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 250138 -960 250250 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 253634 -960 253746 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 257222 -960 257334 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 260718 -960 260830 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 264214 -960 264326 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137070 -960 137182 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 267802 -960 267914 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 271298 -960 271410 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 274886 -960 274998 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 278382 -960 278494 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 281878 -960 281990 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 285466 -960 285578 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 288962 -960 289074 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 292550 -960 292662 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 296046 -960 296158 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 299542 -960 299654 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 140658 -960 140770 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 303130 -960 303242 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 306626 -960 306738 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 310122 -960 310234 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 313710 -960 313822 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 317206 -960 317318 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 320794 -960 320906 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 324290 -960 324402 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 327786 -960 327898 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 331374 -960 331486 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 334870 -960 334982 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144154 -960 144266 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 338458 -960 338570 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 341954 -960 342066 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 359618 -960 359730 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 363114 -960 363226 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 366702 -960 366814 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 370198 -960 370310 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 147650 -960 147762 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 373786 -960 373898 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 377282 -960 377394 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 380778 -960 380890 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 384366 -960 384478 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 387862 -960 387974 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 391450 -960 391562 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 394946 -960 395058 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 398442 -960 398554 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 402030 -960 402142 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 405526 -960 405638 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151238 -960 151350 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 409114 -960 409226 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 412610 -960 412722 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 416106 -960 416218 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 419694 -960 419806 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 423190 -960 423302 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 426778 -960 426890 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 430274 -960 430386 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 433770 -960 433882 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 437358 -960 437470 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 440854 -960 440966 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 154734 -960 154846 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 444350 -960 444462 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 447938 -960 448050 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 451434 -960 451546 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 455022 -960 455134 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 458518 -960 458630 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 462014 -960 462126 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 465602 -960 465714 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 469098 -960 469210 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 472686 -960 472798 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 476182 -960 476294 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158230 -960 158342 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 127686 -960 127798 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 480874 -960 480986 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 484462 -960 484574 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 487958 -960 488070 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 491454 -960 491566 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 495042 -960 495154 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 498538 -960 498650 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 502126 -960 502238 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 505622 -960 505734 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 509118 -960 509230 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 512706 -960 512818 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163014 -960 163126 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 516202 -960 516314 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 519790 -960 519902 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 523286 -960 523398 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 526782 -960 526894 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 530370 -960 530482 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 533866 -960 533978 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 537454 -960 537566 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 540950 -960 541062 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 544446 -960 544558 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 548034 -960 548146 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 166510 -960 166622 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 551530 -960 551642 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 555118 -960 555230 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 558614 -960 558726 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 562110 -960 562222 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 565698 -960 565810 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 569194 -960 569306 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 572782 -960 572894 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170006 -960 170118 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 173594 -960 173706 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177090 -960 177202 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 180678 -960 180790 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184174 -960 184286 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 187670 -960 187782 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191258 -960 191370 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 194754 -960 194866 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131182 -960 131294 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 198342 -960 198454 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 201838 -960 201950 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 205334 -960 205446 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 208922 -960 209034 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 212418 -960 212530 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216006 -960 216118 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 219502 -960 219614 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 222998 -960 223110 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 226586 -960 226698 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 134770 -960 134882 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 240662 -960 240774 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 244250 -960 244362 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 247746 -960 247858 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 251334 -960 251446 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 254830 -960 254942 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 258326 -960 258438 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 261914 -960 262026 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 265410 -960 265522 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138266 -960 138378 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 268998 -960 269110 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 272494 -960 272606 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 275990 -960 276102 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 279578 -960 279690 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 283074 -960 283186 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 286662 -960 286774 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 290158 -960 290270 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 293654 -960 293766 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 297242 -960 297354 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 300738 -960 300850 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 141762 -960 141874 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 304234 -960 304346 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 307822 -960 307934 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 311318 -960 311430 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 314906 -960 315018 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 318402 -960 318514 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 321898 -960 322010 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 325486 -960 325598 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 328982 -960 329094 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 332570 -960 332682 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 336066 -960 336178 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145350 -960 145462 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 339562 -960 339674 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 343150 -960 343262 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 357226 -960 357338 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 360814 -960 360926 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 364310 -960 364422 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 367898 -960 368010 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 371394 -960 371506 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 148846 -960 148958 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 374890 -960 375002 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 378478 -960 378590 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 381974 -960 382086 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 385562 -960 385674 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 389058 -960 389170 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 392554 -960 392666 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 396142 -960 396254 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 399638 -960 399750 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 403226 -960 403338 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 406722 -960 406834 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152342 -960 152454 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 410218 -960 410330 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 413806 -960 413918 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 417302 -960 417414 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 420890 -960 421002 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 424386 -960 424498 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 427882 -960 427994 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 431470 -960 431582 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 434966 -960 435078 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 438554 -960 438666 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 442050 -960 442162 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 155930 -960 156042 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 445546 -960 445658 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 449134 -960 449246 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 452630 -960 452742 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 456126 -960 456238 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 459714 -960 459826 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 463210 -960 463322 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 466798 -960 466910 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 470294 -960 470406 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 473790 -960 473902 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 477378 -960 477490 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 159426 -960 159538 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 577474 -960 577586 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 578670 -960 578782 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 579774 -960 579886 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 580970 -960 581082 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s 73794 561806 254414 562426 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -1894 74414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -1894 110414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -1894 146414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -1894 182414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -1894 218414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -1894 254414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -1894 290414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -1894 326414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -1894 398414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -1894 434414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -1894 470414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -1894 506414 43000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 130308 74414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 130308 110414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 130308 146414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 130308 182414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 130308 218414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 130308 254414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 130308 290414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 130308 326414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 130308 398414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 130308 434414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 130308 470414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 130308 506414 153000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 240308 74414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 240308 110414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 240308 146414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 240308 182414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 240308 218414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 240308 254414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 240308 290414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 240308 326414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 240308 398414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 240308 434414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 240308 470414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 240308 506414 263000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 350308 74414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 350308 110414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 350308 146414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 350308 182414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 350308 218414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 350308 254414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 350308 290414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 350308 326414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 350308 398414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 350308 434414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 350308 470414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 350308 506414 373000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 460308 74414 493000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 460308 110414 493000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 460308 146414 493000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 460308 182414 493000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 460308 218414 493000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 460308 254414 493000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 460308 290414 493000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 460308 326414 533000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -1894 362414 533000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 460308 398414 533000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 557000 74414 573000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 557000 110414 573000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 557000 146414 573000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 557000 182414 573000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 557000 218414 573000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 557000 254414 573000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 460308 470414 583000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 460308 506414 583000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 640099 74414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 640099 110414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 640099 146414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 640099 182414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 640099 218414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 640099 254414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 557000 290414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 648033 326414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 648033 362414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 648033 398414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 460308 434414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 637000 470414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 637000 506414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power bidirectional
rlabel metal2 s 22990 703520 23102 704960 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 77514 565526 258134 566146 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 77514 -3814 78134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 113514 -3814 114134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149514 -3814 150134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 185514 -3814 186134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 221514 -3814 222134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 257514 -3814 258134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 293514 -3814 294134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 329514 -3814 330134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 401514 -3814 402134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 437514 -3814 438134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 473514 -3814 474134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 509514 -3814 510134 43000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 77514 130308 78134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 113514 130308 114134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149514 130308 150134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 185514 130308 186134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 221514 130308 222134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 257514 130308 258134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 293514 130308 294134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 329514 130308 330134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 401514 130308 402134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 437514 130308 438134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 473514 130308 474134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 509514 130308 510134 153000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 77514 240308 78134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 113514 240308 114134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149514 240308 150134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 185514 240308 186134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 221514 240308 222134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 257514 240308 258134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 293514 240308 294134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 329514 240308 330134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 401514 240308 402134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 437514 240308 438134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 473514 240308 474134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 509514 240308 510134 263000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 77514 350308 78134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 113514 350308 114134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149514 350308 150134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 185514 350308 186134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 221514 350308 222134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 257514 350308 258134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 293514 350308 294134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 329514 350308 330134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 401514 350308 402134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 437514 350308 438134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 473514 350308 474134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 509514 350308 510134 373000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 77514 460308 78134 493000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 113514 460308 114134 493000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149514 460308 150134 493000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 185514 460308 186134 493000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 221514 460308 222134 493000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 257514 460308 258134 493000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 293514 460308 294134 493000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 329514 460308 330134 533000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 365514 -3814 366134 533000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 401514 460308 402134 533000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 77514 557000 78134 573000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 113514 557000 114134 573000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149514 557000 150134 573000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 185514 557000 186134 573000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 221514 557000 222134 573000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 257514 557000 258134 573000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 473514 460308 474134 583000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 509514 460308 510134 583000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 77514 640099 78134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 113514 640099 114134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 149514 640099 150134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 185514 640099 186134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 221514 640099 222134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 257514 640099 258134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 293514 557000 294134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 329514 648033 330134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 365514 648033 366134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 401514 648033 402134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 437514 460308 438134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 473514 637000 474134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 509514 637000 510134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 533 nsew power bidirectional
rlabel metal2 s 582166 -960 582278 480 8 vccd2
port 534 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s 81234 137246 513854 137866 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s 81234 567366 261854 567986 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 535 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 81234 -5734 81854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 117234 -5734 117854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 153234 -5734 153854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 189234 -5734 189854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 225234 -5734 225854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 261234 -5734 261854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 297234 -5734 297854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 333234 -5734 333854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 405234 -5734 405854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 441234 -5734 441854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 477234 -5734 477854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 513234 -5734 513854 43000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 81234 130308 81854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 117234 130308 117854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 153234 130308 153854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 189234 130308 189854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 225234 130308 225854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 261234 130308 261854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 297234 130308 297854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 333234 130308 333854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 405234 130308 405854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 441234 130308 441854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 477234 130308 477854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 513234 130308 513854 153000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 81234 240308 81854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 117234 240308 117854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 153234 240308 153854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 189234 240308 189854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 225234 240308 225854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 261234 240308 261854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 297234 240308 297854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 333234 240308 333854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 405234 240308 405854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 441234 240308 441854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 477234 240308 477854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 513234 240308 513854 263000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 81234 350308 81854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 117234 350308 117854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 153234 350308 153854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 189234 350308 189854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 225234 350308 225854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 261234 350308 261854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 297234 350308 297854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 333234 350308 333854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 405234 350308 405854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 441234 350308 441854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 477234 350308 477854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 513234 350308 513854 373000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 81234 460308 81854 493000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 117234 460308 117854 493000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 153234 460308 153854 493000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 189234 460308 189854 493000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 225234 460308 225854 493000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 261234 460308 261854 493000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 297234 460308 297854 493000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 333234 460308 333854 533000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 369234 -5734 369854 533000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 405234 460308 405854 533000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 81234 557000 81854 573000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 117234 557000 117854 573000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 153234 557000 153854 573000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 189234 557000 189854 573000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 225234 557000 225854 573000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 261234 557000 261854 573000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 477234 460308 477854 583000 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 81234 640099 81854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 117234 640099 117854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 153234 640099 153854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 189234 640099 189854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 225234 640099 225854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 261234 640099 261854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 297234 557000 297854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 333234 648033 333854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 369234 648033 369854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 405234 648033 405854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 441234 460308 441854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 477234 637000 477854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 513234 460308 513854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 535 nsew power bidirectional
rlabel metal3 s 583520 684572 584960 684812 6 vdda1
port 536 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s 84954 140966 517574 141586 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s 84954 248966 517574 249586 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s 84954 356966 517574 357586 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s 84954 571086 265574 571706 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 537 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 84954 -7654 85574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 120954 -7654 121574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 156954 -7654 157574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 192954 -7654 193574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 228954 -7654 229574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 264954 -7654 265574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 300954 -7654 301574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 336954 -7654 337574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 408954 -7654 409574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 444954 -7654 445574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 480954 -7654 481574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 516954 -7654 517574 43000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 84954 130308 85574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 120954 130308 121574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 156954 130308 157574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 192954 130308 193574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 228954 130308 229574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 264954 130308 265574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 300954 130308 301574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 336954 130308 337574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 408954 130308 409574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 444954 130308 445574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 480954 130308 481574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 516954 130308 517574 153000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 84954 240308 85574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 120954 240308 121574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 156954 240308 157574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 192954 240308 193574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 228954 240308 229574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 264954 240308 265574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 300954 240308 301574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 336954 240308 337574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 408954 240308 409574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 444954 240308 445574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 480954 240308 481574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 516954 240308 517574 263000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 84954 350308 85574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 120954 350308 121574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 156954 350308 157574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 192954 350308 193574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 228954 350308 229574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 264954 350308 265574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 300954 350308 301574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 336954 350308 337574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 408954 350308 409574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 444954 350308 445574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 480954 350308 481574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 516954 350308 517574 373000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 84954 460308 85574 493000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 120954 460308 121574 493000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 156954 460308 157574 493000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 192954 460308 193574 493000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 228954 460308 229574 493000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 264954 460308 265574 493000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 300954 460308 301574 493000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 336954 460308 337574 533000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 372954 -7654 373574 533000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 408954 460308 409574 533000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 84954 557000 85574 573000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 120954 557000 121574 573000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 156954 557000 157574 573000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 192954 557000 193574 573000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 228954 557000 229574 573000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 264954 557000 265574 573000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 480954 460308 481574 583000 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 84954 640099 85574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 120954 640099 121574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 156954 640099 157574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 192954 640099 193574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 228954 640099 229574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 264954 640099 265574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 300954 557000 301574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 336954 648033 337574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 372954 648033 373574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 408954 648033 409574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 444954 460308 445574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 480954 637000 481574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 516954 460308 517574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 537 nsew power bidirectional
rlabel metal2 s 7626 703520 7738 704960 6 vdda2
port 538 nsew power bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s 63234 477366 279854 477986 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 539 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 63234 -5734 63854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 99234 -5734 99854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 135234 -5734 135854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 171234 -5734 171854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 243234 -5734 243854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 279234 -5734 279854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 315234 -5734 315854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 351234 -5734 351854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 387234 -5734 387854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 423234 -5734 423854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 459234 -5734 459854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 495234 -5734 495854 43000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 63234 130308 63854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 99234 130308 99854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 135234 130308 135854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 171234 130308 171854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 243234 130308 243854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 279234 130308 279854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 315234 130308 315854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 351234 130308 351854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 387234 130308 387854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 423234 130308 423854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 459234 130308 459854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 495234 130308 495854 153000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 63234 240308 63854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 99234 240308 99854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 135234 240308 135854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 171234 240308 171854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 243234 240308 243854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 279234 240308 279854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 315234 240308 315854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 351234 240308 351854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 387234 240308 387854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 423234 240308 423854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 459234 240308 459854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 495234 240308 495854 263000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 63234 350308 63854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 99234 350308 99854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 135234 350308 135854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 171234 350308 171854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 243234 350308 243854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 279234 350308 279854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 315234 350308 315854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 351234 350308 351854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 387234 350308 387854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 423234 350308 423854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 459234 350308 459854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 495234 350308 495854 373000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 63234 460308 63854 493000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 99234 460308 99854 493000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 135234 460308 135854 493000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 171234 460308 171854 493000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 207234 -5734 207854 493000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 243234 460308 243854 493000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 279234 460308 279854 493000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 351234 460308 351854 533000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 387234 460308 387854 533000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 423234 460308 423854 533000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 63234 557000 63854 573000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 99234 557000 99854 573000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 171234 557000 171854 573000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 243234 557000 243854 573000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 279234 557000 279854 573000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 459234 460308 459854 583000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 495234 460308 495854 583000 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 63234 640099 63854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 99234 640099 99854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 135234 557000 135854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 171234 640099 171854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 207234 557000 207854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 243234 640099 243854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 279234 640099 279854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 315234 460308 315854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 351234 648033 351854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 387234 648033 387854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 423234 648033 423854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 459234 637000 459854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 495234 637000 495854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 539 nsew ground bidirectional
rlabel metal2 s 583362 -960 583474 480 8 vssa1
port 540 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 541 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 66954 -7654 67574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 102954 -7654 103574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 138954 -7654 139574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 174954 -7654 175574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 246954 -7654 247574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 282954 -7654 283574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 318954 -7654 319574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 354954 -7654 355574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 390954 -7654 391574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 426954 -7654 427574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 462954 -7654 463574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 498954 -7654 499574 43000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 66954 130308 67574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 102954 130308 103574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 138954 130308 139574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 174954 130308 175574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 246954 130308 247574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 282954 130308 283574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 318954 130308 319574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 354954 130308 355574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 390954 130308 391574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 426954 130308 427574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 462954 130308 463574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 498954 130308 499574 153000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 66954 240308 67574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 102954 240308 103574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 138954 240308 139574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 174954 240308 175574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 246954 240308 247574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 282954 240308 283574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 318954 240308 319574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 354954 240308 355574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 390954 240308 391574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 426954 240308 427574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 462954 240308 463574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 498954 240308 499574 263000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 66954 350308 67574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 102954 350308 103574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 138954 350308 139574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 174954 350308 175574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 246954 350308 247574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 282954 350308 283574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 318954 350308 319574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 354954 350308 355574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 390954 350308 391574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 426954 350308 427574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 462954 350308 463574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 498954 350308 499574 373000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 66954 460308 67574 493000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 102954 460308 103574 493000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 138954 460308 139574 493000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 174954 460308 175574 493000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 210954 -7654 211574 493000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 246954 460308 247574 493000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 282954 460308 283574 493000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 318954 460308 319574 533000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 354954 460308 355574 533000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 390954 460308 391574 533000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 426954 460308 427574 533000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 66954 557000 67574 573000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 102954 557000 103574 573000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 138954 557000 139574 573000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 174954 557000 175574 573000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 246954 557000 247574 573000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 282954 557000 283574 573000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 462954 460308 463574 583000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 498954 460308 499574 583000 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 66954 640099 67574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 102954 640099 103574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 138954 640099 139574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 174954 640099 175574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 210954 557000 211574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 246954 640099 247574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 282954 640099 283574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 318954 648033 319574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 354954 648033 355574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 390954 648033 391574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 426954 648033 427574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 462954 637000 463574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 498954 637000 499574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 541 nsew ground bidirectional
rlabel metal3 s 583520 697356 584960 697596 6 vssa2
port 542 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s 91794 145926 488414 146546 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s 91794 253926 488414 254546 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s 91794 361926 488414 362546 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 543 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 91794 -1894 92414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 127794 -1894 128414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 163794 -1894 164414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 235794 -1894 236414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 271794 -1894 272414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 307794 -1894 308414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 343794 -1894 344414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 379794 -1894 380414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 415794 -1894 416414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 451794 -1894 452414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 487794 -1894 488414 43000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 91794 130308 92414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 127794 130308 128414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 163794 130308 164414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 235794 130308 236414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 271794 130308 272414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 307794 130308 308414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 343794 130308 344414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 379794 130308 380414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 415794 130308 416414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 451794 130308 452414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 487794 130308 488414 153000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 91794 240308 92414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 127794 240308 128414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 163794 240308 164414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 235794 240308 236414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 271794 240308 272414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 307794 240308 308414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 343794 240308 344414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 379794 240308 380414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 415794 240308 416414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 451794 240308 452414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 487794 240308 488414 263000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 91794 350308 92414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 127794 350308 128414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 163794 350308 164414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 235794 350308 236414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 271794 350308 272414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 307794 350308 308414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 343794 350308 344414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 379794 350308 380414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 415794 350308 416414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 451794 350308 452414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 487794 350308 488414 373000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 91794 460308 92414 493000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 127794 460308 128414 493000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 163794 460308 164414 493000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 199794 -1894 200414 493000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 235794 460308 236414 493000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 271794 460308 272414 493000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 343794 460308 344414 533000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 379794 460308 380414 533000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 415794 460308 416414 533000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 91794 557000 92414 573000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 163794 557000 164414 573000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 199794 557000 200414 573000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 235794 557000 236414 573000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 271794 557000 272414 573000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 487794 460308 488414 583000 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 91794 640099 92414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 127794 557000 128414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 163794 640099 164414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 199794 640099 200414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 235794 640099 236414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 271794 640099 272414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 307794 460308 308414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 343794 648033 344414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 379794 648033 380414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 415794 648033 416414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 451794 460308 452414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 487794 637000 488414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 543 nsew ground bidirectional
rlabel metal3 s -960 18716 480 18956 4 vssd1
port 544 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s 59514 365646 492134 366266 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s 59514 475526 276134 476146 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 545 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 59514 -3814 60134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 95514 -3814 96134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 131514 -3814 132134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 167514 -3814 168134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 239514 -3814 240134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 275514 -3814 276134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 311514 -3814 312134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 347514 -3814 348134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 383514 -3814 384134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 419514 -3814 420134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 455514 -3814 456134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 491514 -3814 492134 43000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 59514 130308 60134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 95514 130308 96134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 131514 130308 132134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 167514 130308 168134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 239514 130308 240134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 275514 130308 276134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 311514 130308 312134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 347514 130308 348134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 383514 130308 384134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 419514 130308 420134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 455514 130308 456134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 491514 130308 492134 153000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 59514 240308 60134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 95514 240308 96134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 131514 240308 132134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 167514 240308 168134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 239514 240308 240134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 275514 240308 276134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 311514 240308 312134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 347514 240308 348134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 383514 240308 384134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 419514 240308 420134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 455514 240308 456134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 491514 240308 492134 263000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 59514 350308 60134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 95514 350308 96134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 131514 350308 132134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 167514 350308 168134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 239514 350308 240134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 275514 350308 276134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 311514 350308 312134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 347514 350308 348134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 383514 350308 384134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 419514 350308 420134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 455514 350308 456134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 491514 350308 492134 373000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 59514 460308 60134 493000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 95514 460308 96134 493000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 131514 460308 132134 493000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 167514 460308 168134 493000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 203514 -3814 204134 493000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 239514 460308 240134 493000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 275514 460308 276134 493000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 347514 460308 348134 533000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 383514 460308 384134 533000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 419514 460308 420134 533000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 59514 557000 60134 573000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 95514 557000 96134 573000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 167514 557000 168134 573000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 239514 557000 240134 573000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 275514 557000 276134 573000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 491514 460308 492134 583000 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 59514 640099 60134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 95514 640099 96134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 131514 557000 132134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 167514 640099 168134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 203514 557000 204134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 239514 640099 240134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 275514 640099 276134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 311514 460308 312134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 347514 648033 348134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 383514 648033 384134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 419514 648033 420134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 455514 460308 456134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 491514 637000 492134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 545 nsew ground bidirectional
rlabel metal3 s -960 6204 480 6444 4 vssd2
port 546 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 547 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 548 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 549 nsew signal tristate
rlabel metal2 s 7534 -960 7646 480 8 wbs_adr_i[0]
port 550 nsew signal input
rlabel metal2 s 47554 -960 47666 480 8 wbs_adr_i[10]
port 551 nsew signal input
rlabel metal2 s 51142 -960 51254 480 8 wbs_adr_i[11]
port 552 nsew signal input
rlabel metal2 s 54638 -960 54750 480 8 wbs_adr_i[12]
port 553 nsew signal input
rlabel metal2 s 58226 -960 58338 480 8 wbs_adr_i[13]
port 554 nsew signal input
rlabel metal2 s 61722 -960 61834 480 8 wbs_adr_i[14]
port 555 nsew signal input
rlabel metal2 s 65218 -960 65330 480 8 wbs_adr_i[15]
port 556 nsew signal input
rlabel metal2 s 68806 -960 68918 480 8 wbs_adr_i[16]
port 557 nsew signal input
rlabel metal2 s 72302 -960 72414 480 8 wbs_adr_i[17]
port 558 nsew signal input
rlabel metal2 s 75890 -960 76002 480 8 wbs_adr_i[18]
port 559 nsew signal input
rlabel metal2 s 79386 -960 79498 480 8 wbs_adr_i[19]
port 560 nsew signal input
rlabel metal2 s 12226 -960 12338 480 8 wbs_adr_i[1]
port 561 nsew signal input
rlabel metal2 s 82882 -960 82994 480 8 wbs_adr_i[20]
port 562 nsew signal input
rlabel metal2 s 86470 -960 86582 480 8 wbs_adr_i[21]
port 563 nsew signal input
rlabel metal2 s 89966 -960 90078 480 8 wbs_adr_i[22]
port 564 nsew signal input
rlabel metal2 s 93554 -960 93666 480 8 wbs_adr_i[23]
port 565 nsew signal input
rlabel metal2 s 97050 -960 97162 480 8 wbs_adr_i[24]
port 566 nsew signal input
rlabel metal2 s 100546 -960 100658 480 8 wbs_adr_i[25]
port 567 nsew signal input
rlabel metal2 s 104134 -960 104246 480 8 wbs_adr_i[26]
port 568 nsew signal input
rlabel metal2 s 107630 -960 107742 480 8 wbs_adr_i[27]
port 569 nsew signal input
rlabel metal2 s 111218 -960 111330 480 8 wbs_adr_i[28]
port 570 nsew signal input
rlabel metal2 s 114714 -960 114826 480 8 wbs_adr_i[29]
port 571 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 572 nsew signal input
rlabel metal2 s 118210 -960 118322 480 8 wbs_adr_i[30]
port 573 nsew signal input
rlabel metal2 s 121798 -960 121910 480 8 wbs_adr_i[31]
port 574 nsew signal input
rlabel metal2 s 21702 -960 21814 480 8 wbs_adr_i[3]
port 575 nsew signal input
rlabel metal2 s 26394 -960 26506 480 8 wbs_adr_i[4]
port 576 nsew signal input
rlabel metal2 s 29890 -960 30002 480 8 wbs_adr_i[5]
port 577 nsew signal input
rlabel metal2 s 33478 -960 33590 480 8 wbs_adr_i[6]
port 578 nsew signal input
rlabel metal2 s 36974 -960 37086 480 8 wbs_adr_i[7]
port 579 nsew signal input
rlabel metal2 s 40562 -960 40674 480 8 wbs_adr_i[8]
port 580 nsew signal input
rlabel metal2 s 44058 -960 44170 480 8 wbs_adr_i[9]
port 581 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 582 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 583 nsew signal input
rlabel metal2 s 48750 -960 48862 480 8 wbs_dat_i[10]
port 584 nsew signal input
rlabel metal2 s 52338 -960 52450 480 8 wbs_dat_i[11]
port 585 nsew signal input
rlabel metal2 s 55834 -960 55946 480 8 wbs_dat_i[12]
port 586 nsew signal input
rlabel metal2 s 59330 -960 59442 480 8 wbs_dat_i[13]
port 587 nsew signal input
rlabel metal2 s 62918 -960 63030 480 8 wbs_dat_i[14]
port 588 nsew signal input
rlabel metal2 s 66414 -960 66526 480 8 wbs_dat_i[15]
port 589 nsew signal input
rlabel metal2 s 70002 -960 70114 480 8 wbs_dat_i[16]
port 590 nsew signal input
rlabel metal2 s 73498 -960 73610 480 8 wbs_dat_i[17]
port 591 nsew signal input
rlabel metal2 s 76994 -960 77106 480 8 wbs_dat_i[18]
port 592 nsew signal input
rlabel metal2 s 80582 -960 80694 480 8 wbs_dat_i[19]
port 593 nsew signal input
rlabel metal2 s 13422 -960 13534 480 8 wbs_dat_i[1]
port 594 nsew signal input
rlabel metal2 s 84078 -960 84190 480 8 wbs_dat_i[20]
port 595 nsew signal input
rlabel metal2 s 87666 -960 87778 480 8 wbs_dat_i[21]
port 596 nsew signal input
rlabel metal2 s 91162 -960 91274 480 8 wbs_dat_i[22]
port 597 nsew signal input
rlabel metal2 s 94658 -960 94770 480 8 wbs_dat_i[23]
port 598 nsew signal input
rlabel metal2 s 98246 -960 98358 480 8 wbs_dat_i[24]
port 599 nsew signal input
rlabel metal2 s 101742 -960 101854 480 8 wbs_dat_i[25]
port 600 nsew signal input
rlabel metal2 s 105330 -960 105442 480 8 wbs_dat_i[26]
port 601 nsew signal input
rlabel metal2 s 108826 -960 108938 480 8 wbs_dat_i[27]
port 602 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_dat_i[28]
port 603 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_dat_i[29]
port 604 nsew signal input
rlabel metal2 s 18114 -960 18226 480 8 wbs_dat_i[2]
port 605 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_dat_i[30]
port 606 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_dat_i[31]
port 607 nsew signal input
rlabel metal2 s 22898 -960 23010 480 8 wbs_dat_i[3]
port 608 nsew signal input
rlabel metal2 s 27590 -960 27702 480 8 wbs_dat_i[4]
port 609 nsew signal input
rlabel metal2 s 31086 -960 31198 480 8 wbs_dat_i[5]
port 610 nsew signal input
rlabel metal2 s 34674 -960 34786 480 8 wbs_dat_i[6]
port 611 nsew signal input
rlabel metal2 s 38170 -960 38282 480 8 wbs_dat_i[7]
port 612 nsew signal input
rlabel metal2 s 41666 -960 41778 480 8 wbs_dat_i[8]
port 613 nsew signal input
rlabel metal2 s 45254 -960 45366 480 8 wbs_dat_i[9]
port 614 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 615 nsew signal tristate
rlabel metal2 s 49946 -960 50058 480 8 wbs_dat_o[10]
port 616 nsew signal tristate
rlabel metal2 s 53442 -960 53554 480 8 wbs_dat_o[11]
port 617 nsew signal tristate
rlabel metal2 s 57030 -960 57142 480 8 wbs_dat_o[12]
port 618 nsew signal tristate
rlabel metal2 s 60526 -960 60638 480 8 wbs_dat_o[13]
port 619 nsew signal tristate
rlabel metal2 s 64114 -960 64226 480 8 wbs_dat_o[14]
port 620 nsew signal tristate
rlabel metal2 s 67610 -960 67722 480 8 wbs_dat_o[15]
port 621 nsew signal tristate
rlabel metal2 s 71106 -960 71218 480 8 wbs_dat_o[16]
port 622 nsew signal tristate
rlabel metal2 s 74694 -960 74806 480 8 wbs_dat_o[17]
port 623 nsew signal tristate
rlabel metal2 s 78190 -960 78302 480 8 wbs_dat_o[18]
port 624 nsew signal tristate
rlabel metal2 s 81778 -960 81890 480 8 wbs_dat_o[19]
port 625 nsew signal tristate
rlabel metal2 s 14618 -960 14730 480 8 wbs_dat_o[1]
port 626 nsew signal tristate
rlabel metal2 s 85274 -960 85386 480 8 wbs_dat_o[20]
port 627 nsew signal tristate
rlabel metal2 s 88770 -960 88882 480 8 wbs_dat_o[21]
port 628 nsew signal tristate
rlabel metal2 s 92358 -960 92470 480 8 wbs_dat_o[22]
port 629 nsew signal tristate
rlabel metal2 s 95854 -960 95966 480 8 wbs_dat_o[23]
port 630 nsew signal tristate
rlabel metal2 s 99442 -960 99554 480 8 wbs_dat_o[24]
port 631 nsew signal tristate
rlabel metal2 s 102938 -960 103050 480 8 wbs_dat_o[25]
port 632 nsew signal tristate
rlabel metal2 s 106434 -960 106546 480 8 wbs_dat_o[26]
port 633 nsew signal tristate
rlabel metal2 s 110022 -960 110134 480 8 wbs_dat_o[27]
port 634 nsew signal tristate
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_o[28]
port 635 nsew signal tristate
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_o[29]
port 636 nsew signal tristate
rlabel metal2 s 19310 -960 19422 480 8 wbs_dat_o[2]
port 637 nsew signal tristate
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_o[30]
port 638 nsew signal tristate
rlabel metal2 s 124098 -960 124210 480 8 wbs_dat_o[31]
port 639 nsew signal tristate
rlabel metal2 s 24002 -960 24114 480 8 wbs_dat_o[3]
port 640 nsew signal tristate
rlabel metal2 s 28786 -960 28898 480 8 wbs_dat_o[4]
port 641 nsew signal tristate
rlabel metal2 s 32282 -960 32394 480 8 wbs_dat_o[5]
port 642 nsew signal tristate
rlabel metal2 s 35778 -960 35890 480 8 wbs_dat_o[6]
port 643 nsew signal tristate
rlabel metal2 s 39366 -960 39478 480 8 wbs_dat_o[7]
port 644 nsew signal tristate
rlabel metal2 s 42862 -960 42974 480 8 wbs_dat_o[8]
port 645 nsew signal tristate
rlabel metal2 s 46450 -960 46562 480 8 wbs_dat_o[9]
port 646 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 647 nsew signal input
rlabel metal2 s 15814 -960 15926 480 8 wbs_sel_i[1]
port 648 nsew signal input
rlabel metal2 s 20506 -960 20618 480 8 wbs_sel_i[2]
port 649 nsew signal input
rlabel metal2 s 25198 -960 25310 480 8 wbs_sel_i[3]
port 650 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 651 nsew signal input
rlabel metal2 s 6338 -960 6450 480 8 wbs_we_i
port 652 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
