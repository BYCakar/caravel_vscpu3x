magic
tech sky130A
magscale 1 2
timestamp 1655490044
<< obsli1 >>
rect 61104 495159 509800 640401
<< obsm1 >>
rect 566 3408 580506 700528
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 580502 703610
rect 572 536 580502 703464
rect 710 480 1590 536
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6374 536
rect 6598 480 7570 536
rect 7794 480 8674 536
rect 8898 480 9870 536
rect 10094 480 11066 536
rect 11290 480 12262 536
rect 12486 480 13458 536
rect 13682 480 14654 536
rect 14878 480 15850 536
rect 16074 480 16954 536
rect 17178 480 18150 536
rect 18374 480 19346 536
rect 19570 480 20542 536
rect 20766 480 21738 536
rect 21962 480 22934 536
rect 23158 480 24130 536
rect 24354 480 25234 536
rect 25458 480 26430 536
rect 26654 480 27626 536
rect 27850 480 28822 536
rect 29046 480 30018 536
rect 30242 480 31214 536
rect 31438 480 32318 536
rect 32542 480 33514 536
rect 33738 480 34710 536
rect 34934 480 35906 536
rect 36130 480 37102 536
rect 37326 480 38298 536
rect 38522 480 39494 536
rect 39718 480 40598 536
rect 40822 480 41794 536
rect 42018 480 42990 536
rect 43214 480 44186 536
rect 44410 480 45382 536
rect 45606 480 46578 536
rect 46802 480 47774 536
rect 47998 480 48878 536
rect 49102 480 50074 536
rect 50298 480 51270 536
rect 51494 480 52466 536
rect 52690 480 53662 536
rect 53886 480 54858 536
rect 55082 480 55962 536
rect 56186 480 57158 536
rect 57382 480 58354 536
rect 58578 480 59550 536
rect 59774 480 60746 536
rect 60970 480 61942 536
rect 62166 480 63138 536
rect 63362 480 64242 536
rect 64466 480 65438 536
rect 65662 480 66634 536
rect 66858 480 67830 536
rect 68054 480 69026 536
rect 69250 480 70222 536
rect 70446 480 71418 536
rect 71642 480 72522 536
rect 72746 480 73718 536
rect 73942 480 74914 536
rect 75138 480 76110 536
rect 76334 480 77306 536
rect 77530 480 78502 536
rect 78726 480 79606 536
rect 79830 480 80802 536
rect 81026 480 81998 536
rect 82222 480 83194 536
rect 83418 480 84390 536
rect 84614 480 85586 536
rect 85810 480 86782 536
rect 87006 480 87886 536
rect 88110 480 89082 536
rect 89306 480 90278 536
rect 90502 480 91474 536
rect 91698 480 92670 536
rect 92894 480 93866 536
rect 94090 480 95062 536
rect 95286 480 96166 536
rect 96390 480 97362 536
rect 97586 480 98558 536
rect 98782 480 99754 536
rect 99978 480 100950 536
rect 101174 480 102146 536
rect 102370 480 103250 536
rect 103474 480 104446 536
rect 104670 480 105642 536
rect 105866 480 106838 536
rect 107062 480 108034 536
rect 108258 480 109230 536
rect 109454 480 110426 536
rect 110650 480 111530 536
rect 111754 480 112726 536
rect 112950 480 113922 536
rect 114146 480 115118 536
rect 115342 480 116314 536
rect 116538 480 117510 536
rect 117734 480 118706 536
rect 118930 480 119810 536
rect 120034 480 121006 536
rect 121230 480 122202 536
rect 122426 480 123398 536
rect 123622 480 124594 536
rect 124818 480 125790 536
rect 126014 480 126894 536
rect 127118 480 128090 536
rect 128314 480 129286 536
rect 129510 480 130482 536
rect 130706 480 131678 536
rect 131902 480 132874 536
rect 133098 480 134070 536
rect 134294 480 135174 536
rect 135398 480 136370 536
rect 136594 480 137566 536
rect 137790 480 138762 536
rect 138986 480 139958 536
rect 140182 480 141154 536
rect 141378 480 142350 536
rect 142574 480 143454 536
rect 143678 480 144650 536
rect 144874 480 145846 536
rect 146070 480 147042 536
rect 147266 480 148238 536
rect 148462 480 149434 536
rect 149658 480 150538 536
rect 150762 480 151734 536
rect 151958 480 152930 536
rect 153154 480 154126 536
rect 154350 480 155322 536
rect 155546 480 156518 536
rect 156742 480 157714 536
rect 157938 480 158818 536
rect 159042 480 160014 536
rect 160238 480 161210 536
rect 161434 480 162406 536
rect 162630 480 163602 536
rect 163826 480 164798 536
rect 165022 480 165994 536
rect 166218 480 167098 536
rect 167322 480 168294 536
rect 168518 480 169490 536
rect 169714 480 170686 536
rect 170910 480 171882 536
rect 172106 480 173078 536
rect 173302 480 174182 536
rect 174406 480 175378 536
rect 175602 480 176574 536
rect 176798 480 177770 536
rect 177994 480 178966 536
rect 179190 480 180162 536
rect 180386 480 181358 536
rect 181582 480 182462 536
rect 182686 480 183658 536
rect 183882 480 184854 536
rect 185078 480 186050 536
rect 186274 480 187246 536
rect 187470 480 188442 536
rect 188666 480 189638 536
rect 189862 480 190742 536
rect 190966 480 191938 536
rect 192162 480 193134 536
rect 193358 480 194330 536
rect 194554 480 195526 536
rect 195750 480 196722 536
rect 196946 480 197826 536
rect 198050 480 199022 536
rect 199246 480 200218 536
rect 200442 480 201414 536
rect 201638 480 202610 536
rect 202834 480 203806 536
rect 204030 480 205002 536
rect 205226 480 206106 536
rect 206330 480 207302 536
rect 207526 480 208498 536
rect 208722 480 209694 536
rect 209918 480 210890 536
rect 211114 480 212086 536
rect 212310 480 213282 536
rect 213506 480 214386 536
rect 214610 480 215582 536
rect 215806 480 216778 536
rect 217002 480 217974 536
rect 218198 480 219170 536
rect 219394 480 220366 536
rect 220590 480 221470 536
rect 221694 480 222666 536
rect 222890 480 223862 536
rect 224086 480 225058 536
rect 225282 480 226254 536
rect 226478 480 227450 536
rect 227674 480 228646 536
rect 228870 480 229750 536
rect 229974 480 230946 536
rect 231170 480 232142 536
rect 232366 480 233338 536
rect 233562 480 234534 536
rect 234758 480 235730 536
rect 235954 480 236926 536
rect 237150 480 238030 536
rect 238254 480 239226 536
rect 239450 480 240422 536
rect 240646 480 241618 536
rect 241842 480 242814 536
rect 243038 480 244010 536
rect 244234 480 245114 536
rect 245338 480 246310 536
rect 246534 480 247506 536
rect 247730 480 248702 536
rect 248926 480 249898 536
rect 250122 480 251094 536
rect 251318 480 252290 536
rect 252514 480 253394 536
rect 253618 480 254590 536
rect 254814 480 255786 536
rect 256010 480 256982 536
rect 257206 480 258178 536
rect 258402 480 259374 536
rect 259598 480 260570 536
rect 260794 480 261674 536
rect 261898 480 262870 536
rect 263094 480 264066 536
rect 264290 480 265262 536
rect 265486 480 266458 536
rect 266682 480 267654 536
rect 267878 480 268758 536
rect 268982 480 269954 536
rect 270178 480 271150 536
rect 271374 480 272346 536
rect 272570 480 273542 536
rect 273766 480 274738 536
rect 274962 480 275934 536
rect 276158 480 277038 536
rect 277262 480 278234 536
rect 278458 480 279430 536
rect 279654 480 280626 536
rect 280850 480 281822 536
rect 282046 480 283018 536
rect 283242 480 284214 536
rect 284438 480 285318 536
rect 285542 480 286514 536
rect 286738 480 287710 536
rect 287934 480 288906 536
rect 289130 480 290102 536
rect 290326 480 291298 536
rect 291522 480 292494 536
rect 292718 480 293598 536
rect 293822 480 294794 536
rect 295018 480 295990 536
rect 296214 480 297186 536
rect 297410 480 298382 536
rect 298606 480 299578 536
rect 299802 480 300682 536
rect 300906 480 301878 536
rect 302102 480 303074 536
rect 303298 480 304270 536
rect 304494 480 305466 536
rect 305690 480 306662 536
rect 306886 480 307858 536
rect 308082 480 308962 536
rect 309186 480 310158 536
rect 310382 480 311354 536
rect 311578 480 312550 536
rect 312774 480 313746 536
rect 313970 480 314942 536
rect 315166 480 316138 536
rect 316362 480 317242 536
rect 317466 480 318438 536
rect 318662 480 319634 536
rect 319858 480 320830 536
rect 321054 480 322026 536
rect 322250 480 323222 536
rect 323446 480 324326 536
rect 324550 480 325522 536
rect 325746 480 326718 536
rect 326942 480 327914 536
rect 328138 480 329110 536
rect 329334 480 330306 536
rect 330530 480 331502 536
rect 331726 480 332606 536
rect 332830 480 333802 536
rect 334026 480 334998 536
rect 335222 480 336194 536
rect 336418 480 337390 536
rect 337614 480 338586 536
rect 338810 480 339782 536
rect 340006 480 340886 536
rect 341110 480 342082 536
rect 342306 480 343278 536
rect 343502 480 344474 536
rect 344698 480 345670 536
rect 345894 480 346866 536
rect 347090 480 347970 536
rect 348194 480 349166 536
rect 349390 480 350362 536
rect 350586 480 351558 536
rect 351782 480 352754 536
rect 352978 480 353950 536
rect 354174 480 355146 536
rect 355370 480 356250 536
rect 356474 480 357446 536
rect 357670 480 358642 536
rect 358866 480 359838 536
rect 360062 480 361034 536
rect 361258 480 362230 536
rect 362454 480 363426 536
rect 363650 480 364530 536
rect 364754 480 365726 536
rect 365950 480 366922 536
rect 367146 480 368118 536
rect 368342 480 369314 536
rect 369538 480 370510 536
rect 370734 480 371614 536
rect 371838 480 372810 536
rect 373034 480 374006 536
rect 374230 480 375202 536
rect 375426 480 376398 536
rect 376622 480 377594 536
rect 377818 480 378790 536
rect 379014 480 379894 536
rect 380118 480 381090 536
rect 381314 480 382286 536
rect 382510 480 383482 536
rect 383706 480 384678 536
rect 384902 480 385874 536
rect 386098 480 387070 536
rect 387294 480 388174 536
rect 388398 480 389370 536
rect 389594 480 390566 536
rect 390790 480 391762 536
rect 391986 480 392958 536
rect 393182 480 394154 536
rect 394378 480 395258 536
rect 395482 480 396454 536
rect 396678 480 397650 536
rect 397874 480 398846 536
rect 399070 480 400042 536
rect 400266 480 401238 536
rect 401462 480 402434 536
rect 402658 480 403538 536
rect 403762 480 404734 536
rect 404958 480 405930 536
rect 406154 480 407126 536
rect 407350 480 408322 536
rect 408546 480 409518 536
rect 409742 480 410714 536
rect 410938 480 411818 536
rect 412042 480 413014 536
rect 413238 480 414210 536
rect 414434 480 415406 536
rect 415630 480 416602 536
rect 416826 480 417798 536
rect 418022 480 418902 536
rect 419126 480 420098 536
rect 420322 480 421294 536
rect 421518 480 422490 536
rect 422714 480 423686 536
rect 423910 480 424882 536
rect 425106 480 426078 536
rect 426302 480 427182 536
rect 427406 480 428378 536
rect 428602 480 429574 536
rect 429798 480 430770 536
rect 430994 480 431966 536
rect 432190 480 433162 536
rect 433386 480 434358 536
rect 434582 480 435462 536
rect 435686 480 436658 536
rect 436882 480 437854 536
rect 438078 480 439050 536
rect 439274 480 440246 536
rect 440470 480 441442 536
rect 441666 480 442546 536
rect 442770 480 443742 536
rect 443966 480 444938 536
rect 445162 480 446134 536
rect 446358 480 447330 536
rect 447554 480 448526 536
rect 448750 480 449722 536
rect 449946 480 450826 536
rect 451050 480 452022 536
rect 452246 480 453218 536
rect 453442 480 454414 536
rect 454638 480 455610 536
rect 455834 480 456806 536
rect 457030 480 458002 536
rect 458226 480 459106 536
rect 459330 480 460302 536
rect 460526 480 461498 536
rect 461722 480 462694 536
rect 462918 480 463890 536
rect 464114 480 465086 536
rect 465310 480 466190 536
rect 466414 480 467386 536
rect 467610 480 468582 536
rect 468806 480 469778 536
rect 470002 480 470974 536
rect 471198 480 472170 536
rect 472394 480 473366 536
rect 473590 480 474470 536
rect 474694 480 475666 536
rect 475890 480 476862 536
rect 477086 480 478058 536
rect 478282 480 479254 536
rect 479478 480 480450 536
rect 480674 480 481646 536
rect 481870 480 482750 536
rect 482974 480 483946 536
rect 484170 480 485142 536
rect 485366 480 486338 536
rect 486562 480 487534 536
rect 487758 480 488730 536
rect 488954 480 489834 536
rect 490058 480 491030 536
rect 491254 480 492226 536
rect 492450 480 493422 536
rect 493646 480 494618 536
rect 494842 480 495814 536
rect 496038 480 497010 536
rect 497234 480 498114 536
rect 498338 480 499310 536
rect 499534 480 500506 536
rect 500730 480 501702 536
rect 501926 480 502898 536
rect 503122 480 504094 536
rect 504318 480 505290 536
rect 505514 480 506394 536
rect 506618 480 507590 536
rect 507814 480 508786 536
rect 509010 480 509982 536
rect 510206 480 511178 536
rect 511402 480 512374 536
rect 512598 480 513478 536
rect 513702 480 514674 536
rect 514898 480 515870 536
rect 516094 480 517066 536
rect 517290 480 518262 536
rect 518486 480 519458 536
rect 519682 480 520654 536
rect 520878 480 521758 536
rect 521982 480 522954 536
rect 523178 480 524150 536
rect 524374 480 525346 536
rect 525570 480 526542 536
rect 526766 480 527738 536
rect 527962 480 528934 536
rect 529158 480 530038 536
rect 530262 480 531234 536
rect 531458 480 532430 536
rect 532654 480 533626 536
rect 533850 480 534822 536
rect 535046 480 536018 536
rect 536242 480 537122 536
rect 537346 480 538318 536
rect 538542 480 539514 536
rect 539738 480 540710 536
rect 540934 480 541906 536
rect 542130 480 543102 536
rect 543326 480 544298 536
rect 544522 480 545402 536
rect 545626 480 546598 536
rect 546822 480 547794 536
rect 548018 480 548990 536
rect 549214 480 550186 536
rect 550410 480 551382 536
rect 551606 480 552578 536
rect 552802 480 553682 536
rect 553906 480 554878 536
rect 555102 480 556074 536
rect 556298 480 557270 536
rect 557494 480 558466 536
rect 558690 480 559662 536
rect 559886 480 560766 536
rect 560990 480 561962 536
rect 562186 480 563158 536
rect 563382 480 564354 536
rect 564578 480 565550 536
rect 565774 480 566746 536
rect 566970 480 567942 536
rect 568166 480 569046 536
rect 569270 480 570242 536
rect 570466 480 571438 536
rect 571662 480 572634 536
rect 572858 480 573830 536
rect 574054 480 575026 536
rect 575250 480 576222 536
rect 576446 480 577326 536
rect 577550 480 578522 536
rect 578746 480 579718 536
rect 579942 480 580502 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 560 684084 583520 684317
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19588 583440 19988
rect 480 19580 583520 19588
rect 560 19180 583520 19580
rect 480 6796 583520 19180
rect 480 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 480 3299 583520 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 -5734 9854 709670
rect 11794 -1894 12414 705830
rect 12954 -7654 13574 711590
rect 15514 -3814 16134 707750
rect 19234 -5734 19854 709670
rect 21794 -1894 22414 705830
rect 22954 -7654 23574 711590
rect 25514 -3814 26134 707750
rect 29234 -5734 29854 709670
rect 31794 -1894 32414 705830
rect 32954 -7654 33574 711590
rect 35514 -3814 36134 707750
rect 39234 -5734 39854 709670
rect 41794 -1894 42414 705830
rect 42954 -7654 43574 711590
rect 45514 -3814 46134 707750
rect 49234 -5734 49854 709670
rect 51794 -1894 52414 705830
rect 52954 -7654 53574 711590
rect 55514 -3814 56134 707750
rect 59234 636033 59854 709670
rect 61794 636033 62414 705830
rect 62954 636033 63574 711590
rect 65514 636033 66134 707750
rect 69234 636033 69854 709670
rect 71794 636033 72414 705830
rect 72954 636033 73574 711590
rect 75514 636033 76134 707750
rect 79234 636033 79854 709670
rect 81794 636033 82414 705830
rect 82954 636033 83574 711590
rect 85514 636033 86134 707750
rect 89234 636033 89854 709670
rect 91794 636033 92414 705830
rect 92954 636033 93574 711590
rect 95514 636033 96134 707750
rect 99234 636033 99854 709670
rect 101794 636033 102414 705830
rect 102954 636033 103574 711590
rect 105514 636033 106134 707750
rect 109234 636033 109854 709670
rect 111794 636033 112414 705830
rect 112954 636033 113574 711590
rect 115514 636033 116134 707750
rect 119234 636033 119854 709670
rect 121794 636033 122414 705830
rect 122954 636033 123574 711590
rect 125514 636033 126134 707750
rect 129234 636033 129854 709670
rect 131794 636033 132414 705830
rect 132954 636033 133574 711590
rect 135514 636033 136134 707750
rect 139234 636033 139854 709670
rect 141794 636033 142414 705830
rect 142954 636033 143574 711590
rect 145514 636033 146134 707750
rect 149234 636033 149854 709670
rect 151794 636033 152414 705830
rect 152954 636033 153574 711590
rect 155514 636033 156134 707750
rect 159234 636033 159854 709670
rect 161794 636033 162414 705830
rect 162954 636033 163574 711590
rect 165514 636033 166134 707750
rect 169234 636033 169854 709670
rect 59234 466308 59854 521000
rect 61794 466308 62414 521000
rect 62954 466308 63574 521000
rect 65514 466308 66134 521000
rect 69234 466308 69854 521000
rect 71794 466308 72414 521000
rect 72954 466308 73574 521000
rect 75514 466308 76134 521000
rect 79234 466308 79854 521000
rect 81794 466308 82414 521000
rect 82954 466308 83574 521000
rect 85514 466308 86134 521000
rect 89234 466308 89854 521000
rect 91794 466308 92414 521000
rect 92954 466308 93574 521000
rect 95514 466308 96134 521000
rect 99234 466308 99854 521000
rect 101794 466308 102414 521000
rect 102954 466308 103574 521000
rect 105514 466308 106134 521000
rect 109234 466308 109854 521000
rect 111794 466308 112414 521000
rect 112954 466308 113574 521000
rect 115514 466308 116134 521000
rect 119234 466308 119854 521000
rect 121794 466308 122414 521000
rect 122954 466308 123574 521000
rect 125514 466308 126134 521000
rect 129234 466308 129854 521000
rect 131794 466308 132414 521000
rect 132954 466308 133574 521000
rect 135514 466308 136134 521000
rect 139234 466308 139854 521000
rect 141794 466308 142414 521000
rect 142954 466308 143574 521000
rect 145514 466308 146134 521000
rect 149234 466308 149854 521000
rect 151794 466308 152414 521000
rect 152954 466308 153574 521000
rect 155514 466308 156134 521000
rect 159234 466308 159854 521000
rect 161794 466308 162414 521000
rect 162954 466308 163574 521000
rect 165514 466308 166134 521000
rect 169234 466308 169854 521000
rect 171794 466308 172414 705830
rect 172954 466308 173574 711590
rect 175514 466308 176134 707750
rect 179234 466308 179854 709670
rect 181794 466308 182414 705830
rect 182954 466308 183574 711590
rect 185514 466308 186134 707750
rect 189234 466308 189854 709670
rect 191794 466308 192414 705830
rect 192954 466308 193574 711590
rect 195514 466308 196134 707750
rect 199234 642000 199854 709670
rect 201794 642000 202414 705830
rect 202954 642000 203574 711590
rect 205514 642000 206134 707750
rect 209234 642000 209854 709670
rect 211794 642000 212414 705830
rect 212954 642000 213574 711590
rect 215514 642000 216134 707750
rect 219234 642000 219854 709670
rect 221794 642000 222414 705830
rect 222954 642000 223574 711590
rect 225514 642000 226134 707750
rect 229234 642000 229854 709670
rect 231794 642000 232414 705830
rect 232954 642000 233574 711590
rect 235514 642000 236134 707750
rect 239234 642000 239854 709670
rect 241794 642000 242414 705830
rect 242954 642000 243574 711590
rect 245514 642000 246134 707750
rect 249234 642000 249854 709670
rect 251794 642000 252414 705830
rect 252954 642000 253574 711590
rect 255514 642000 256134 707750
rect 259234 642000 259854 709670
rect 261794 642000 262414 705830
rect 262954 642000 263574 711590
rect 265514 642000 266134 707750
rect 269234 642000 269854 709670
rect 271794 642000 272414 705830
rect 272954 642000 273574 711590
rect 275514 642000 276134 707750
rect 279234 642000 279854 709670
rect 281794 642000 282414 705830
rect 282954 642000 283574 711590
rect 285514 642000 286134 707750
rect 289234 642000 289854 709670
rect 291794 642000 292414 705830
rect 292954 642000 293574 711590
rect 295514 642000 296134 707750
rect 299234 642000 299854 709670
rect 301794 642000 302414 705830
rect 302954 642000 303574 711590
rect 305514 642000 306134 707750
rect 309234 642000 309854 709670
rect 311794 642000 312414 705830
rect 312954 642000 313574 711590
rect 315514 642000 316134 707750
rect 319234 642000 319854 709670
rect 321794 642000 322414 705830
rect 59234 359308 59854 379000
rect 61794 359308 62414 379000
rect 62954 359308 63574 379000
rect 65514 359308 66134 379000
rect 69234 359308 69854 379000
rect 71794 359308 72414 379000
rect 72954 359308 73574 379000
rect 75514 359308 76134 379000
rect 79234 359308 79854 379000
rect 81794 359308 82414 379000
rect 82954 359308 83574 379000
rect 85514 359308 86134 379000
rect 89234 359308 89854 379000
rect 91794 359308 92414 379000
rect 92954 359308 93574 379000
rect 95514 359308 96134 379000
rect 99234 359308 99854 379000
rect 101794 359308 102414 379000
rect 102954 359308 103574 379000
rect 105514 359308 106134 379000
rect 109234 359308 109854 379000
rect 111794 359308 112414 379000
rect 112954 359308 113574 379000
rect 115514 359308 116134 379000
rect 119234 359308 119854 379000
rect 121794 359308 122414 379000
rect 122954 359308 123574 379000
rect 125514 359308 126134 379000
rect 129234 359308 129854 379000
rect 131794 359308 132414 379000
rect 132954 359308 133574 379000
rect 135514 359308 136134 379000
rect 139234 359308 139854 379000
rect 141794 359308 142414 379000
rect 142954 359308 143574 379000
rect 145514 359308 146134 379000
rect 149234 359308 149854 379000
rect 151794 359308 152414 379000
rect 152954 359308 153574 379000
rect 155514 359308 156134 379000
rect 159234 359308 159854 379000
rect 161794 359308 162414 379000
rect 162954 359308 163574 379000
rect 165514 359308 166134 379000
rect 169234 359308 169854 379000
rect 171794 359308 172414 379000
rect 172954 359308 173574 379000
rect 175514 359308 176134 379000
rect 179234 359308 179854 379000
rect 181794 359308 182414 379000
rect 182954 359308 183574 379000
rect 185514 359308 186134 379000
rect 189234 359308 189854 379000
rect 191794 359308 192414 379000
rect 192954 359308 193574 379000
rect 195514 359308 196134 379000
rect 59234 252308 59854 272000
rect 61794 252308 62414 272000
rect 62954 252308 63574 272000
rect 65514 252308 66134 272000
rect 69234 252308 69854 272000
rect 71794 252308 72414 272000
rect 72954 252308 73574 272000
rect 75514 252308 76134 272000
rect 79234 252308 79854 272000
rect 81794 252308 82414 272000
rect 82954 252308 83574 272000
rect 85514 252308 86134 272000
rect 89234 252308 89854 272000
rect 91794 252308 92414 272000
rect 92954 252308 93574 272000
rect 95514 252308 96134 272000
rect 99234 252308 99854 272000
rect 101794 252308 102414 272000
rect 102954 252308 103574 272000
rect 105514 252308 106134 272000
rect 109234 252308 109854 272000
rect 111794 252308 112414 272000
rect 112954 252308 113574 272000
rect 115514 252308 116134 272000
rect 119234 252308 119854 272000
rect 121794 252308 122414 272000
rect 122954 252308 123574 272000
rect 125514 252308 126134 272000
rect 129234 252308 129854 272000
rect 131794 252308 132414 272000
rect 132954 252308 133574 272000
rect 135514 252308 136134 272000
rect 139234 252308 139854 272000
rect 141794 252308 142414 272000
rect 142954 252308 143574 272000
rect 145514 252308 146134 272000
rect 149234 252308 149854 272000
rect 151794 252308 152414 272000
rect 152954 252308 153574 272000
rect 155514 252308 156134 272000
rect 159234 252308 159854 272000
rect 161794 252308 162414 272000
rect 162954 252308 163574 272000
rect 165514 252308 166134 272000
rect 169234 252308 169854 272000
rect 171794 252308 172414 272000
rect 172954 252308 173574 272000
rect 175514 252308 176134 272000
rect 179234 252308 179854 272000
rect 181794 252308 182414 272000
rect 182954 252308 183574 272000
rect 185514 252308 186134 272000
rect 189234 252308 189854 272000
rect 191794 252308 192414 272000
rect 192954 252308 193574 272000
rect 195514 252308 196134 272000
rect 59234 145308 59854 165000
rect 61794 145308 62414 165000
rect 62954 145308 63574 165000
rect 65514 145308 66134 165000
rect 69234 145308 69854 165000
rect 71794 145308 72414 165000
rect 72954 145308 73574 165000
rect 75514 145308 76134 165000
rect 79234 145308 79854 165000
rect 81794 145308 82414 165000
rect 82954 145308 83574 165000
rect 85514 145308 86134 165000
rect 89234 145308 89854 165000
rect 91794 145308 92414 165000
rect 92954 145308 93574 165000
rect 95514 145308 96134 165000
rect 99234 145308 99854 165000
rect 101794 145308 102414 165000
rect 102954 145308 103574 165000
rect 105514 145308 106134 165000
rect 109234 145308 109854 165000
rect 111794 145308 112414 165000
rect 112954 145308 113574 165000
rect 115514 145308 116134 165000
rect 119234 145308 119854 165000
rect 121794 145308 122414 165000
rect 122954 145308 123574 165000
rect 125514 145308 126134 165000
rect 129234 145308 129854 165000
rect 131794 145308 132414 165000
rect 132954 145308 133574 165000
rect 135514 145308 136134 165000
rect 139234 145308 139854 165000
rect 141794 145308 142414 165000
rect 142954 145308 143574 165000
rect 145514 145308 146134 165000
rect 149234 145308 149854 165000
rect 151794 145308 152414 165000
rect 152954 145308 153574 165000
rect 155514 145308 156134 165000
rect 159234 145308 159854 165000
rect 161794 145308 162414 165000
rect 162954 145308 163574 165000
rect 165514 145308 166134 165000
rect 169234 145308 169854 165000
rect 171794 145308 172414 165000
rect 172954 145308 173574 165000
rect 175514 145308 176134 165000
rect 179234 145308 179854 165000
rect 181794 145308 182414 165000
rect 182954 145308 183574 165000
rect 185514 145308 186134 165000
rect 189234 145308 189854 165000
rect 191794 145308 192414 165000
rect 192954 145308 193574 165000
rect 195514 145308 196134 165000
rect 59234 -5734 59854 58000
rect 61794 -1894 62414 58000
rect 62954 -7654 63574 58000
rect 65514 -3814 66134 58000
rect 69234 -5734 69854 58000
rect 71794 -1894 72414 58000
rect 72954 -7654 73574 58000
rect 75514 -3814 76134 58000
rect 79234 -5734 79854 58000
rect 81794 -1894 82414 58000
rect 82954 -7654 83574 58000
rect 85514 -3814 86134 58000
rect 89234 -5734 89854 58000
rect 91794 -1894 92414 58000
rect 92954 -7654 93574 58000
rect 95514 -3814 96134 58000
rect 99234 -5734 99854 58000
rect 101794 -1894 102414 58000
rect 102954 -7654 103574 58000
rect 105514 -3814 106134 58000
rect 109234 -5734 109854 58000
rect 111794 -1894 112414 58000
rect 112954 -7654 113574 58000
rect 115514 -3814 116134 58000
rect 119234 -5734 119854 58000
rect 121794 -1894 122414 58000
rect 122954 -7654 123574 58000
rect 125514 -3814 126134 58000
rect 129234 -5734 129854 58000
rect 131794 -1894 132414 58000
rect 132954 -7654 133574 58000
rect 135514 -3814 136134 58000
rect 139234 -5734 139854 58000
rect 141794 -1894 142414 58000
rect 142954 -7654 143574 58000
rect 145514 -3814 146134 58000
rect 149234 -5734 149854 58000
rect 151794 -1894 152414 58000
rect 152954 -7654 153574 58000
rect 155514 -3814 156134 58000
rect 159234 -5734 159854 58000
rect 161794 -1894 162414 58000
rect 162954 -7654 163574 58000
rect 165514 -3814 166134 58000
rect 169234 -5734 169854 58000
rect 171794 -1894 172414 58000
rect 172954 -7654 173574 58000
rect 175514 -3814 176134 58000
rect 179234 -5734 179854 58000
rect 181794 -1894 182414 58000
rect 182954 -7654 183574 58000
rect 185514 -3814 186134 58000
rect 189234 -5734 189854 58000
rect 191794 -1894 192414 58000
rect 192954 -7654 193574 58000
rect 195514 -3814 196134 58000
rect 199234 -5734 199854 491000
rect 201794 -1894 202414 491000
rect 202954 -7654 203574 491000
rect 205514 -3814 206134 491000
rect 209234 -5734 209854 491000
rect 211794 -1894 212414 491000
rect 212954 -7654 213574 491000
rect 215514 -3814 216134 491000
rect 219234 466308 219854 491000
rect 221794 466308 222414 491000
rect 222954 466308 223574 491000
rect 225514 466308 226134 491000
rect 229234 466308 229854 491000
rect 231794 466308 232414 491000
rect 232954 466308 233574 491000
rect 235514 466308 236134 491000
rect 239234 466308 239854 491000
rect 241794 466308 242414 491000
rect 242954 466308 243574 491000
rect 245514 466308 246134 491000
rect 249234 466308 249854 491000
rect 251794 466308 252414 491000
rect 252954 466308 253574 491000
rect 255514 466308 256134 491000
rect 259234 466308 259854 491000
rect 261794 466308 262414 491000
rect 262954 466308 263574 491000
rect 265514 466308 266134 491000
rect 269234 466308 269854 491000
rect 271794 466308 272414 491000
rect 272954 466308 273574 491000
rect 275514 466308 276134 491000
rect 279234 466308 279854 491000
rect 281794 466308 282414 491000
rect 282954 466308 283574 491000
rect 285514 466308 286134 491000
rect 289234 466308 289854 491000
rect 291794 466308 292414 491000
rect 292954 466308 293574 491000
rect 295514 466308 296134 491000
rect 299234 466308 299854 491000
rect 301794 466308 302414 491000
rect 302954 466308 303574 491000
rect 305514 466308 306134 491000
rect 309234 466308 309854 491000
rect 311794 466308 312414 491000
rect 312954 466308 313574 491000
rect 315514 466308 316134 491000
rect 319234 466308 319854 491000
rect 321794 466308 322414 491000
rect 322954 466308 323574 711590
rect 325514 466308 326134 707750
rect 329234 466308 329854 709670
rect 331794 466308 332414 705830
rect 332954 466308 333574 711590
rect 335514 466308 336134 707750
rect 339234 466308 339854 709670
rect 341794 466308 342414 705830
rect 342954 466308 343574 711590
rect 345514 466308 346134 707750
rect 349234 466308 349854 709670
rect 351794 466308 352414 705830
rect 352954 645099 353574 711590
rect 355514 645099 356134 707750
rect 359234 645099 359854 709670
rect 361794 645099 362414 705830
rect 362954 645099 363574 711590
rect 365514 645099 366134 707750
rect 369234 645099 369854 709670
rect 371794 645099 372414 705830
rect 372954 645099 373574 711590
rect 375514 645099 376134 707750
rect 379234 645099 379854 709670
rect 381794 645099 382414 705830
rect 382954 645099 383574 711590
rect 385514 645099 386134 707750
rect 389234 645099 389854 709670
rect 391794 645099 392414 705830
rect 392954 645099 393574 711590
rect 395514 645099 396134 707750
rect 399234 645099 399854 709670
rect 401794 645099 402414 705830
rect 402954 645099 403574 711590
rect 405514 645099 406134 707750
rect 409234 645099 409854 709670
rect 411794 645099 412414 705830
rect 412954 645099 413574 711590
rect 415514 645099 416134 707750
rect 352954 558099 353574 578000
rect 355514 558099 356134 578000
rect 359234 558099 359854 578000
rect 361794 558099 362414 578000
rect 362954 558099 363574 578000
rect 365514 558099 366134 578000
rect 369234 558099 369854 578000
rect 371794 558099 372414 578000
rect 372954 558099 373574 578000
rect 375514 558099 376134 578000
rect 379234 558099 379854 578000
rect 381794 558099 382414 578000
rect 382954 558099 383574 578000
rect 385514 558099 386134 578000
rect 389234 558099 389854 578000
rect 391794 558099 392414 578000
rect 392954 558099 393574 578000
rect 395514 558099 396134 578000
rect 399234 558099 399854 578000
rect 401794 558099 402414 578000
rect 402954 558099 403574 578000
rect 405514 558099 406134 578000
rect 409234 558099 409854 578000
rect 411794 558099 412414 578000
rect 412954 558099 413574 578000
rect 415514 558099 416134 578000
rect 352954 466308 353574 491000
rect 355514 466308 356134 491000
rect 219234 359308 219854 379000
rect 221794 359308 222414 379000
rect 222954 359308 223574 379000
rect 225514 359308 226134 379000
rect 229234 359308 229854 379000
rect 231794 359308 232414 379000
rect 232954 359308 233574 379000
rect 235514 359308 236134 379000
rect 239234 359308 239854 379000
rect 241794 359308 242414 379000
rect 242954 359308 243574 379000
rect 245514 359308 246134 379000
rect 249234 359308 249854 379000
rect 251794 359308 252414 379000
rect 252954 359308 253574 379000
rect 255514 359308 256134 379000
rect 259234 359308 259854 379000
rect 261794 359308 262414 379000
rect 262954 359308 263574 379000
rect 265514 359308 266134 379000
rect 269234 359308 269854 379000
rect 271794 359308 272414 379000
rect 272954 359308 273574 379000
rect 275514 359308 276134 379000
rect 279234 359308 279854 379000
rect 281794 359308 282414 379000
rect 282954 359308 283574 379000
rect 285514 359308 286134 379000
rect 289234 359308 289854 379000
rect 291794 359308 292414 379000
rect 292954 359308 293574 379000
rect 295514 359308 296134 379000
rect 299234 359308 299854 379000
rect 301794 359308 302414 379000
rect 302954 359308 303574 379000
rect 305514 359308 306134 379000
rect 309234 359308 309854 379000
rect 311794 359308 312414 379000
rect 312954 359308 313574 379000
rect 315514 359308 316134 379000
rect 319234 359308 319854 379000
rect 321794 359308 322414 379000
rect 322954 359308 323574 379000
rect 325514 359308 326134 379000
rect 329234 359308 329854 379000
rect 331794 359308 332414 379000
rect 332954 359308 333574 379000
rect 335514 359308 336134 379000
rect 339234 359308 339854 379000
rect 341794 359308 342414 379000
rect 342954 359308 343574 379000
rect 345514 359308 346134 379000
rect 349234 359308 349854 379000
rect 351794 359308 352414 379000
rect 352954 359308 353574 379000
rect 355514 359308 356134 379000
rect 219234 252308 219854 272000
rect 221794 252308 222414 272000
rect 222954 252308 223574 272000
rect 225514 252308 226134 272000
rect 229234 252308 229854 272000
rect 231794 252308 232414 272000
rect 232954 252308 233574 272000
rect 235514 252308 236134 272000
rect 239234 252308 239854 272000
rect 241794 252308 242414 272000
rect 242954 252308 243574 272000
rect 245514 252308 246134 272000
rect 249234 252308 249854 272000
rect 251794 252308 252414 272000
rect 252954 252308 253574 272000
rect 255514 252308 256134 272000
rect 259234 252308 259854 272000
rect 261794 252308 262414 272000
rect 262954 252308 263574 272000
rect 265514 252308 266134 272000
rect 269234 252308 269854 272000
rect 271794 252308 272414 272000
rect 272954 252308 273574 272000
rect 275514 252308 276134 272000
rect 279234 252308 279854 272000
rect 281794 252308 282414 272000
rect 282954 252308 283574 272000
rect 285514 252308 286134 272000
rect 289234 252308 289854 272000
rect 291794 252308 292414 272000
rect 292954 252308 293574 272000
rect 295514 252308 296134 272000
rect 299234 252308 299854 272000
rect 301794 252308 302414 272000
rect 302954 252308 303574 272000
rect 305514 252308 306134 272000
rect 309234 252308 309854 272000
rect 311794 252308 312414 272000
rect 312954 252308 313574 272000
rect 315514 252308 316134 272000
rect 319234 252308 319854 272000
rect 321794 252308 322414 272000
rect 322954 252308 323574 272000
rect 325514 252308 326134 272000
rect 329234 252308 329854 272000
rect 331794 252308 332414 272000
rect 332954 252308 333574 272000
rect 335514 252308 336134 272000
rect 339234 252308 339854 272000
rect 341794 252308 342414 272000
rect 342954 252308 343574 272000
rect 345514 252308 346134 272000
rect 349234 252308 349854 272000
rect 351794 252308 352414 272000
rect 352954 252308 353574 272000
rect 355514 252308 356134 272000
rect 219234 145308 219854 165000
rect 221794 145308 222414 165000
rect 222954 145308 223574 165000
rect 225514 145308 226134 165000
rect 229234 145308 229854 165000
rect 231794 145308 232414 165000
rect 232954 145308 233574 165000
rect 235514 145308 236134 165000
rect 239234 145308 239854 165000
rect 241794 145308 242414 165000
rect 242954 145308 243574 165000
rect 245514 145308 246134 165000
rect 249234 145308 249854 165000
rect 251794 145308 252414 165000
rect 252954 145308 253574 165000
rect 255514 145308 256134 165000
rect 259234 145308 259854 165000
rect 261794 145308 262414 165000
rect 262954 145308 263574 165000
rect 265514 145308 266134 165000
rect 269234 145308 269854 165000
rect 271794 145308 272414 165000
rect 272954 145308 273574 165000
rect 275514 145308 276134 165000
rect 279234 145308 279854 165000
rect 281794 145308 282414 165000
rect 282954 145308 283574 165000
rect 285514 145308 286134 165000
rect 289234 145308 289854 165000
rect 291794 145308 292414 165000
rect 292954 145308 293574 165000
rect 295514 145308 296134 165000
rect 299234 145308 299854 165000
rect 301794 145308 302414 165000
rect 302954 145308 303574 165000
rect 305514 145308 306134 165000
rect 309234 145308 309854 165000
rect 311794 145308 312414 165000
rect 312954 145308 313574 165000
rect 315514 145308 316134 165000
rect 319234 145308 319854 165000
rect 321794 145308 322414 165000
rect 322954 145308 323574 165000
rect 325514 145308 326134 165000
rect 329234 145308 329854 165000
rect 331794 145308 332414 165000
rect 332954 145308 333574 165000
rect 335514 145308 336134 165000
rect 339234 145308 339854 165000
rect 341794 145308 342414 165000
rect 342954 145308 343574 165000
rect 345514 145308 346134 165000
rect 349234 145308 349854 165000
rect 351794 145308 352414 165000
rect 352954 145308 353574 165000
rect 355514 145308 356134 165000
rect 219234 -5734 219854 58000
rect 221794 -1894 222414 58000
rect 222954 -7654 223574 58000
rect 225514 -3814 226134 58000
rect 229234 -5734 229854 58000
rect 231794 -1894 232414 58000
rect 232954 -7654 233574 58000
rect 235514 -3814 236134 58000
rect 239234 -5734 239854 58000
rect 241794 -1894 242414 58000
rect 242954 -7654 243574 58000
rect 245514 -3814 246134 58000
rect 249234 -5734 249854 58000
rect 251794 -1894 252414 58000
rect 252954 -7654 253574 58000
rect 255514 -3814 256134 58000
rect 259234 -5734 259854 58000
rect 261794 -1894 262414 58000
rect 262954 -7654 263574 58000
rect 265514 -3814 266134 58000
rect 269234 -5734 269854 58000
rect 271794 -1894 272414 58000
rect 272954 -7654 273574 58000
rect 275514 -3814 276134 58000
rect 279234 -5734 279854 58000
rect 281794 -1894 282414 58000
rect 282954 -7654 283574 58000
rect 285514 -3814 286134 58000
rect 289234 -5734 289854 58000
rect 291794 -1894 292414 58000
rect 292954 -7654 293574 58000
rect 295514 -3814 296134 58000
rect 299234 -5734 299854 58000
rect 301794 -1894 302414 58000
rect 302954 -7654 303574 58000
rect 305514 -3814 306134 58000
rect 309234 -5734 309854 58000
rect 311794 -1894 312414 58000
rect 312954 -7654 313574 58000
rect 315514 -3814 316134 58000
rect 319234 -5734 319854 58000
rect 321794 -1894 322414 58000
rect 322954 -7654 323574 58000
rect 325514 -3814 326134 58000
rect 329234 -5734 329854 58000
rect 331794 -1894 332414 58000
rect 332954 -7654 333574 58000
rect 335514 -3814 336134 58000
rect 339234 -5734 339854 58000
rect 341794 -1894 342414 58000
rect 342954 -7654 343574 58000
rect 345514 -3814 346134 58000
rect 349234 -5734 349854 58000
rect 351794 -1894 352414 58000
rect 352954 -7654 353574 58000
rect 355514 -3814 356134 58000
rect 359234 -5734 359854 491000
rect 361794 -1894 362414 491000
rect 362954 -7654 363574 491000
rect 365514 -3814 366134 491000
rect 369234 -5734 369854 491000
rect 371794 -1894 372414 491000
rect 372954 -7654 373574 491000
rect 375514 -3814 376134 491000
rect 379234 466308 379854 491000
rect 381794 466308 382414 491000
rect 382954 466308 383574 491000
rect 385514 466308 386134 491000
rect 389234 466308 389854 491000
rect 391794 466308 392414 491000
rect 392954 466308 393574 491000
rect 395514 466308 396134 491000
rect 399234 466308 399854 491000
rect 401794 466308 402414 491000
rect 402954 466308 403574 491000
rect 405514 466308 406134 491000
rect 409234 466308 409854 491000
rect 411794 466308 412414 491000
rect 412954 466308 413574 491000
rect 415514 466308 416134 491000
rect 419234 466308 419854 709670
rect 421794 466308 422414 705830
rect 422954 466308 423574 711590
rect 425514 466308 426134 707750
rect 429234 466308 429854 709670
rect 431794 466308 432414 705830
rect 432954 466308 433574 711590
rect 435514 466308 436134 707750
rect 439234 466308 439854 709670
rect 441794 466308 442414 705830
rect 442954 466308 443574 711590
rect 445514 466308 446134 707750
rect 449234 645099 449854 709670
rect 451794 645099 452414 705830
rect 452954 645099 453574 711590
rect 455514 645099 456134 707750
rect 459234 645099 459854 709670
rect 461794 645099 462414 705830
rect 462954 645099 463574 711590
rect 465514 645099 466134 707750
rect 469234 645099 469854 709670
rect 471794 645099 472414 705830
rect 472954 645099 473574 711590
rect 475514 645099 476134 707750
rect 479234 645099 479854 709670
rect 481794 645099 482414 705830
rect 482954 645099 483574 711590
rect 485514 645099 486134 707750
rect 489234 645099 489854 709670
rect 491794 645099 492414 705830
rect 492954 645099 493574 711590
rect 495514 645099 496134 707750
rect 499234 645099 499854 709670
rect 501794 645099 502414 705830
rect 502954 645099 503574 711590
rect 505514 645099 506134 707750
rect 509234 645099 509854 709670
rect 511794 645099 512414 705830
rect 512954 645099 513574 711590
rect 449234 555000 449854 578000
rect 451794 555000 452414 578000
rect 452954 555000 453574 578000
rect 455514 555000 456134 578000
rect 459234 555000 459854 578000
rect 461794 555000 462414 578000
rect 462954 555000 463574 578000
rect 465514 555000 466134 578000
rect 469234 555000 469854 578000
rect 471794 555000 472414 578000
rect 472954 555000 473574 578000
rect 475514 555000 476134 578000
rect 479234 555000 479854 578000
rect 481794 555000 482414 578000
rect 482954 555000 483574 578000
rect 485514 555000 486134 578000
rect 489234 555000 489854 578000
rect 491794 555000 492414 578000
rect 492954 555000 493574 578000
rect 495514 555000 496134 578000
rect 499234 555000 499854 578000
rect 501794 555000 502414 578000
rect 449234 466308 449854 501000
rect 451794 466308 452414 501000
rect 452954 466308 453574 501000
rect 455514 466308 456134 501000
rect 459234 466308 459854 501000
rect 461794 466308 462414 501000
rect 462954 466308 463574 501000
rect 465514 466308 466134 501000
rect 469234 466308 469854 501000
rect 471794 466308 472414 501000
rect 472954 466308 473574 501000
rect 475514 466308 476134 501000
rect 479234 466308 479854 501000
rect 481794 466308 482414 501000
rect 482954 466308 483574 501000
rect 485514 466308 486134 501000
rect 489234 466308 489854 501000
rect 491794 466308 492414 501000
rect 492954 466308 493574 501000
rect 495514 466308 496134 501000
rect 499234 466308 499854 501000
rect 501794 466308 502414 501000
rect 502954 466308 503574 578000
rect 505514 466308 506134 578000
rect 509234 466308 509854 578000
rect 511794 466308 512414 578000
rect 512954 466308 513574 578000
rect 515514 466308 516134 707750
rect 379234 359308 379854 379000
rect 381794 359308 382414 379000
rect 382954 359308 383574 379000
rect 385514 359308 386134 379000
rect 389234 359308 389854 379000
rect 391794 359308 392414 379000
rect 392954 359308 393574 379000
rect 395514 359308 396134 379000
rect 399234 359308 399854 379000
rect 401794 359308 402414 379000
rect 402954 359308 403574 379000
rect 405514 359308 406134 379000
rect 409234 359308 409854 379000
rect 411794 359308 412414 379000
rect 412954 359308 413574 379000
rect 415514 359308 416134 379000
rect 419234 359308 419854 379000
rect 421794 359308 422414 379000
rect 422954 359308 423574 379000
rect 425514 359308 426134 379000
rect 429234 359308 429854 379000
rect 431794 359308 432414 379000
rect 432954 359308 433574 379000
rect 435514 359308 436134 379000
rect 439234 359308 439854 379000
rect 441794 359308 442414 379000
rect 442954 359308 443574 379000
rect 445514 359308 446134 379000
rect 449234 359308 449854 379000
rect 451794 359308 452414 379000
rect 452954 359308 453574 379000
rect 455514 359308 456134 379000
rect 459234 359308 459854 379000
rect 461794 359308 462414 379000
rect 462954 359308 463574 379000
rect 465514 359308 466134 379000
rect 469234 359308 469854 379000
rect 471794 359308 472414 379000
rect 472954 359308 473574 379000
rect 475514 359308 476134 379000
rect 479234 359308 479854 379000
rect 481794 359308 482414 379000
rect 482954 359308 483574 379000
rect 485514 359308 486134 379000
rect 489234 359308 489854 379000
rect 491794 359308 492414 379000
rect 492954 359308 493574 379000
rect 495514 359308 496134 379000
rect 499234 359308 499854 379000
rect 501794 359308 502414 379000
rect 502954 359308 503574 379000
rect 505514 359308 506134 379000
rect 509234 359308 509854 379000
rect 511794 359308 512414 379000
rect 512954 359308 513574 379000
rect 515514 359308 516134 379000
rect 379234 252308 379854 272000
rect 381794 252308 382414 272000
rect 382954 252308 383574 272000
rect 385514 252308 386134 272000
rect 389234 252308 389854 272000
rect 391794 252308 392414 272000
rect 392954 252308 393574 272000
rect 395514 252308 396134 272000
rect 399234 252308 399854 272000
rect 401794 252308 402414 272000
rect 402954 252308 403574 272000
rect 405514 252308 406134 272000
rect 409234 252308 409854 272000
rect 411794 252308 412414 272000
rect 412954 252308 413574 272000
rect 415514 252308 416134 272000
rect 419234 252308 419854 272000
rect 421794 252308 422414 272000
rect 422954 252308 423574 272000
rect 425514 252308 426134 272000
rect 429234 252308 429854 272000
rect 431794 252308 432414 272000
rect 432954 252308 433574 272000
rect 435514 252308 436134 272000
rect 439234 252308 439854 272000
rect 441794 252308 442414 272000
rect 442954 252308 443574 272000
rect 445514 252308 446134 272000
rect 449234 252308 449854 272000
rect 451794 252308 452414 272000
rect 452954 252308 453574 272000
rect 455514 252308 456134 272000
rect 459234 252308 459854 272000
rect 461794 252308 462414 272000
rect 462954 252308 463574 272000
rect 465514 252308 466134 272000
rect 469234 252308 469854 272000
rect 471794 252308 472414 272000
rect 472954 252308 473574 272000
rect 475514 252308 476134 272000
rect 479234 252308 479854 272000
rect 481794 252308 482414 272000
rect 482954 252308 483574 272000
rect 485514 252308 486134 272000
rect 489234 252308 489854 272000
rect 491794 252308 492414 272000
rect 492954 252308 493574 272000
rect 495514 252308 496134 272000
rect 499234 252308 499854 272000
rect 501794 252308 502414 272000
rect 502954 252308 503574 272000
rect 505514 252308 506134 272000
rect 509234 252308 509854 272000
rect 511794 252308 512414 272000
rect 512954 252308 513574 272000
rect 515514 252308 516134 272000
rect 379234 145308 379854 165000
rect 381794 145308 382414 165000
rect 382954 145308 383574 165000
rect 385514 145308 386134 165000
rect 389234 145308 389854 165000
rect 391794 145308 392414 165000
rect 392954 145308 393574 165000
rect 395514 145308 396134 165000
rect 399234 145308 399854 165000
rect 401794 145308 402414 165000
rect 402954 145308 403574 165000
rect 405514 145308 406134 165000
rect 409234 145308 409854 165000
rect 411794 145308 412414 165000
rect 412954 145308 413574 165000
rect 415514 145308 416134 165000
rect 419234 145308 419854 165000
rect 421794 145308 422414 165000
rect 422954 145308 423574 165000
rect 425514 145308 426134 165000
rect 429234 145308 429854 165000
rect 431794 145308 432414 165000
rect 432954 145308 433574 165000
rect 435514 145308 436134 165000
rect 439234 145308 439854 165000
rect 441794 145308 442414 165000
rect 442954 145308 443574 165000
rect 445514 145308 446134 165000
rect 449234 145308 449854 165000
rect 451794 145308 452414 165000
rect 452954 145308 453574 165000
rect 455514 145308 456134 165000
rect 459234 145308 459854 165000
rect 461794 145308 462414 165000
rect 462954 145308 463574 165000
rect 465514 145308 466134 165000
rect 469234 145308 469854 165000
rect 471794 145308 472414 165000
rect 472954 145308 473574 165000
rect 475514 145308 476134 165000
rect 479234 145308 479854 165000
rect 481794 145308 482414 165000
rect 482954 145308 483574 165000
rect 485514 145308 486134 165000
rect 489234 145308 489854 165000
rect 491794 145308 492414 165000
rect 492954 145308 493574 165000
rect 495514 145308 496134 165000
rect 499234 145308 499854 165000
rect 501794 145308 502414 165000
rect 502954 145308 503574 165000
rect 505514 145308 506134 165000
rect 509234 145308 509854 165000
rect 511794 145308 512414 165000
rect 512954 145308 513574 165000
rect 515514 145308 516134 165000
rect 379234 -5734 379854 58000
rect 381794 -1894 382414 58000
rect 382954 -7654 383574 58000
rect 385514 -3814 386134 58000
rect 389234 -5734 389854 58000
rect 391794 -1894 392414 58000
rect 392954 -7654 393574 58000
rect 395514 -3814 396134 58000
rect 399234 -5734 399854 58000
rect 401794 -1894 402414 58000
rect 402954 -7654 403574 58000
rect 405514 -3814 406134 58000
rect 409234 -5734 409854 58000
rect 411794 -1894 412414 58000
rect 412954 -7654 413574 58000
rect 415514 -3814 416134 58000
rect 419234 -5734 419854 58000
rect 421794 -1894 422414 58000
rect 422954 -7654 423574 58000
rect 425514 -3814 426134 58000
rect 429234 -5734 429854 58000
rect 431794 -1894 432414 58000
rect 432954 -7654 433574 58000
rect 435514 -3814 436134 58000
rect 439234 -5734 439854 58000
rect 441794 -1894 442414 58000
rect 442954 -7654 443574 58000
rect 445514 -3814 446134 58000
rect 449234 -5734 449854 58000
rect 451794 -1894 452414 58000
rect 452954 -7654 453574 58000
rect 455514 -3814 456134 58000
rect 459234 -5734 459854 58000
rect 461794 -1894 462414 58000
rect 462954 -7654 463574 58000
rect 465514 -3814 466134 58000
rect 469234 -5734 469854 58000
rect 471794 -1894 472414 58000
rect 472954 -7654 473574 58000
rect 475514 -3814 476134 58000
rect 479234 -5734 479854 58000
rect 481794 -1894 482414 58000
rect 482954 -7654 483574 58000
rect 485514 -3814 486134 58000
rect 489234 -5734 489854 58000
rect 491794 -1894 492414 58000
rect 492954 -7654 493574 58000
rect 495514 -3814 496134 58000
rect 499234 -5734 499854 58000
rect 501794 -1894 502414 58000
rect 502954 -7654 503574 58000
rect 505514 -3814 506134 58000
rect 509234 -5734 509854 58000
rect 511794 -1894 512414 58000
rect 512954 -7654 513574 58000
rect 515514 -3814 516134 58000
rect 519234 -5734 519854 709670
rect 521794 -1894 522414 705830
rect 522954 -7654 523574 711590
rect 525514 -3814 526134 707750
rect 529234 -5734 529854 709670
rect 531794 -1894 532414 705830
rect 532954 -7654 533574 711590
rect 535514 -3814 536134 707750
rect 539234 -5734 539854 709670
rect 541794 -1894 542414 705830
rect 542954 -7654 543574 711590
rect 545514 -3814 546134 707750
rect 549234 -5734 549854 709670
rect 551794 -1894 552414 705830
rect 552954 -7654 553574 711590
rect 555514 -3814 556134 707750
rect 559234 -5734 559854 709670
rect 561794 -1894 562414 705830
rect 562954 -7654 563574 711590
rect 565514 -3814 566134 707750
rect 569234 -5734 569854 709670
rect 571794 -1894 572414 705830
rect 572954 -7654 573574 711590
rect 575514 -3814 576134 707750
rect 579234 -5734 579854 709670
rect 581794 -1894 582414 705830
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 54891 3299 55434 640661
rect 56214 635953 59154 640661
rect 59934 635953 61714 640661
rect 62494 635953 62874 640661
rect 63654 635953 65434 640661
rect 66214 635953 69154 640661
rect 69934 635953 71714 640661
rect 72494 635953 72874 640661
rect 73654 635953 75434 640661
rect 76214 635953 79154 640661
rect 79934 635953 81714 640661
rect 82494 635953 82874 640661
rect 83654 635953 85434 640661
rect 86214 635953 89154 640661
rect 89934 635953 91714 640661
rect 92494 635953 92874 640661
rect 93654 635953 95434 640661
rect 96214 635953 99154 640661
rect 99934 635953 101714 640661
rect 102494 635953 102874 640661
rect 103654 635953 105434 640661
rect 106214 635953 109154 640661
rect 109934 635953 111714 640661
rect 112494 635953 112874 640661
rect 113654 635953 115434 640661
rect 116214 635953 119154 640661
rect 119934 635953 121714 640661
rect 122494 635953 122874 640661
rect 123654 635953 125434 640661
rect 126214 635953 129154 640661
rect 129934 635953 131714 640661
rect 132494 635953 132874 640661
rect 133654 635953 135434 640661
rect 136214 635953 139154 640661
rect 139934 635953 141714 640661
rect 142494 635953 142874 640661
rect 143654 635953 145434 640661
rect 146214 635953 149154 640661
rect 149934 635953 151714 640661
rect 152494 635953 152874 640661
rect 153654 635953 155434 640661
rect 156214 635953 159154 640661
rect 159934 635953 161714 640661
rect 162494 635953 162874 640661
rect 163654 635953 165434 640661
rect 166214 635953 169154 640661
rect 169934 635953 171714 640661
rect 56214 521080 171714 635953
rect 56214 466228 59154 521080
rect 59934 466228 61714 521080
rect 62494 466228 62874 521080
rect 63654 466228 65434 521080
rect 66214 466228 69154 521080
rect 69934 466228 71714 521080
rect 72494 466228 72874 521080
rect 73654 466228 75434 521080
rect 76214 466228 79154 521080
rect 79934 466228 81714 521080
rect 82494 466228 82874 521080
rect 83654 466228 85434 521080
rect 86214 466228 89154 521080
rect 89934 466228 91714 521080
rect 92494 466228 92874 521080
rect 93654 466228 95434 521080
rect 96214 466228 99154 521080
rect 99934 466228 101714 521080
rect 102494 466228 102874 521080
rect 103654 466228 105434 521080
rect 106214 466228 109154 521080
rect 109934 466228 111714 521080
rect 112494 466228 112874 521080
rect 113654 466228 115434 521080
rect 116214 466228 119154 521080
rect 119934 466228 121714 521080
rect 122494 466228 122874 521080
rect 123654 466228 125434 521080
rect 126214 466228 129154 521080
rect 129934 466228 131714 521080
rect 132494 466228 132874 521080
rect 133654 466228 135434 521080
rect 136214 466228 139154 521080
rect 139934 466228 141714 521080
rect 142494 466228 142874 521080
rect 143654 466228 145434 521080
rect 146214 466228 149154 521080
rect 149934 466228 151714 521080
rect 152494 466228 152874 521080
rect 153654 466228 155434 521080
rect 156214 466228 159154 521080
rect 159934 466228 161714 521080
rect 162494 466228 162874 521080
rect 163654 466228 165434 521080
rect 166214 466228 169154 521080
rect 169934 466228 171714 521080
rect 172494 466228 172874 640661
rect 173654 466228 175434 640661
rect 176214 466228 179154 640661
rect 179934 466228 181714 640661
rect 182494 466228 182874 640661
rect 183654 466228 185434 640661
rect 186214 466228 189154 640661
rect 189934 466228 191714 640661
rect 192494 466228 192874 640661
rect 193654 466228 195434 640661
rect 196214 491080 322874 640661
rect 196214 466228 199154 491080
rect 56214 379080 199154 466228
rect 56214 359228 59154 379080
rect 59934 359228 61714 379080
rect 62494 359228 62874 379080
rect 63654 359228 65434 379080
rect 66214 359228 69154 379080
rect 69934 359228 71714 379080
rect 72494 359228 72874 379080
rect 73654 359228 75434 379080
rect 76214 359228 79154 379080
rect 79934 359228 81714 379080
rect 82494 359228 82874 379080
rect 83654 359228 85434 379080
rect 86214 359228 89154 379080
rect 89934 359228 91714 379080
rect 92494 359228 92874 379080
rect 93654 359228 95434 379080
rect 96214 359228 99154 379080
rect 99934 359228 101714 379080
rect 102494 359228 102874 379080
rect 103654 359228 105434 379080
rect 106214 359228 109154 379080
rect 109934 359228 111714 379080
rect 112494 359228 112874 379080
rect 113654 359228 115434 379080
rect 116214 359228 119154 379080
rect 119934 359228 121714 379080
rect 122494 359228 122874 379080
rect 123654 359228 125434 379080
rect 126214 359228 129154 379080
rect 129934 359228 131714 379080
rect 132494 359228 132874 379080
rect 133654 359228 135434 379080
rect 136214 359228 139154 379080
rect 139934 359228 141714 379080
rect 142494 359228 142874 379080
rect 143654 359228 145434 379080
rect 146214 359228 149154 379080
rect 149934 359228 151714 379080
rect 152494 359228 152874 379080
rect 153654 359228 155434 379080
rect 156214 359228 159154 379080
rect 159934 359228 161714 379080
rect 162494 359228 162874 379080
rect 163654 359228 165434 379080
rect 166214 359228 169154 379080
rect 169934 359228 171714 379080
rect 172494 359228 172874 379080
rect 173654 359228 175434 379080
rect 176214 359228 179154 379080
rect 179934 359228 181714 379080
rect 182494 359228 182874 379080
rect 183654 359228 185434 379080
rect 186214 359228 189154 379080
rect 189934 359228 191714 379080
rect 192494 359228 192874 379080
rect 193654 359228 195434 379080
rect 196214 359228 199154 379080
rect 56214 272080 199154 359228
rect 56214 252228 59154 272080
rect 59934 252228 61714 272080
rect 62494 252228 62874 272080
rect 63654 252228 65434 272080
rect 66214 252228 69154 272080
rect 69934 252228 71714 272080
rect 72494 252228 72874 272080
rect 73654 252228 75434 272080
rect 76214 252228 79154 272080
rect 79934 252228 81714 272080
rect 82494 252228 82874 272080
rect 83654 252228 85434 272080
rect 86214 252228 89154 272080
rect 89934 252228 91714 272080
rect 92494 252228 92874 272080
rect 93654 252228 95434 272080
rect 96214 252228 99154 272080
rect 99934 252228 101714 272080
rect 102494 252228 102874 272080
rect 103654 252228 105434 272080
rect 106214 252228 109154 272080
rect 109934 252228 111714 272080
rect 112494 252228 112874 272080
rect 113654 252228 115434 272080
rect 116214 252228 119154 272080
rect 119934 252228 121714 272080
rect 122494 252228 122874 272080
rect 123654 252228 125434 272080
rect 126214 252228 129154 272080
rect 129934 252228 131714 272080
rect 132494 252228 132874 272080
rect 133654 252228 135434 272080
rect 136214 252228 139154 272080
rect 139934 252228 141714 272080
rect 142494 252228 142874 272080
rect 143654 252228 145434 272080
rect 146214 252228 149154 272080
rect 149934 252228 151714 272080
rect 152494 252228 152874 272080
rect 153654 252228 155434 272080
rect 156214 252228 159154 272080
rect 159934 252228 161714 272080
rect 162494 252228 162874 272080
rect 163654 252228 165434 272080
rect 166214 252228 169154 272080
rect 169934 252228 171714 272080
rect 172494 252228 172874 272080
rect 173654 252228 175434 272080
rect 176214 252228 179154 272080
rect 179934 252228 181714 272080
rect 182494 252228 182874 272080
rect 183654 252228 185434 272080
rect 186214 252228 189154 272080
rect 189934 252228 191714 272080
rect 192494 252228 192874 272080
rect 193654 252228 195434 272080
rect 196214 252228 199154 272080
rect 56214 165080 199154 252228
rect 56214 145228 59154 165080
rect 59934 145228 61714 165080
rect 62494 145228 62874 165080
rect 63654 145228 65434 165080
rect 66214 145228 69154 165080
rect 69934 145228 71714 165080
rect 72494 145228 72874 165080
rect 73654 145228 75434 165080
rect 76214 145228 79154 165080
rect 79934 145228 81714 165080
rect 82494 145228 82874 165080
rect 83654 145228 85434 165080
rect 86214 145228 89154 165080
rect 89934 145228 91714 165080
rect 92494 145228 92874 165080
rect 93654 145228 95434 165080
rect 96214 145228 99154 165080
rect 99934 145228 101714 165080
rect 102494 145228 102874 165080
rect 103654 145228 105434 165080
rect 106214 145228 109154 165080
rect 109934 145228 111714 165080
rect 112494 145228 112874 165080
rect 113654 145228 115434 165080
rect 116214 145228 119154 165080
rect 119934 145228 121714 165080
rect 122494 145228 122874 165080
rect 123654 145228 125434 165080
rect 126214 145228 129154 165080
rect 129934 145228 131714 165080
rect 132494 145228 132874 165080
rect 133654 145228 135434 165080
rect 136214 145228 139154 165080
rect 139934 145228 141714 165080
rect 142494 145228 142874 165080
rect 143654 145228 145434 165080
rect 146214 145228 149154 165080
rect 149934 145228 151714 165080
rect 152494 145228 152874 165080
rect 153654 145228 155434 165080
rect 156214 145228 159154 165080
rect 159934 145228 161714 165080
rect 162494 145228 162874 165080
rect 163654 145228 165434 165080
rect 166214 145228 169154 165080
rect 169934 145228 171714 165080
rect 172494 145228 172874 165080
rect 173654 145228 175434 165080
rect 176214 145228 179154 165080
rect 179934 145228 181714 165080
rect 182494 145228 182874 165080
rect 183654 145228 185434 165080
rect 186214 145228 189154 165080
rect 189934 145228 191714 165080
rect 192494 145228 192874 165080
rect 193654 145228 195434 165080
rect 196214 145228 199154 165080
rect 56214 58080 199154 145228
rect 56214 3299 59154 58080
rect 59934 3299 61714 58080
rect 62494 3299 62874 58080
rect 63654 3299 65434 58080
rect 66214 3299 69154 58080
rect 69934 3299 71714 58080
rect 72494 3299 72874 58080
rect 73654 3299 75434 58080
rect 76214 3299 79154 58080
rect 79934 3299 81714 58080
rect 82494 3299 82874 58080
rect 83654 3299 85434 58080
rect 86214 3299 89154 58080
rect 89934 3299 91714 58080
rect 92494 3299 92874 58080
rect 93654 3299 95434 58080
rect 96214 3299 99154 58080
rect 99934 3299 101714 58080
rect 102494 3299 102874 58080
rect 103654 3299 105434 58080
rect 106214 3299 109154 58080
rect 109934 3299 111714 58080
rect 112494 3299 112874 58080
rect 113654 3299 115434 58080
rect 116214 3299 119154 58080
rect 119934 3299 121714 58080
rect 122494 3299 122874 58080
rect 123654 3299 125434 58080
rect 126214 3299 129154 58080
rect 129934 3299 131714 58080
rect 132494 3299 132874 58080
rect 133654 3299 135434 58080
rect 136214 3299 139154 58080
rect 139934 3299 141714 58080
rect 142494 3299 142874 58080
rect 143654 3299 145434 58080
rect 146214 3299 149154 58080
rect 149934 3299 151714 58080
rect 152494 3299 152874 58080
rect 153654 3299 155434 58080
rect 156214 3299 159154 58080
rect 159934 3299 161714 58080
rect 162494 3299 162874 58080
rect 163654 3299 165434 58080
rect 166214 3299 169154 58080
rect 169934 3299 171714 58080
rect 172494 3299 172874 58080
rect 173654 3299 175434 58080
rect 176214 3299 179154 58080
rect 179934 3299 181714 58080
rect 182494 3299 182874 58080
rect 183654 3299 185434 58080
rect 186214 3299 189154 58080
rect 189934 3299 191714 58080
rect 192494 3299 192874 58080
rect 193654 3299 195434 58080
rect 196214 3299 199154 58080
rect 199934 3299 201714 491080
rect 202494 3299 202874 491080
rect 203654 3299 205434 491080
rect 206214 3299 209154 491080
rect 209934 3299 211714 491080
rect 212494 3299 212874 491080
rect 213654 3299 215434 491080
rect 216214 466228 219154 491080
rect 219934 466228 221714 491080
rect 222494 466228 222874 491080
rect 223654 466228 225434 491080
rect 226214 466228 229154 491080
rect 229934 466228 231714 491080
rect 232494 466228 232874 491080
rect 233654 466228 235434 491080
rect 236214 466228 239154 491080
rect 239934 466228 241714 491080
rect 242494 466228 242874 491080
rect 243654 466228 245434 491080
rect 246214 466228 249154 491080
rect 249934 466228 251714 491080
rect 252494 466228 252874 491080
rect 253654 466228 255434 491080
rect 256214 466228 259154 491080
rect 259934 466228 261714 491080
rect 262494 466228 262874 491080
rect 263654 466228 265434 491080
rect 266214 466228 269154 491080
rect 269934 466228 271714 491080
rect 272494 466228 272874 491080
rect 273654 466228 275434 491080
rect 276214 466228 279154 491080
rect 279934 466228 281714 491080
rect 282494 466228 282874 491080
rect 283654 466228 285434 491080
rect 286214 466228 289154 491080
rect 289934 466228 291714 491080
rect 292494 466228 292874 491080
rect 293654 466228 295434 491080
rect 296214 466228 299154 491080
rect 299934 466228 301714 491080
rect 302494 466228 302874 491080
rect 303654 466228 305434 491080
rect 306214 466228 309154 491080
rect 309934 466228 311714 491080
rect 312494 466228 312874 491080
rect 313654 466228 315434 491080
rect 316214 466228 319154 491080
rect 319934 466228 321714 491080
rect 322494 466228 322874 491080
rect 323654 466228 325434 640661
rect 326214 466228 329154 640661
rect 329934 466228 331714 640661
rect 332494 466228 332874 640661
rect 333654 466228 335434 640661
rect 336214 466228 339154 640661
rect 339934 466228 341714 640661
rect 342494 466228 342874 640661
rect 343654 466228 345434 640661
rect 346214 466228 349154 640661
rect 349934 466228 351714 640661
rect 352494 578080 419154 640661
rect 352494 558019 352874 578080
rect 353654 558019 355434 578080
rect 356214 558019 359154 578080
rect 359934 558019 361714 578080
rect 362494 558019 362874 578080
rect 363654 558019 365434 578080
rect 366214 558019 369154 578080
rect 369934 558019 371714 578080
rect 372494 558019 372874 578080
rect 373654 558019 375434 578080
rect 376214 558019 379154 578080
rect 379934 558019 381714 578080
rect 382494 558019 382874 578080
rect 383654 558019 385434 578080
rect 386214 558019 389154 578080
rect 389934 558019 391714 578080
rect 392494 558019 392874 578080
rect 393654 558019 395434 578080
rect 396214 558019 399154 578080
rect 399934 558019 401714 578080
rect 402494 558019 402874 578080
rect 403654 558019 405434 578080
rect 406214 558019 409154 578080
rect 409934 558019 411714 578080
rect 412494 558019 412874 578080
rect 413654 558019 415434 578080
rect 416214 558019 419154 578080
rect 352494 491080 419154 558019
rect 352494 466228 352874 491080
rect 353654 466228 355434 491080
rect 356214 466228 359154 491080
rect 216214 379080 359154 466228
rect 216214 359228 219154 379080
rect 219934 359228 221714 379080
rect 222494 359228 222874 379080
rect 223654 359228 225434 379080
rect 226214 359228 229154 379080
rect 229934 359228 231714 379080
rect 232494 359228 232874 379080
rect 233654 359228 235434 379080
rect 236214 359228 239154 379080
rect 239934 359228 241714 379080
rect 242494 359228 242874 379080
rect 243654 359228 245434 379080
rect 246214 359228 249154 379080
rect 249934 359228 251714 379080
rect 252494 359228 252874 379080
rect 253654 359228 255434 379080
rect 256214 359228 259154 379080
rect 259934 359228 261714 379080
rect 262494 359228 262874 379080
rect 263654 359228 265434 379080
rect 266214 359228 269154 379080
rect 269934 359228 271714 379080
rect 272494 359228 272874 379080
rect 273654 359228 275434 379080
rect 276214 359228 279154 379080
rect 279934 359228 281714 379080
rect 282494 359228 282874 379080
rect 283654 359228 285434 379080
rect 286214 359228 289154 379080
rect 289934 359228 291714 379080
rect 292494 359228 292874 379080
rect 293654 359228 295434 379080
rect 296214 359228 299154 379080
rect 299934 359228 301714 379080
rect 302494 359228 302874 379080
rect 303654 359228 305434 379080
rect 306214 359228 309154 379080
rect 309934 359228 311714 379080
rect 312494 359228 312874 379080
rect 313654 359228 315434 379080
rect 316214 359228 319154 379080
rect 319934 359228 321714 379080
rect 322494 359228 322874 379080
rect 323654 359228 325434 379080
rect 326214 359228 329154 379080
rect 329934 359228 331714 379080
rect 332494 359228 332874 379080
rect 333654 359228 335434 379080
rect 336214 359228 339154 379080
rect 339934 359228 341714 379080
rect 342494 359228 342874 379080
rect 343654 359228 345434 379080
rect 346214 359228 349154 379080
rect 349934 359228 351714 379080
rect 352494 359228 352874 379080
rect 353654 359228 355434 379080
rect 356214 359228 359154 379080
rect 216214 272080 359154 359228
rect 216214 252228 219154 272080
rect 219934 252228 221714 272080
rect 222494 252228 222874 272080
rect 223654 252228 225434 272080
rect 226214 252228 229154 272080
rect 229934 252228 231714 272080
rect 232494 252228 232874 272080
rect 233654 252228 235434 272080
rect 236214 252228 239154 272080
rect 239934 252228 241714 272080
rect 242494 252228 242874 272080
rect 243654 252228 245434 272080
rect 246214 252228 249154 272080
rect 249934 252228 251714 272080
rect 252494 252228 252874 272080
rect 253654 252228 255434 272080
rect 256214 252228 259154 272080
rect 259934 252228 261714 272080
rect 262494 252228 262874 272080
rect 263654 252228 265434 272080
rect 266214 252228 269154 272080
rect 269934 252228 271714 272080
rect 272494 252228 272874 272080
rect 273654 252228 275434 272080
rect 276214 252228 279154 272080
rect 279934 252228 281714 272080
rect 282494 252228 282874 272080
rect 283654 252228 285434 272080
rect 286214 252228 289154 272080
rect 289934 252228 291714 272080
rect 292494 252228 292874 272080
rect 293654 252228 295434 272080
rect 296214 252228 299154 272080
rect 299934 252228 301714 272080
rect 302494 252228 302874 272080
rect 303654 252228 305434 272080
rect 306214 252228 309154 272080
rect 309934 252228 311714 272080
rect 312494 252228 312874 272080
rect 313654 252228 315434 272080
rect 316214 252228 319154 272080
rect 319934 252228 321714 272080
rect 322494 252228 322874 272080
rect 323654 252228 325434 272080
rect 326214 252228 329154 272080
rect 329934 252228 331714 272080
rect 332494 252228 332874 272080
rect 333654 252228 335434 272080
rect 336214 252228 339154 272080
rect 339934 252228 341714 272080
rect 342494 252228 342874 272080
rect 343654 252228 345434 272080
rect 346214 252228 349154 272080
rect 349934 252228 351714 272080
rect 352494 252228 352874 272080
rect 353654 252228 355434 272080
rect 356214 252228 359154 272080
rect 216214 165080 359154 252228
rect 216214 145228 219154 165080
rect 219934 145228 221714 165080
rect 222494 145228 222874 165080
rect 223654 145228 225434 165080
rect 226214 145228 229154 165080
rect 229934 145228 231714 165080
rect 232494 145228 232874 165080
rect 233654 145228 235434 165080
rect 236214 145228 239154 165080
rect 239934 145228 241714 165080
rect 242494 145228 242874 165080
rect 243654 145228 245434 165080
rect 246214 145228 249154 165080
rect 249934 145228 251714 165080
rect 252494 145228 252874 165080
rect 253654 145228 255434 165080
rect 256214 145228 259154 165080
rect 259934 145228 261714 165080
rect 262494 145228 262874 165080
rect 263654 145228 265434 165080
rect 266214 145228 269154 165080
rect 269934 145228 271714 165080
rect 272494 145228 272874 165080
rect 273654 145228 275434 165080
rect 276214 145228 279154 165080
rect 279934 145228 281714 165080
rect 282494 145228 282874 165080
rect 283654 145228 285434 165080
rect 286214 145228 289154 165080
rect 289934 145228 291714 165080
rect 292494 145228 292874 165080
rect 293654 145228 295434 165080
rect 296214 145228 299154 165080
rect 299934 145228 301714 165080
rect 302494 145228 302874 165080
rect 303654 145228 305434 165080
rect 306214 145228 309154 165080
rect 309934 145228 311714 165080
rect 312494 145228 312874 165080
rect 313654 145228 315434 165080
rect 316214 145228 319154 165080
rect 319934 145228 321714 165080
rect 322494 145228 322874 165080
rect 323654 145228 325434 165080
rect 326214 145228 329154 165080
rect 329934 145228 331714 165080
rect 332494 145228 332874 165080
rect 333654 145228 335434 165080
rect 336214 145228 339154 165080
rect 339934 145228 341714 165080
rect 342494 145228 342874 165080
rect 343654 145228 345434 165080
rect 346214 145228 349154 165080
rect 349934 145228 351714 165080
rect 352494 145228 352874 165080
rect 353654 145228 355434 165080
rect 356214 145228 359154 165080
rect 216214 58080 359154 145228
rect 216214 3299 219154 58080
rect 219934 3299 221714 58080
rect 222494 3299 222874 58080
rect 223654 3299 225434 58080
rect 226214 3299 229154 58080
rect 229934 3299 231714 58080
rect 232494 3299 232874 58080
rect 233654 3299 235434 58080
rect 236214 3299 239154 58080
rect 239934 3299 241714 58080
rect 242494 3299 242874 58080
rect 243654 3299 245434 58080
rect 246214 3299 249154 58080
rect 249934 3299 251714 58080
rect 252494 3299 252874 58080
rect 253654 3299 255434 58080
rect 256214 3299 259154 58080
rect 259934 3299 261714 58080
rect 262494 3299 262874 58080
rect 263654 3299 265434 58080
rect 266214 3299 269154 58080
rect 269934 3299 271714 58080
rect 272494 3299 272874 58080
rect 273654 3299 275434 58080
rect 276214 3299 279154 58080
rect 279934 3299 281714 58080
rect 282494 3299 282874 58080
rect 283654 3299 285434 58080
rect 286214 3299 289154 58080
rect 289934 3299 291714 58080
rect 292494 3299 292874 58080
rect 293654 3299 295434 58080
rect 296214 3299 299154 58080
rect 299934 3299 301714 58080
rect 302494 3299 302874 58080
rect 303654 3299 305434 58080
rect 306214 3299 309154 58080
rect 309934 3299 311714 58080
rect 312494 3299 312874 58080
rect 313654 3299 315434 58080
rect 316214 3299 319154 58080
rect 319934 3299 321714 58080
rect 322494 3299 322874 58080
rect 323654 3299 325434 58080
rect 326214 3299 329154 58080
rect 329934 3299 331714 58080
rect 332494 3299 332874 58080
rect 333654 3299 335434 58080
rect 336214 3299 339154 58080
rect 339934 3299 341714 58080
rect 342494 3299 342874 58080
rect 343654 3299 345434 58080
rect 346214 3299 349154 58080
rect 349934 3299 351714 58080
rect 352494 3299 352874 58080
rect 353654 3299 355434 58080
rect 356214 3299 359154 58080
rect 359934 3299 361714 491080
rect 362494 3299 362874 491080
rect 363654 3299 365434 491080
rect 366214 3299 369154 491080
rect 369934 3299 371714 491080
rect 372494 3299 372874 491080
rect 373654 3299 375434 491080
rect 376214 466228 379154 491080
rect 379934 466228 381714 491080
rect 382494 466228 382874 491080
rect 383654 466228 385434 491080
rect 386214 466228 389154 491080
rect 389934 466228 391714 491080
rect 392494 466228 392874 491080
rect 393654 466228 395434 491080
rect 396214 466228 399154 491080
rect 399934 466228 401714 491080
rect 402494 466228 402874 491080
rect 403654 466228 405434 491080
rect 406214 466228 409154 491080
rect 409934 466228 411714 491080
rect 412494 466228 412874 491080
rect 413654 466228 415434 491080
rect 416214 466228 419154 491080
rect 419934 466228 421714 640661
rect 422494 466228 422874 640661
rect 423654 466228 425434 640661
rect 426214 466228 429154 640661
rect 429934 466228 431714 640661
rect 432494 466228 432874 640661
rect 433654 466228 435434 640661
rect 436214 466228 439154 640661
rect 439934 466228 441714 640661
rect 442494 466228 442874 640661
rect 443654 466228 445434 640661
rect 446214 578080 515434 640661
rect 446214 554920 449154 578080
rect 449934 554920 451714 578080
rect 452494 554920 452874 578080
rect 453654 554920 455434 578080
rect 456214 554920 459154 578080
rect 459934 554920 461714 578080
rect 462494 554920 462874 578080
rect 463654 554920 465434 578080
rect 466214 554920 469154 578080
rect 469934 554920 471714 578080
rect 472494 554920 472874 578080
rect 473654 554920 475434 578080
rect 476214 554920 479154 578080
rect 479934 554920 481714 578080
rect 482494 554920 482874 578080
rect 483654 554920 485434 578080
rect 486214 554920 489154 578080
rect 489934 554920 491714 578080
rect 492494 554920 492874 578080
rect 493654 554920 495434 578080
rect 496214 554920 499154 578080
rect 499934 554920 501714 578080
rect 502494 554920 502874 578080
rect 446214 501080 502874 554920
rect 446214 466228 449154 501080
rect 449934 466228 451714 501080
rect 452494 466228 452874 501080
rect 453654 466228 455434 501080
rect 456214 466228 459154 501080
rect 459934 466228 461714 501080
rect 462494 466228 462874 501080
rect 463654 466228 465434 501080
rect 466214 466228 469154 501080
rect 469934 466228 471714 501080
rect 472494 466228 472874 501080
rect 473654 466228 475434 501080
rect 476214 466228 479154 501080
rect 479934 466228 481714 501080
rect 482494 466228 482874 501080
rect 483654 466228 485434 501080
rect 486214 466228 489154 501080
rect 489934 466228 491714 501080
rect 492494 466228 492874 501080
rect 493654 466228 495434 501080
rect 496214 466228 499154 501080
rect 499934 466228 501714 501080
rect 502494 466228 502874 501080
rect 503654 466228 505434 578080
rect 506214 466228 509154 578080
rect 509934 466228 511714 578080
rect 512494 466228 512874 578080
rect 513654 466228 515434 578080
rect 516214 466228 517533 640661
rect 376214 379080 517533 466228
rect 376214 359228 379154 379080
rect 379934 359228 381714 379080
rect 382494 359228 382874 379080
rect 383654 359228 385434 379080
rect 386214 359228 389154 379080
rect 389934 359228 391714 379080
rect 392494 359228 392874 379080
rect 393654 359228 395434 379080
rect 396214 359228 399154 379080
rect 399934 359228 401714 379080
rect 402494 359228 402874 379080
rect 403654 359228 405434 379080
rect 406214 359228 409154 379080
rect 409934 359228 411714 379080
rect 412494 359228 412874 379080
rect 413654 359228 415434 379080
rect 416214 359228 419154 379080
rect 419934 359228 421714 379080
rect 422494 359228 422874 379080
rect 423654 359228 425434 379080
rect 426214 359228 429154 379080
rect 429934 359228 431714 379080
rect 432494 359228 432874 379080
rect 433654 359228 435434 379080
rect 436214 359228 439154 379080
rect 439934 359228 441714 379080
rect 442494 359228 442874 379080
rect 443654 359228 445434 379080
rect 446214 359228 449154 379080
rect 449934 359228 451714 379080
rect 452494 359228 452874 379080
rect 453654 359228 455434 379080
rect 456214 359228 459154 379080
rect 459934 359228 461714 379080
rect 462494 359228 462874 379080
rect 463654 359228 465434 379080
rect 466214 359228 469154 379080
rect 469934 359228 471714 379080
rect 472494 359228 472874 379080
rect 473654 359228 475434 379080
rect 476214 359228 479154 379080
rect 479934 359228 481714 379080
rect 482494 359228 482874 379080
rect 483654 359228 485434 379080
rect 486214 359228 489154 379080
rect 489934 359228 491714 379080
rect 492494 359228 492874 379080
rect 493654 359228 495434 379080
rect 496214 359228 499154 379080
rect 499934 359228 501714 379080
rect 502494 359228 502874 379080
rect 503654 359228 505434 379080
rect 506214 359228 509154 379080
rect 509934 359228 511714 379080
rect 512494 359228 512874 379080
rect 513654 359228 515434 379080
rect 516214 359228 517533 379080
rect 376214 272080 517533 359228
rect 376214 252228 379154 272080
rect 379934 252228 381714 272080
rect 382494 252228 382874 272080
rect 383654 252228 385434 272080
rect 386214 252228 389154 272080
rect 389934 252228 391714 272080
rect 392494 252228 392874 272080
rect 393654 252228 395434 272080
rect 396214 252228 399154 272080
rect 399934 252228 401714 272080
rect 402494 252228 402874 272080
rect 403654 252228 405434 272080
rect 406214 252228 409154 272080
rect 409934 252228 411714 272080
rect 412494 252228 412874 272080
rect 413654 252228 415434 272080
rect 416214 252228 419154 272080
rect 419934 252228 421714 272080
rect 422494 252228 422874 272080
rect 423654 252228 425434 272080
rect 426214 252228 429154 272080
rect 429934 252228 431714 272080
rect 432494 252228 432874 272080
rect 433654 252228 435434 272080
rect 436214 252228 439154 272080
rect 439934 252228 441714 272080
rect 442494 252228 442874 272080
rect 443654 252228 445434 272080
rect 446214 252228 449154 272080
rect 449934 252228 451714 272080
rect 452494 252228 452874 272080
rect 453654 252228 455434 272080
rect 456214 252228 459154 272080
rect 459934 252228 461714 272080
rect 462494 252228 462874 272080
rect 463654 252228 465434 272080
rect 466214 252228 469154 272080
rect 469934 252228 471714 272080
rect 472494 252228 472874 272080
rect 473654 252228 475434 272080
rect 476214 252228 479154 272080
rect 479934 252228 481714 272080
rect 482494 252228 482874 272080
rect 483654 252228 485434 272080
rect 486214 252228 489154 272080
rect 489934 252228 491714 272080
rect 492494 252228 492874 272080
rect 493654 252228 495434 272080
rect 496214 252228 499154 272080
rect 499934 252228 501714 272080
rect 502494 252228 502874 272080
rect 503654 252228 505434 272080
rect 506214 252228 509154 272080
rect 509934 252228 511714 272080
rect 512494 252228 512874 272080
rect 513654 252228 515434 272080
rect 516214 252228 517533 272080
rect 376214 165080 517533 252228
rect 376214 145228 379154 165080
rect 379934 145228 381714 165080
rect 382494 145228 382874 165080
rect 383654 145228 385434 165080
rect 386214 145228 389154 165080
rect 389934 145228 391714 165080
rect 392494 145228 392874 165080
rect 393654 145228 395434 165080
rect 396214 145228 399154 165080
rect 399934 145228 401714 165080
rect 402494 145228 402874 165080
rect 403654 145228 405434 165080
rect 406214 145228 409154 165080
rect 409934 145228 411714 165080
rect 412494 145228 412874 165080
rect 413654 145228 415434 165080
rect 416214 145228 419154 165080
rect 419934 145228 421714 165080
rect 422494 145228 422874 165080
rect 423654 145228 425434 165080
rect 426214 145228 429154 165080
rect 429934 145228 431714 165080
rect 432494 145228 432874 165080
rect 433654 145228 435434 165080
rect 436214 145228 439154 165080
rect 439934 145228 441714 165080
rect 442494 145228 442874 165080
rect 443654 145228 445434 165080
rect 446214 145228 449154 165080
rect 449934 145228 451714 165080
rect 452494 145228 452874 165080
rect 453654 145228 455434 165080
rect 456214 145228 459154 165080
rect 459934 145228 461714 165080
rect 462494 145228 462874 165080
rect 463654 145228 465434 165080
rect 466214 145228 469154 165080
rect 469934 145228 471714 165080
rect 472494 145228 472874 165080
rect 473654 145228 475434 165080
rect 476214 145228 479154 165080
rect 479934 145228 481714 165080
rect 482494 145228 482874 165080
rect 483654 145228 485434 165080
rect 486214 145228 489154 165080
rect 489934 145228 491714 165080
rect 492494 145228 492874 165080
rect 493654 145228 495434 165080
rect 496214 145228 499154 165080
rect 499934 145228 501714 165080
rect 502494 145228 502874 165080
rect 503654 145228 505434 165080
rect 506214 145228 509154 165080
rect 509934 145228 511714 165080
rect 512494 145228 512874 165080
rect 513654 145228 515434 165080
rect 516214 145228 517533 165080
rect 376214 58080 517533 145228
rect 376214 3299 379154 58080
rect 379934 3299 381714 58080
rect 382494 3299 382874 58080
rect 383654 3299 385434 58080
rect 386214 3299 389154 58080
rect 389934 3299 391714 58080
rect 392494 3299 392874 58080
rect 393654 3299 395434 58080
rect 396214 3299 399154 58080
rect 399934 3299 401714 58080
rect 402494 3299 402874 58080
rect 403654 3299 405434 58080
rect 406214 3299 409154 58080
rect 409934 3299 411714 58080
rect 412494 3299 412874 58080
rect 413654 3299 415434 58080
rect 416214 3299 419154 58080
rect 419934 3299 421714 58080
rect 422494 3299 422874 58080
rect 423654 3299 425434 58080
rect 426214 3299 429154 58080
rect 429934 3299 431714 58080
rect 432494 3299 432874 58080
rect 433654 3299 435434 58080
rect 436214 3299 439154 58080
rect 439934 3299 441714 58080
rect 442494 3299 442874 58080
rect 443654 3299 445434 58080
rect 446214 3299 449154 58080
rect 449934 3299 451714 58080
rect 452494 3299 452874 58080
rect 453654 3299 455434 58080
rect 456214 3299 459154 58080
rect 459934 3299 461714 58080
rect 462494 3299 462874 58080
rect 463654 3299 465434 58080
rect 466214 3299 469154 58080
rect 469934 3299 471714 58080
rect 472494 3299 472874 58080
rect 473654 3299 475434 58080
rect 476214 3299 479154 58080
rect 479934 3299 481714 58080
rect 482494 3299 482874 58080
rect 483654 3299 485434 58080
rect 486214 3299 489154 58080
rect 489934 3299 491714 58080
rect 492494 3299 492874 58080
rect 493654 3299 495434 58080
rect 496214 3299 499154 58080
rect 499934 3299 501714 58080
rect 502494 3299 502874 58080
rect 503654 3299 505434 58080
rect 506214 3299 509154 58080
rect 509934 3299 511714 58080
rect 512494 3299 512874 58080
rect 513654 3299 515434 58080
rect 516214 3299 517533 58080
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -6806 700306 590730 700926
rect -4886 696586 588810 697206
rect -8726 694026 592650 694646
rect -2966 692866 586890 693486
rect -6806 690306 590730 690926
rect -4886 686586 588810 687206
rect -8726 684026 592650 684646
rect -2966 682866 586890 683486
rect -6806 680306 590730 680926
rect -4886 676586 588810 677206
rect -8726 674026 592650 674646
rect -2966 672866 586890 673486
rect -6806 670306 590730 670926
rect -4886 666586 588810 667206
rect -8726 664026 592650 664646
rect -2966 662866 586890 663486
rect -6806 660306 590730 660926
rect -4886 656586 588810 657206
rect -8726 654026 592650 654646
rect -2966 652866 586890 653486
rect -6806 650306 590730 650926
rect -4886 646586 588810 647206
rect -8726 644026 592650 644646
rect -2966 642866 586890 643486
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -8726 634026 592650 634646
rect -2966 632866 586890 633486
rect -6806 630306 590730 630926
rect -4886 626586 588810 627206
rect -8726 624026 592650 624646
rect -2966 622866 586890 623486
rect -6806 620306 590730 620926
rect -4886 616586 588810 617206
rect -8726 614026 592650 614646
rect -2966 612866 586890 613486
rect -6806 610306 590730 610926
rect -4886 606586 588810 607206
rect -8726 604026 592650 604646
rect -2966 602866 586890 603486
rect -6806 600306 590730 600926
rect -4886 596586 588810 597206
rect -8726 594026 592650 594646
rect -2966 592866 586890 593486
rect -6806 590306 590730 590926
rect -4886 586586 588810 587206
rect -8726 584026 592650 584646
rect -2966 582866 586890 583486
rect -6806 580306 590730 580926
rect -4886 576586 588810 577206
rect -8726 574026 592650 574646
rect -2966 572866 586890 573486
rect -6806 570306 590730 570926
rect -4886 566586 588810 567206
rect -8726 564026 592650 564646
rect -2966 562866 586890 563486
rect -6806 560306 590730 560926
rect -4886 556586 588810 557206
rect -8726 554026 592650 554646
rect -2966 552866 586890 553486
rect -6806 550306 590730 550926
rect -4886 546586 588810 547206
rect -8726 544026 592650 544646
rect -2966 542866 586890 543486
rect -6806 540306 590730 540926
rect -4886 536586 588810 537206
rect -8726 534026 592650 534646
rect -2966 532866 586890 533486
rect -6806 530306 590730 530926
rect -4886 526586 588810 527206
rect -8726 524026 592650 524646
rect -2966 522866 586890 523486
rect -6806 520306 590730 520926
rect -4886 516586 588810 517206
rect -8726 514026 592650 514646
rect -2966 512866 586890 513486
rect -6806 510306 590730 510926
rect -4886 506586 588810 507206
rect -8726 504026 592650 504646
rect -2966 502866 586890 503486
rect -6806 500306 590730 500926
rect -4886 496586 588810 497206
rect -8726 494026 592650 494646
rect -2966 492866 586890 493486
rect -6806 490306 590730 490926
rect -4886 486586 588810 487206
rect -8726 484026 592650 484646
rect -2966 482866 586890 483486
rect -6806 480306 590730 480926
rect -4886 476586 588810 477206
rect -8726 474026 592650 474646
rect -2966 472866 586890 473486
rect -6806 470306 590730 470926
rect -4886 466586 588810 467206
rect -8726 464026 592650 464646
rect -2966 462866 586890 463486
rect -6806 460306 590730 460926
rect -4886 456586 588810 457206
rect -8726 454026 592650 454646
rect -2966 452866 586890 453486
rect -6806 450306 590730 450926
rect -4886 446586 588810 447206
rect -8726 444026 592650 444646
rect -2966 442866 586890 443486
rect -6806 440306 590730 440926
rect -4886 436586 588810 437206
rect -8726 434026 592650 434646
rect -2966 432866 586890 433486
rect -6806 430306 590730 430926
rect -4886 426586 588810 427206
rect -8726 424026 592650 424646
rect -2966 422866 586890 423486
rect -6806 420306 590730 420926
rect -4886 416586 588810 417206
rect -8726 414026 592650 414646
rect -2966 412866 586890 413486
rect -6806 410306 590730 410926
rect -4886 406586 588810 407206
rect -8726 404026 592650 404646
rect -2966 402866 586890 403486
rect -6806 400306 590730 400926
rect -4886 396586 588810 397206
rect -8726 394026 592650 394646
rect -2966 392866 586890 393486
rect -6806 390306 590730 390926
rect -4886 386586 588810 387206
rect -8726 384026 592650 384646
rect -2966 382866 586890 383486
rect -6806 380306 590730 380926
rect -4886 376586 588810 377206
rect -8726 374026 592650 374646
rect -2966 372866 586890 373486
rect -6806 370306 590730 370926
rect -4886 366586 588810 367206
rect -8726 364026 592650 364646
rect -2966 362866 586890 363486
rect -6806 360306 590730 360926
rect -4886 356586 588810 357206
rect -8726 354026 592650 354646
rect -2966 352866 586890 353486
rect -6806 350306 590730 350926
rect -4886 346586 588810 347206
rect -8726 344026 592650 344646
rect -2966 342866 586890 343486
rect -6806 340306 590730 340926
rect -4886 336586 588810 337206
rect -8726 334026 592650 334646
rect -2966 332866 586890 333486
rect -6806 330306 590730 330926
rect -4886 326586 588810 327206
rect -8726 324026 592650 324646
rect -2966 322866 586890 323486
rect -6806 320306 590730 320926
rect -4886 316586 588810 317206
rect -8726 314026 592650 314646
rect -2966 312866 586890 313486
rect -6806 310306 590730 310926
rect -4886 306586 588810 307206
rect -8726 304026 592650 304646
rect -2966 302866 586890 303486
rect -6806 300306 590730 300926
rect -4886 296586 588810 297206
rect -8726 294026 592650 294646
rect -2966 292866 586890 293486
rect -6806 290306 590730 290926
rect -4886 286586 588810 287206
rect -8726 284026 592650 284646
rect -2966 282866 586890 283486
rect -6806 280306 590730 280926
rect -4886 276586 588810 277206
rect -8726 274026 592650 274646
rect -2966 272866 586890 273486
rect -6806 270306 590730 270926
rect -4886 266586 588810 267206
rect -8726 264026 592650 264646
rect -2966 262866 586890 263486
rect -6806 260306 590730 260926
rect -4886 256586 588810 257206
rect -8726 254026 592650 254646
rect -2966 252866 586890 253486
rect -6806 250306 590730 250926
rect -4886 246586 588810 247206
rect -8726 244026 592650 244646
rect -2966 242866 586890 243486
rect -6806 240306 590730 240926
rect -4886 236586 588810 237206
rect -8726 234026 592650 234646
rect -2966 232866 586890 233486
rect -6806 230306 590730 230926
rect -4886 226586 588810 227206
rect -8726 224026 592650 224646
rect -2966 222866 586890 223486
rect -6806 220306 590730 220926
rect -4886 216586 588810 217206
rect -8726 214026 592650 214646
rect -2966 212866 586890 213486
rect -6806 210306 590730 210926
rect -4886 206586 588810 207206
rect -8726 204026 592650 204646
rect -2966 202866 586890 203486
rect -6806 200306 590730 200926
rect -4886 196586 588810 197206
rect -8726 194026 592650 194646
rect -2966 192866 586890 193486
rect -6806 190306 590730 190926
rect -4886 186586 588810 187206
rect -8726 184026 592650 184646
rect -2966 182866 586890 183486
rect -6806 180306 590730 180926
rect -4886 176586 588810 177206
rect -8726 174026 592650 174646
rect -2966 172866 586890 173486
rect -6806 170306 590730 170926
rect -4886 166586 588810 167206
rect -8726 164026 592650 164646
rect -2966 162866 586890 163486
rect -6806 160306 590730 160926
rect -4886 156586 588810 157206
rect -8726 154026 592650 154646
rect -2966 152866 586890 153486
rect -6806 150306 590730 150926
rect -4886 146586 588810 147206
rect -8726 144026 592650 144646
rect -2966 142866 586890 143486
rect -6806 140306 590730 140926
rect -4886 136586 588810 137206
rect -8726 134026 592650 134646
rect -2966 132866 586890 133486
rect -6806 130306 590730 130926
rect -4886 126586 588810 127206
rect -8726 124026 592650 124646
rect -2966 122866 586890 123486
rect -6806 120306 590730 120926
rect -4886 116586 588810 117206
rect -8726 114026 592650 114646
rect -2966 112866 586890 113486
rect -6806 110306 590730 110926
rect -4886 106586 588810 107206
rect -8726 104026 592650 104646
rect -2966 102866 586890 103486
rect -6806 100306 590730 100926
rect -4886 96586 588810 97206
rect -8726 94026 592650 94646
rect -2966 92866 586890 93486
rect -6806 90306 590730 90926
rect -4886 86586 588810 87206
rect -8726 84026 592650 84646
rect -2966 82866 586890 83486
rect -6806 80306 590730 80926
rect -4886 76586 588810 77206
rect -8726 74026 592650 74646
rect -2966 72866 586890 73486
rect -6806 70306 590730 70926
rect -4886 66586 588810 67206
rect -8726 64026 592650 64646
rect -2966 62866 586890 63486
rect -6806 60306 590730 60926
rect -4886 56586 588810 57206
rect -8726 54026 592650 54646
rect -2966 52866 586890 53486
rect -6806 50306 590730 50926
rect -4886 46586 588810 47206
rect -8726 44026 592650 44646
rect -2966 42866 586890 43486
rect -6806 40306 590730 40926
rect -4886 36586 588810 37206
rect -8726 34026 592650 34646
rect -2966 32866 586890 33486
rect -6806 30306 590730 30926
rect -4886 26586 588810 27206
rect -8726 24026 592650 24646
rect -2966 22866 586890 23486
rect -6806 20306 590730 20926
rect -4886 16586 588810 17206
rect -8726 14026 592650 14646
rect -2966 12866 586890 13486
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 22866 586890 23486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 42866 586890 43486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 62866 586890 63486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 82866 586890 83486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 102866 586890 103486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 122866 586890 123486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 142866 586890 143486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 162866 586890 163486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 202866 586890 203486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 222866 586890 223486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 242866 586890 243486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 262866 586890 263486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 282866 586890 283486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 302866 586890 303486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 322866 586890 323486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 342866 586890 343486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 382866 586890 383486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 402866 586890 403486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 422866 586890 423486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 442866 586890 443486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 462866 586890 463486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 482866 586890 483486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 502866 586890 503486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 522866 586890 523486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 562866 586890 563486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 582866 586890 583486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 602866 586890 603486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 622866 586890 623486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 642866 586890 643486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 662866 586890 663486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 682866 586890 683486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 -1894 62414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 -1894 82414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 -1894 102414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 -1894 122414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 -1894 142414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 -1894 162414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 -1894 222414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 -1894 242414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 -1894 262414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 -1894 282414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 -1894 302414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 -1894 322414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 341794 -1894 342414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 -1894 382414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 -1894 402414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 -1894 422414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 -1894 442414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 -1894 462414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 -1894 482414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 -1894 502414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 145308 62414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 145308 82414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 145308 102414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 145308 122414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 145308 142414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 145308 162414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 145308 182414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 145308 222414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 145308 242414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 145308 262414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 145308 282414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 145308 302414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 145308 322414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 341794 145308 342414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 145308 382414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 145308 402414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 145308 422414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 145308 442414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 145308 462414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 145308 482414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 145308 502414 165000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 252308 62414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 252308 82414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 252308 102414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 252308 122414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 252308 142414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 252308 162414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 252308 182414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 252308 222414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 252308 242414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 252308 262414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 252308 282414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 252308 302414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 252308 322414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 341794 252308 342414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 252308 382414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 252308 402414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 252308 422414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 252308 442414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 252308 462414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 252308 482414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 252308 502414 272000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 359308 62414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 359308 82414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 359308 102414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 359308 122414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 359308 142414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 359308 162414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 359308 182414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 359308 222414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 359308 242414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 359308 262414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 359308 282414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 359308 302414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 359308 322414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 341794 359308 342414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 359308 382414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 359308 402414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 359308 422414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 359308 442414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 359308 462414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 359308 482414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 359308 502414 379000 6 vccd1
port 532 nsew power input
rlabel metal4 s 201794 -1894 202414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 466308 222414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 466308 242414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 466308 262414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 466308 282414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 466308 302414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 466308 322414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 -1894 362414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 466308 382414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 466308 402414 491000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 466308 462414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 466308 482414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 466308 502414 501000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 466308 62414 521000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 466308 82414 521000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 466308 102414 521000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 466308 122414 521000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 466308 142414 521000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 466308 162414 521000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 558099 362414 578000 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 558099 382414 578000 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 558099 402414 578000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 555000 462414 578000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 555000 482414 578000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 555000 502414 578000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 21794 -1894 22414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 41794 -1894 42414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 636033 62414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 636033 82414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 636033 102414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 636033 122414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 636033 142414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 636033 162414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 466308 182414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 201794 642000 202414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 642000 222414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 642000 242414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 642000 262414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 642000 282414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 642000 302414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 642000 322414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 341794 466308 342414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 645099 362414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 645099 382414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 645099 402414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 466308 422414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 466308 442414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 645099 462414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 645099 482414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 645099 502414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 521794 -1894 522414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 561794 -1894 562414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 581794 -1894 582414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 26586 588810 27206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 46586 588810 47206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 66586 588810 67206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 86586 588810 87206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 106586 588810 107206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 126586 588810 127206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 146586 588810 147206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 166586 588810 167206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 206586 588810 207206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 226586 588810 227206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 246586 588810 247206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 266586 588810 267206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 286586 588810 287206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 306586 588810 307206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 326586 588810 327206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 346586 588810 347206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 386586 588810 387206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 406586 588810 407206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 426586 588810 427206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 446586 588810 447206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 466586 588810 467206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 486586 588810 487206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 506586 588810 507206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 526586 588810 527206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 566586 588810 567206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 586586 588810 587206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 606586 588810 607206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 626586 588810 627206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 646586 588810 647206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 666586 588810 667206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 686586 588810 687206 6 vccd2
port 533 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 -3814 66134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 -3814 86134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 -3814 106134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 -3814 126134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 -3814 146134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 -3814 166134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 -3814 226134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 -3814 246134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 -3814 266134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 -3814 286134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 -3814 306134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 -3814 326134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 345514 -3814 346134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 -3814 386134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 -3814 406134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 -3814 426134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 -3814 446134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 -3814 466134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 -3814 486134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 -3814 506134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 145308 66134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 145308 86134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 145308 106134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 145308 126134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 145308 146134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 145308 166134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 145308 186134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 145308 226134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 145308 246134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 145308 266134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 145308 286134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 145308 306134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 145308 326134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 345514 145308 346134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 145308 386134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 145308 406134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 145308 426134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 145308 446134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 145308 466134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 145308 486134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 145308 506134 165000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 252308 66134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 252308 86134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 252308 106134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 252308 126134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 252308 146134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 252308 166134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 252308 186134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 252308 226134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 252308 246134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 252308 266134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 252308 286134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 252308 306134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 252308 326134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 345514 252308 346134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 252308 386134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 252308 406134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 252308 426134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 252308 446134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 252308 466134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 252308 486134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 252308 506134 272000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 359308 66134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 359308 86134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 359308 106134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 359308 126134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 359308 146134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 359308 166134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 359308 186134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 359308 226134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 359308 246134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 359308 266134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 359308 286134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 359308 306134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 359308 326134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 345514 359308 346134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 359308 386134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 359308 406134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 359308 426134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 359308 446134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 359308 466134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 359308 486134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 359308 506134 379000 6 vccd2
port 533 nsew power input
rlabel metal4 s 205514 -3814 206134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 466308 226134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 466308 246134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 466308 266134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 466308 286134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 466308 306134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 -3814 366134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 466308 386134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 466308 406134 491000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 466308 466134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 466308 486134 501000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 466308 66134 521000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 466308 86134 521000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 466308 106134 521000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 466308 126134 521000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 466308 146134 521000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 466308 166134 521000 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 558099 366134 578000 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 558099 386134 578000 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 558099 406134 578000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 555000 466134 578000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 555000 486134 578000 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 466308 506134 578000 6 vccd2
port 533 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 25514 -3814 26134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 45514 -3814 46134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 636033 66134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 636033 86134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 636033 106134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 636033 126134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 636033 146134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 636033 166134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 466308 186134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 205514 642000 206134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 642000 226134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 642000 246134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 642000 266134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 642000 286134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 642000 306134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 466308 326134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 345514 466308 346134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 645099 366134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 645099 386134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 645099 406134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 466308 426134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 466308 446134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 645099 466134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 645099 486134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 645099 506134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 525514 -3814 526134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 565514 -3814 566134 707750 6 vccd2
port 533 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 30306 590730 30926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 50306 590730 50926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 70306 590730 70926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 90306 590730 90926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 110306 590730 110926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 130306 590730 130926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 150306 590730 150926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 170306 590730 170926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 210306 590730 210926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 230306 590730 230926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 250306 590730 250926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 270306 590730 270926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 290306 590730 290926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 310306 590730 310926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 330306 590730 330926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 350306 590730 350926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 390306 590730 390926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 410306 590730 410926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 430306 590730 430926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 450306 590730 450926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 470306 590730 470926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 490306 590730 490926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 510306 590730 510926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 530306 590730 530926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 570306 590730 570926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 590306 590730 590926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 610306 590730 610926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 630306 590730 630926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 650306 590730 650926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 670306 590730 670926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 690306 590730 690926 6 vdda1
port 534 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 -5734 69854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 -5734 89854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 -5734 109854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 -5734 129854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 -5734 149854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 169234 -5734 169854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 -5734 229854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 -5734 249854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 -5734 269854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 -5734 289854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 -5734 309854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 -5734 329854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 349234 -5734 349854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 -5734 389854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 -5734 409854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 -5734 429854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 -5734 449854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 -5734 469854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 -5734 489854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 -5734 509854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 145308 69854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 145308 89854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 145308 109854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 145308 129854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 145308 149854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 169234 145308 169854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 145308 189854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 145308 229854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 145308 249854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 145308 269854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 145308 289854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 145308 309854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 145308 329854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 349234 145308 349854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 145308 389854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 145308 409854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 145308 429854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 145308 449854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 145308 469854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 145308 489854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 145308 509854 165000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 252308 69854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 252308 89854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 252308 109854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 252308 129854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 252308 149854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 169234 252308 169854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 252308 189854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 252308 229854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 252308 249854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 252308 269854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 252308 289854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 252308 309854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 252308 329854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 349234 252308 349854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 252308 389854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 252308 409854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 252308 429854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 252308 449854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 252308 469854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 252308 489854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 252308 509854 272000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 359308 69854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 359308 89854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 359308 109854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 359308 129854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 359308 149854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 169234 359308 169854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 359308 189854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 359308 229854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 359308 249854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 359308 269854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 359308 289854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 359308 309854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 359308 329854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 349234 359308 349854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 359308 389854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 359308 409854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 359308 429854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 359308 449854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 359308 469854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 359308 489854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 359308 509854 379000 6 vdda1
port 534 nsew power input
rlabel metal4 s 209234 -5734 209854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 466308 229854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 466308 249854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 466308 269854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 466308 289854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 466308 309854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 -5734 369854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 466308 389854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 466308 409854 491000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 466308 449854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 466308 469854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 466308 489854 501000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 466308 69854 521000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 466308 89854 521000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 466308 109854 521000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 466308 129854 521000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 466308 149854 521000 6 vdda1
port 534 nsew power input
rlabel metal4 s 169234 466308 169854 521000 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 558099 369854 578000 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 558099 389854 578000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 558099 409854 578000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 555000 449854 578000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 555000 469854 578000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 555000 489854 578000 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 466308 509854 578000 6 vdda1
port 534 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 29234 -5734 29854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 49234 -5734 49854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 636033 69854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 636033 89854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 636033 109854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 636033 129854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 636033 149854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 169234 636033 169854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 466308 189854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 209234 642000 209854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 642000 229854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 642000 249854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 642000 269854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 642000 289854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 642000 309854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 466308 329854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 349234 466308 349854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 645099 369854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 645099 389854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 645099 409854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 466308 429854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 645099 449854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 645099 469854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 645099 489854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 645099 509854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 529234 -5734 529854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 569234 -5734 569854 709670 6 vdda1
port 534 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 34026 592650 34646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 54026 592650 54646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 74026 592650 74646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 94026 592650 94646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 114026 592650 114646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 134026 592650 134646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 154026 592650 154646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 174026 592650 174646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 214026 592650 214646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 234026 592650 234646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 254026 592650 254646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 274026 592650 274646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 294026 592650 294646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 314026 592650 314646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 334026 592650 334646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 354026 592650 354646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 394026 592650 394646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 414026 592650 414646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 434026 592650 434646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 454026 592650 454646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 474026 592650 474646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 494026 592650 494646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 514026 592650 514646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 534026 592650 534646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 574026 592650 574646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 594026 592650 594646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 614026 592650 614646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 634026 592650 634646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 654026 592650 654646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 674026 592650 674646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 694026 592650 694646 6 vdda2
port 535 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 -7654 73574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 -7654 93574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 -7654 113574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 -7654 133574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 -7654 153574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 172954 -7654 173574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 -7654 233574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 -7654 253574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 -7654 273574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 -7654 293574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 -7654 313574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 -7654 333574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 -7654 353574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 -7654 393574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 -7654 413574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 -7654 433574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 -7654 453574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 -7654 473574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 -7654 493574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 -7654 513574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 145308 73574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 145308 93574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 145308 113574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 145308 133574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 145308 153574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 172954 145308 173574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 145308 193574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 145308 233574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 145308 253574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 145308 273574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 145308 293574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 145308 313574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 145308 333574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 145308 353574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 145308 393574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 145308 413574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 145308 433574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 145308 453574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 145308 473574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 145308 493574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 145308 513574 165000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 252308 73574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 252308 93574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 252308 113574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 252308 133574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 252308 153574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 172954 252308 173574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 252308 193574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 252308 233574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 252308 253574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 252308 273574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 252308 293574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 252308 313574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 252308 333574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 252308 353574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 252308 393574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 252308 413574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 252308 433574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 252308 453574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 252308 473574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 252308 493574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 252308 513574 272000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 359308 73574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 359308 93574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 359308 113574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 359308 133574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 359308 153574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 172954 359308 173574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 359308 193574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 359308 233574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 359308 253574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 359308 273574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 359308 293574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 359308 313574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 359308 333574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 359308 353574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 359308 393574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 359308 413574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 359308 433574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 359308 453574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 359308 473574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 359308 493574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 359308 513574 379000 6 vdda2
port 535 nsew power input
rlabel metal4 s 212954 -7654 213574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 466308 233574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 466308 253574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 466308 273574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 466308 293574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 466308 313574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 466308 353574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 -7654 373574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 466308 393574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 466308 413574 491000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 466308 453574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 466308 473574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 466308 493574 501000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 466308 73574 521000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 466308 93574 521000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 466308 113574 521000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 466308 133574 521000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 466308 153574 521000 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 558099 353574 578000 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 558099 373574 578000 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 558099 393574 578000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 558099 413574 578000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 555000 453574 578000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 555000 473574 578000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 555000 493574 578000 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 466308 513574 578000 6 vdda2
port 535 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 32954 -7654 33574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 52954 -7654 53574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 636033 73574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 636033 93574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 636033 113574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 636033 133574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 636033 153574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 172954 466308 173574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 466308 193574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 212954 642000 213574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 642000 233574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 642000 253574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 642000 273574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 642000 293574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 642000 313574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 466308 333574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 645099 353574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 645099 373574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 645099 393574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 645099 413574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 466308 433574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 645099 453574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 645099 473574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 645099 493574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 645099 513574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 532954 -7654 533574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 572954 -7654 573574 711590 6 vdda2
port 535 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 20306 590730 20926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 40306 590730 40926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 60306 590730 60926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 80306 590730 80926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 120306 590730 120926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 140306 590730 140926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 160306 590730 160926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 180306 590730 180926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 200306 590730 200926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 220306 590730 220926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 240306 590730 240926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 260306 590730 260926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 300306 590730 300926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 320306 590730 320926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 340306 590730 340926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 360306 590730 360926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 380306 590730 380926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 400306 590730 400926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 420306 590730 420926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 440306 590730 440926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 480306 590730 480926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 500306 590730 500926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 520306 590730 520926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 540306 590730 540926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 560306 590730 560926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 580306 590730 580926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 600306 590730 600926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 620306 590730 620926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 660306 590730 660926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 680306 590730 680926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 700306 590730 700926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 -5734 59854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 -5734 79854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 -5734 119854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 -5734 139854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 -5734 159854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 179234 -5734 179854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 -5734 219854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 -5734 239854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 -5734 259854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 -5734 299854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 -5734 319854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 339234 -5734 339854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 -5734 379854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 -5734 399854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 -5734 419854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 -5734 439854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 -5734 479854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 -5734 499854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 145308 59854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 145308 79854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 145308 99854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 145308 119854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 145308 139854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 145308 159854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 179234 145308 179854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 145308 219854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 145308 239854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 145308 259854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 145308 279854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 145308 299854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 145308 319854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 339234 145308 339854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 145308 379854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 145308 399854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 145308 419854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 145308 439854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 145308 459854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 145308 479854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 145308 499854 165000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 252308 59854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 252308 79854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 252308 99854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 252308 119854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 252308 139854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 252308 159854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 179234 252308 179854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 252308 219854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 252308 239854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 252308 259854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 252308 279854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 252308 299854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 252308 319854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 339234 252308 339854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 252308 379854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 252308 399854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 252308 419854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 252308 439854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 252308 459854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 252308 479854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 252308 499854 272000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 359308 59854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 359308 79854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 359308 99854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 359308 119854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 359308 139854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 359308 159854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 179234 359308 179854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 359308 219854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 359308 239854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 359308 259854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 359308 279854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 359308 299854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 359308 319854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 339234 359308 339854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 359308 379854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 359308 399854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 359308 419854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 359308 439854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 359308 459854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 359308 479854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 359308 499854 379000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 199234 -5734 199854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 466308 219854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 466308 239854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 466308 259854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 466308 279854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 466308 299854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 466308 319854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 359234 -5734 359854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 466308 379854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 466308 399854 491000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 466308 459854 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 466308 479854 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 466308 499854 501000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 466308 59854 521000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 466308 79854 521000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 466308 99854 521000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 466308 119854 521000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 466308 139854 521000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 466308 159854 521000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 359234 558099 359854 578000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 558099 379854 578000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 558099 399854 578000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 555000 459854 578000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 555000 479854 578000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 555000 499854 578000 6 vssa1
port 536 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground input
rlabel metal4 s 19234 -5734 19854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 39234 -5734 39854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 636033 59854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 636033 79854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 636033 99854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 636033 119854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 636033 139854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 636033 159854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 179234 466308 179854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 199234 642000 199854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 642000 219854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 642000 239854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 642000 259854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 642000 279854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 642000 299854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 642000 319854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 339234 466308 339854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 359234 645099 359854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 645099 379854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 645099 399854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 466308 419854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 466308 439854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 645099 459854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 645099 479854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 645099 499854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 519234 -5734 519854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 539234 -5734 539854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 559234 -5734 559854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 579234 -5734 579854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 24026 592650 24646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 44026 592650 44646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 64026 592650 64646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 84026 592650 84646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 124026 592650 124646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 144026 592650 144646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 164026 592650 164646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 184026 592650 184646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 204026 592650 204646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 224026 592650 224646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 244026 592650 244646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 264026 592650 264646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 304026 592650 304646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 324026 592650 324646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 344026 592650 344646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 364026 592650 364646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 384026 592650 384646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 404026 592650 404646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 424026 592650 424646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 444026 592650 444646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 484026 592650 484646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 504026 592650 504646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 524026 592650 524646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 544026 592650 544646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 564026 592650 564646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 584026 592650 584646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 604026 592650 604646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 624026 592650 624646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 664026 592650 664646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 684026 592650 684646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 -7654 63574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 -7654 83574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 -7654 123574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 -7654 143574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 -7654 163574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 182954 -7654 183574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 -7654 223574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 -7654 243574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 -7654 263574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 -7654 303574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 -7654 323574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 342954 -7654 343574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 -7654 383574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 -7654 403574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 -7654 423574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 -7654 443574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 -7654 483574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 -7654 503574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 145308 63574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 145308 83574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 145308 103574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 145308 123574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 145308 143574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 145308 163574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 182954 145308 183574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 145308 223574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 145308 243574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 145308 263574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 145308 283574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 145308 303574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 145308 323574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 342954 145308 343574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 145308 383574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 145308 403574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 145308 423574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 145308 443574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 145308 463574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 145308 483574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 145308 503574 165000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 252308 63574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 252308 83574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 252308 103574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 252308 123574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 252308 143574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 252308 163574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 182954 252308 183574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 252308 223574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 252308 243574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 252308 263574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 252308 283574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 252308 303574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 252308 323574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 342954 252308 343574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 252308 383574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 252308 403574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 252308 423574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 252308 443574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 252308 463574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 252308 483574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 252308 503574 272000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 359308 63574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 359308 83574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 359308 103574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 359308 123574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 359308 143574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 359308 163574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 182954 359308 183574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 359308 223574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 359308 243574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 359308 263574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 359308 283574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 359308 303574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 359308 323574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 342954 359308 343574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 359308 383574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 359308 403574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 359308 423574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 359308 443574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 359308 463574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 359308 483574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 359308 503574 379000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 202954 -7654 203574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 466308 223574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 466308 243574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 466308 263574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 466308 283574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 466308 303574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 362954 -7654 363574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 466308 383574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 466308 403574 491000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 466308 463574 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 466308 483574 501000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 466308 63574 521000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 466308 83574 521000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 466308 103574 521000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 466308 123574 521000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 466308 143574 521000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 466308 163574 521000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 362954 558099 363574 578000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 558099 383574 578000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 558099 403574 578000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 555000 463574 578000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 555000 483574 578000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 466308 503574 578000 6 vssa2
port 537 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground input
rlabel metal4 s 22954 -7654 23574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 42954 -7654 43574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 636033 63574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 636033 83574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 636033 103574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 636033 123574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 636033 143574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 636033 163574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 182954 466308 183574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 202954 642000 203574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 642000 223574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 642000 243574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 642000 263574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 642000 283574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 642000 303574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 466308 323574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 342954 466308 343574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 362954 645099 363574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 645099 383574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 645099 403574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 466308 423574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 466308 443574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 645099 463574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 645099 483574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 645099 503574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 522954 -7654 523574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 542954 -7654 543574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 562954 -7654 563574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 12866 586890 13486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 32866 586890 33486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 52866 586890 53486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 72866 586890 73486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 112866 586890 113486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 132866 586890 133486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 152866 586890 153486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 172866 586890 173486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 192866 586890 193486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 212866 586890 213486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 232866 586890 233486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 252866 586890 253486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 292866 586890 293486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 312866 586890 313486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 332866 586890 333486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 352866 586890 353486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 372866 586890 373486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 392866 586890 393486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 412866 586890 413486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 432866 586890 433486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 472866 586890 473486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 492866 586890 493486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 512866 586890 513486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 532866 586890 533486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 552866 586890 553486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 572866 586890 573486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 592866 586890 593486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 612866 586890 613486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 652866 586890 653486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 672866 586890 673486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 692866 586890 693486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 -1894 72414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 -1894 112414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 -1894 132414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 -1894 152414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 171794 -1894 172414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 191794 -1894 192414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 -1894 232414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 -1894 252414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 -1894 292414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 -1894 312414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 -1894 332414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 -1894 352414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 -1894 392414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 -1894 412414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 -1894 432414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 -1894 472414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 -1894 492414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 -1894 512414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 145308 72414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 145308 92414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 145308 112414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 145308 132414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 145308 152414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 171794 145308 172414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 191794 145308 192414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 145308 232414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 145308 252414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 145308 272414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 145308 292414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 145308 312414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 145308 332414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 145308 352414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 145308 392414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 145308 412414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 145308 432414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 145308 452414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 145308 472414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 145308 492414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 145308 512414 165000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 252308 72414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 252308 92414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 252308 112414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 252308 132414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 252308 152414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 171794 252308 172414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 191794 252308 192414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 252308 232414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 252308 252414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 252308 272414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 252308 292414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 252308 312414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 252308 332414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 252308 352414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 252308 392414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 252308 412414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 252308 432414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 252308 452414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 252308 472414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 252308 492414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 252308 512414 272000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 359308 72414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 359308 92414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 359308 112414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 359308 132414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 359308 152414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 171794 359308 172414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 191794 359308 192414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 359308 232414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 359308 252414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 359308 272414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 359308 292414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 359308 312414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 359308 332414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 359308 352414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 359308 392414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 359308 412414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 359308 432414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 359308 452414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 359308 472414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 359308 492414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 359308 512414 379000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211794 -1894 212414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 466308 232414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 466308 252414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 466308 272414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 466308 292414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 466308 312414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 371794 -1894 372414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 466308 392414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 466308 412414 491000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 466308 452414 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 466308 472414 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 466308 492414 501000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 466308 72414 521000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 466308 92414 521000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 466308 112414 521000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 466308 132414 521000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 466308 152414 521000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 371794 558099 372414 578000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 558099 392414 578000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 558099 412414 578000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 555000 452414 578000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 555000 472414 578000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 555000 492414 578000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 466308 512414 578000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground input
rlabel metal4 s 11794 -1894 12414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 31794 -1894 32414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 51794 -1894 52414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 636033 72414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 636033 92414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 636033 112414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 636033 132414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 636033 152414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 171794 466308 172414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 191794 466308 192414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211794 642000 212414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 642000 232414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 642000 252414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 642000 272414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 642000 292414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 642000 312414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 466308 332414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 466308 352414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 371794 645099 372414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 645099 392414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 645099 412414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 466308 432414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 645099 452414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 645099 472414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 645099 492414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 645099 512414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 531794 -1894 532414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 551794 -1894 552414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 571794 -1894 572414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 16586 588810 17206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 36586 588810 37206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 56586 588810 57206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 76586 588810 77206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 116586 588810 117206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 136586 588810 137206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 156586 588810 157206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 176586 588810 177206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 196586 588810 197206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 216586 588810 217206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 236586 588810 237206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 256586 588810 257206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 296586 588810 297206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 316586 588810 317206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 336586 588810 337206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 356586 588810 357206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 376586 588810 377206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 396586 588810 397206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 416586 588810 417206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 436586 588810 437206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 476586 588810 477206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 496586 588810 497206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 516586 588810 517206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 536586 588810 537206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 556586 588810 557206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 576586 588810 577206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 596586 588810 597206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 616586 588810 617206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 656586 588810 657206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 676586 588810 677206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 696586 588810 697206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 -3814 76134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 -3814 116134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 -3814 136134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 -3814 156134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 175514 -3814 176134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 195514 -3814 196134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 -3814 236134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 -3814 256134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 -3814 296134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 -3814 316134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 -3814 336134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 -3814 356134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 -3814 396134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 -3814 416134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 -3814 436134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 -3814 476134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 -3814 496134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 515514 -3814 516134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 145308 76134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 145308 96134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 145308 116134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 145308 136134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 145308 156134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 175514 145308 176134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 195514 145308 196134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 145308 236134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 145308 256134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 145308 276134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 145308 296134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 145308 316134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 145308 336134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 145308 356134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 145308 396134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 145308 416134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 145308 436134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 145308 456134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 145308 476134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 145308 496134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 515514 145308 516134 165000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 252308 76134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 252308 96134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 252308 116134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 252308 136134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 252308 156134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 175514 252308 176134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 195514 252308 196134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 252308 236134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 252308 256134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 252308 276134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 252308 296134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 252308 316134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 252308 336134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 252308 356134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 252308 396134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 252308 416134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 252308 436134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 252308 456134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 252308 476134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 252308 496134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 515514 252308 516134 272000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 359308 76134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 359308 96134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 359308 116134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 359308 136134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 359308 156134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 175514 359308 176134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 195514 359308 196134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 359308 236134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 359308 256134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 359308 276134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 359308 296134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 359308 316134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 359308 336134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 359308 356134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 359308 396134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 359308 416134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 359308 436134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 359308 456134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 359308 476134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 359308 496134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 515514 359308 516134 379000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215514 -3814 216134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 466308 236134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 466308 256134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 466308 276134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 466308 296134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 466308 316134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 466308 356134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 375514 -3814 376134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 466308 396134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 466308 416134 491000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 466308 456134 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 466308 476134 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 466308 496134 501000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 466308 76134 521000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 466308 96134 521000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 466308 116134 521000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 466308 136134 521000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 466308 156134 521000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 558099 356134 578000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 375514 558099 376134 578000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 558099 396134 578000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 558099 416134 578000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 555000 456134 578000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 555000 476134 578000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 555000 496134 578000 6 vssd2
port 539 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground input
rlabel metal4 s 15514 -3814 16134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 35514 -3814 36134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 55514 -3814 56134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 636033 76134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 636033 96134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 636033 116134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 636033 136134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 636033 156134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 175514 466308 176134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 195514 466308 196134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215514 642000 216134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 642000 236134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 642000 256134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 642000 276134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 642000 296134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 642000 316134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 466308 336134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 645099 356134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 375514 645099 376134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 645099 396134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 645099 416134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 466308 436134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 645099 456134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 645099 476134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 645099 496134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 515514 466308 516134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 535514 -3814 536134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 555514 -3814 556134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 575514 -3814 576134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 95497000
string GDS_FILE /home/burak/asic_tools/caravel_vscpu3x/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 90644312
<< end >>

