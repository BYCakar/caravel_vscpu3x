magic
tech sky130A
magscale 1 2
timestamp 1655395919
<< obsli1 >>
rect 61104 482159 508852 628817
<< obsm1 >>
rect 566 3408 580506 700392
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 580502 703610
rect 572 536 580502 703464
rect 710 480 1590 536
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6374 536
rect 6598 480 7570 536
rect 7794 480 8674 536
rect 8898 480 9870 536
rect 10094 480 11066 536
rect 11290 480 12262 536
rect 12486 480 13458 536
rect 13682 480 14654 536
rect 14878 480 15850 536
rect 16074 480 16954 536
rect 17178 480 18150 536
rect 18374 480 19346 536
rect 19570 480 20542 536
rect 20766 480 21738 536
rect 21962 480 22934 536
rect 23158 480 24130 536
rect 24354 480 25234 536
rect 25458 480 26430 536
rect 26654 480 27626 536
rect 27850 480 28822 536
rect 29046 480 30018 536
rect 30242 480 31214 536
rect 31438 480 32318 536
rect 32542 480 33514 536
rect 33738 480 34710 536
rect 34934 480 35906 536
rect 36130 480 37102 536
rect 37326 480 38298 536
rect 38522 480 39494 536
rect 39718 480 40598 536
rect 40822 480 41794 536
rect 42018 480 42990 536
rect 43214 480 44186 536
rect 44410 480 45382 536
rect 45606 480 46578 536
rect 46802 480 47774 536
rect 47998 480 48878 536
rect 49102 480 50074 536
rect 50298 480 51270 536
rect 51494 480 52466 536
rect 52690 480 53662 536
rect 53886 480 54858 536
rect 55082 480 55962 536
rect 56186 480 57158 536
rect 57382 480 58354 536
rect 58578 480 59550 536
rect 59774 480 60746 536
rect 60970 480 61942 536
rect 62166 480 63138 536
rect 63362 480 64242 536
rect 64466 480 65438 536
rect 65662 480 66634 536
rect 66858 480 67830 536
rect 68054 480 69026 536
rect 69250 480 70222 536
rect 70446 480 71418 536
rect 71642 480 72522 536
rect 72746 480 73718 536
rect 73942 480 74914 536
rect 75138 480 76110 536
rect 76334 480 77306 536
rect 77530 480 78502 536
rect 78726 480 79606 536
rect 79830 480 80802 536
rect 81026 480 81998 536
rect 82222 480 83194 536
rect 83418 480 84390 536
rect 84614 480 85586 536
rect 85810 480 86782 536
rect 87006 480 87886 536
rect 88110 480 89082 536
rect 89306 480 90278 536
rect 90502 480 91474 536
rect 91698 480 92670 536
rect 92894 480 93866 536
rect 94090 480 95062 536
rect 95286 480 96166 536
rect 96390 480 97362 536
rect 97586 480 98558 536
rect 98782 480 99754 536
rect 99978 480 100950 536
rect 101174 480 102146 536
rect 102370 480 103250 536
rect 103474 480 104446 536
rect 104670 480 105642 536
rect 105866 480 106838 536
rect 107062 480 108034 536
rect 108258 480 109230 536
rect 109454 480 110426 536
rect 110650 480 111530 536
rect 111754 480 112726 536
rect 112950 480 113922 536
rect 114146 480 115118 536
rect 115342 480 116314 536
rect 116538 480 117510 536
rect 117734 480 118706 536
rect 118930 480 119810 536
rect 120034 480 121006 536
rect 121230 480 122202 536
rect 122426 480 123398 536
rect 123622 480 124594 536
rect 124818 480 125790 536
rect 126014 480 126894 536
rect 127118 480 128090 536
rect 128314 480 129286 536
rect 129510 480 130482 536
rect 130706 480 131678 536
rect 131902 480 132874 536
rect 133098 480 134070 536
rect 134294 480 135174 536
rect 135398 480 136370 536
rect 136594 480 137566 536
rect 137790 480 138762 536
rect 138986 480 139958 536
rect 140182 480 141154 536
rect 141378 480 142350 536
rect 142574 480 143454 536
rect 143678 480 144650 536
rect 144874 480 145846 536
rect 146070 480 147042 536
rect 147266 480 148238 536
rect 148462 480 149434 536
rect 149658 480 150538 536
rect 150762 480 151734 536
rect 151958 480 152930 536
rect 153154 480 154126 536
rect 154350 480 155322 536
rect 155546 480 156518 536
rect 156742 480 157714 536
rect 157938 480 158818 536
rect 159042 480 160014 536
rect 160238 480 161210 536
rect 161434 480 162406 536
rect 162630 480 163602 536
rect 163826 480 164798 536
rect 165022 480 165994 536
rect 166218 480 167098 536
rect 167322 480 168294 536
rect 168518 480 169490 536
rect 169714 480 170686 536
rect 170910 480 171882 536
rect 172106 480 173078 536
rect 173302 480 174182 536
rect 174406 480 175378 536
rect 175602 480 176574 536
rect 176798 480 177770 536
rect 177994 480 178966 536
rect 179190 480 180162 536
rect 180386 480 181358 536
rect 181582 480 182462 536
rect 182686 480 183658 536
rect 183882 480 184854 536
rect 185078 480 186050 536
rect 186274 480 187246 536
rect 187470 480 188442 536
rect 188666 480 189638 536
rect 189862 480 190742 536
rect 190966 480 191938 536
rect 192162 480 193134 536
rect 193358 480 194330 536
rect 194554 480 195526 536
rect 195750 480 196722 536
rect 196946 480 197826 536
rect 198050 480 199022 536
rect 199246 480 200218 536
rect 200442 480 201414 536
rect 201638 480 202610 536
rect 202834 480 203806 536
rect 204030 480 205002 536
rect 205226 480 206106 536
rect 206330 480 207302 536
rect 207526 480 208498 536
rect 208722 480 209694 536
rect 209918 480 210890 536
rect 211114 480 212086 536
rect 212310 480 213282 536
rect 213506 480 214386 536
rect 214610 480 215582 536
rect 215806 480 216778 536
rect 217002 480 217974 536
rect 218198 480 219170 536
rect 219394 480 220366 536
rect 220590 480 221470 536
rect 221694 480 222666 536
rect 222890 480 223862 536
rect 224086 480 225058 536
rect 225282 480 226254 536
rect 226478 480 227450 536
rect 227674 480 228646 536
rect 228870 480 229750 536
rect 229974 480 230946 536
rect 231170 480 232142 536
rect 232366 480 233338 536
rect 233562 480 234534 536
rect 234758 480 235730 536
rect 235954 480 236926 536
rect 237150 480 238030 536
rect 238254 480 239226 536
rect 239450 480 240422 536
rect 240646 480 241618 536
rect 241842 480 242814 536
rect 243038 480 244010 536
rect 244234 480 245114 536
rect 245338 480 246310 536
rect 246534 480 247506 536
rect 247730 480 248702 536
rect 248926 480 249898 536
rect 250122 480 251094 536
rect 251318 480 252290 536
rect 252514 480 253394 536
rect 253618 480 254590 536
rect 254814 480 255786 536
rect 256010 480 256982 536
rect 257206 480 258178 536
rect 258402 480 259374 536
rect 259598 480 260570 536
rect 260794 480 261674 536
rect 261898 480 262870 536
rect 263094 480 264066 536
rect 264290 480 265262 536
rect 265486 480 266458 536
rect 266682 480 267654 536
rect 267878 480 268758 536
rect 268982 480 269954 536
rect 270178 480 271150 536
rect 271374 480 272346 536
rect 272570 480 273542 536
rect 273766 480 274738 536
rect 274962 480 275934 536
rect 276158 480 277038 536
rect 277262 480 278234 536
rect 278458 480 279430 536
rect 279654 480 280626 536
rect 280850 480 281822 536
rect 282046 480 283018 536
rect 283242 480 284214 536
rect 284438 480 285318 536
rect 285542 480 286514 536
rect 286738 480 287710 536
rect 287934 480 288906 536
rect 289130 480 290102 536
rect 290326 480 291298 536
rect 291522 480 292494 536
rect 292718 480 293598 536
rect 293822 480 294794 536
rect 295018 480 295990 536
rect 296214 480 297186 536
rect 297410 480 298382 536
rect 298606 480 299578 536
rect 299802 480 300682 536
rect 300906 480 301878 536
rect 302102 480 303074 536
rect 303298 480 304270 536
rect 304494 480 305466 536
rect 305690 480 306662 536
rect 306886 480 307858 536
rect 308082 480 308962 536
rect 309186 480 310158 536
rect 310382 480 311354 536
rect 311578 480 312550 536
rect 312774 480 313746 536
rect 313970 480 314942 536
rect 315166 480 316138 536
rect 316362 480 317242 536
rect 317466 480 318438 536
rect 318662 480 319634 536
rect 319858 480 320830 536
rect 321054 480 322026 536
rect 322250 480 323222 536
rect 323446 480 324326 536
rect 324550 480 325522 536
rect 325746 480 326718 536
rect 326942 480 327914 536
rect 328138 480 329110 536
rect 329334 480 330306 536
rect 330530 480 331502 536
rect 331726 480 332606 536
rect 332830 480 333802 536
rect 334026 480 334998 536
rect 335222 480 336194 536
rect 336418 480 337390 536
rect 337614 480 338586 536
rect 338810 480 339782 536
rect 340006 480 340886 536
rect 341110 480 342082 536
rect 342306 480 343278 536
rect 343502 480 344474 536
rect 344698 480 345670 536
rect 345894 480 346866 536
rect 347090 480 347970 536
rect 348194 480 349166 536
rect 349390 480 350362 536
rect 350586 480 351558 536
rect 351782 480 352754 536
rect 352978 480 353950 536
rect 354174 480 355146 536
rect 355370 480 356250 536
rect 356474 480 357446 536
rect 357670 480 358642 536
rect 358866 480 359838 536
rect 360062 480 361034 536
rect 361258 480 362230 536
rect 362454 480 363426 536
rect 363650 480 364530 536
rect 364754 480 365726 536
rect 365950 480 366922 536
rect 367146 480 368118 536
rect 368342 480 369314 536
rect 369538 480 370510 536
rect 370734 480 371614 536
rect 371838 480 372810 536
rect 373034 480 374006 536
rect 374230 480 375202 536
rect 375426 480 376398 536
rect 376622 480 377594 536
rect 377818 480 378790 536
rect 379014 480 379894 536
rect 380118 480 381090 536
rect 381314 480 382286 536
rect 382510 480 383482 536
rect 383706 480 384678 536
rect 384902 480 385874 536
rect 386098 480 387070 536
rect 387294 480 388174 536
rect 388398 480 389370 536
rect 389594 480 390566 536
rect 390790 480 391762 536
rect 391986 480 392958 536
rect 393182 480 394154 536
rect 394378 480 395258 536
rect 395482 480 396454 536
rect 396678 480 397650 536
rect 397874 480 398846 536
rect 399070 480 400042 536
rect 400266 480 401238 536
rect 401462 480 402434 536
rect 402658 480 403538 536
rect 403762 480 404734 536
rect 404958 480 405930 536
rect 406154 480 407126 536
rect 407350 480 408322 536
rect 408546 480 409518 536
rect 409742 480 410714 536
rect 410938 480 411818 536
rect 412042 480 413014 536
rect 413238 480 414210 536
rect 414434 480 415406 536
rect 415630 480 416602 536
rect 416826 480 417798 536
rect 418022 480 418902 536
rect 419126 480 420098 536
rect 420322 480 421294 536
rect 421518 480 422490 536
rect 422714 480 423686 536
rect 423910 480 424882 536
rect 425106 480 426078 536
rect 426302 480 427182 536
rect 427406 480 428378 536
rect 428602 480 429574 536
rect 429798 480 430770 536
rect 430994 480 431966 536
rect 432190 480 433162 536
rect 433386 480 434358 536
rect 434582 480 435462 536
rect 435686 480 436658 536
rect 436882 480 437854 536
rect 438078 480 439050 536
rect 439274 480 440246 536
rect 440470 480 441442 536
rect 441666 480 442546 536
rect 442770 480 443742 536
rect 443966 480 444938 536
rect 445162 480 446134 536
rect 446358 480 447330 536
rect 447554 480 448526 536
rect 448750 480 449722 536
rect 449946 480 450826 536
rect 451050 480 452022 536
rect 452246 480 453218 536
rect 453442 480 454414 536
rect 454638 480 455610 536
rect 455834 480 456806 536
rect 457030 480 458002 536
rect 458226 480 459106 536
rect 459330 480 460302 536
rect 460526 480 461498 536
rect 461722 480 462694 536
rect 462918 480 463890 536
rect 464114 480 465086 536
rect 465310 480 466190 536
rect 466414 480 467386 536
rect 467610 480 468582 536
rect 468806 480 469778 536
rect 470002 480 470974 536
rect 471198 480 472170 536
rect 472394 480 473366 536
rect 473590 480 474470 536
rect 474694 480 475666 536
rect 475890 480 476862 536
rect 477086 480 478058 536
rect 478282 480 479254 536
rect 479478 480 480450 536
rect 480674 480 481646 536
rect 481870 480 482750 536
rect 482974 480 483946 536
rect 484170 480 485142 536
rect 485366 480 486338 536
rect 486562 480 487534 536
rect 487758 480 488730 536
rect 488954 480 489834 536
rect 490058 480 491030 536
rect 491254 480 492226 536
rect 492450 480 493422 536
rect 493646 480 494618 536
rect 494842 480 495814 536
rect 496038 480 497010 536
rect 497234 480 498114 536
rect 498338 480 499310 536
rect 499534 480 500506 536
rect 500730 480 501702 536
rect 501926 480 502898 536
rect 503122 480 504094 536
rect 504318 480 505290 536
rect 505514 480 506394 536
rect 506618 480 507590 536
rect 507814 480 508786 536
rect 509010 480 509982 536
rect 510206 480 511178 536
rect 511402 480 512374 536
rect 512598 480 513478 536
rect 513702 480 514674 536
rect 514898 480 515870 536
rect 516094 480 517066 536
rect 517290 480 518262 536
rect 518486 480 519458 536
rect 519682 480 520654 536
rect 520878 480 521758 536
rect 521982 480 522954 536
rect 523178 480 524150 536
rect 524374 480 525346 536
rect 525570 480 526542 536
rect 526766 480 527738 536
rect 527962 480 528934 536
rect 529158 480 530038 536
rect 530262 480 531234 536
rect 531458 480 532430 536
rect 532654 480 533626 536
rect 533850 480 534822 536
rect 535046 480 536018 536
rect 536242 480 537122 536
rect 537346 480 538318 536
rect 538542 480 539514 536
rect 539738 480 540710 536
rect 540934 480 541906 536
rect 542130 480 543102 536
rect 543326 480 544298 536
rect 544522 480 545402 536
rect 545626 480 546598 536
rect 546822 480 547794 536
rect 548018 480 548990 536
rect 549214 480 550186 536
rect 550410 480 551382 536
rect 551606 480 552578 536
rect 552802 480 553682 536
rect 553906 480 554878 536
rect 555102 480 556074 536
rect 556298 480 557270 536
rect 557494 480 558466 536
rect 558690 480 559662 536
rect 559886 480 560766 536
rect 560990 480 561962 536
rect 562186 480 563158 536
rect 563382 480 564354 536
rect 564578 480 565550 536
rect 565774 480 566746 536
rect 566970 480 567942 536
rect 568166 480 569046 536
rect 569270 480 570242 536
rect 570466 480 571438 536
rect 571662 480 572634 536
rect 572858 480 573830 536
rect 574054 480 575026 536
rect 575250 480 576222 536
rect 576446 480 577326 536
rect 577550 480 578522 536
rect 578746 480 579718 536
rect 579942 480 580502 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 560 684084 583520 684317
rect 246 684076 583520 684084
rect 246 683676 583440 684076
rect 246 671428 583520 683676
rect 560 671028 583520 671428
rect 246 670884 583520 671028
rect 246 670484 583440 670884
rect 246 658372 583520 670484
rect 560 657972 583520 658372
rect 246 657556 583520 657972
rect 246 657156 583440 657556
rect 246 645316 583520 657156
rect 560 644916 583520 645316
rect 246 644228 583520 644916
rect 246 643828 583440 644228
rect 246 632260 583520 643828
rect 560 631860 583520 632260
rect 246 631036 583520 631860
rect 246 630636 583440 631036
rect 246 619340 583520 630636
rect 560 618940 583520 619340
rect 246 617708 583520 618940
rect 246 617308 583440 617708
rect 246 606284 583520 617308
rect 560 605884 583520 606284
rect 246 604380 583520 605884
rect 246 603980 583440 604380
rect 246 593228 583520 603980
rect 560 592828 583520 593228
rect 246 591188 583520 592828
rect 246 590788 583440 591188
rect 246 580172 583520 590788
rect 560 579772 583520 580172
rect 246 577860 583520 579772
rect 246 577460 583440 577860
rect 246 567116 583520 577460
rect 560 566716 583520 567116
rect 246 564532 583520 566716
rect 246 564132 583440 564532
rect 246 554060 583520 564132
rect 560 553660 583520 554060
rect 246 551340 583520 553660
rect 246 550940 583440 551340
rect 246 541004 583520 550940
rect 560 540604 583520 541004
rect 246 538012 583520 540604
rect 246 537612 583440 538012
rect 246 528084 583520 537612
rect 560 527684 583520 528084
rect 246 524684 583520 527684
rect 246 524284 583440 524684
rect 246 515028 583520 524284
rect 560 514628 583520 515028
rect 246 511492 583520 514628
rect 246 511092 583440 511492
rect 246 501972 583520 511092
rect 560 501572 583520 501972
rect 246 498164 583520 501572
rect 246 497764 583440 498164
rect 246 488916 583520 497764
rect 560 488516 583520 488916
rect 246 484836 583520 488516
rect 246 484436 583440 484836
rect 246 475860 583520 484436
rect 560 475460 583520 475860
rect 246 471644 583520 475460
rect 246 471244 583440 471644
rect 246 462804 583520 471244
rect 560 462404 583520 462804
rect 246 458316 583520 462404
rect 246 457916 583440 458316
rect 246 449748 583520 457916
rect 560 449348 583520 449748
rect 246 444988 583520 449348
rect 246 444588 583440 444988
rect 246 436828 583520 444588
rect 560 436428 583520 436828
rect 246 431796 583520 436428
rect 246 431396 583440 431796
rect 246 423772 583520 431396
rect 560 423372 583520 423772
rect 246 418468 583520 423372
rect 246 418068 583440 418468
rect 246 410716 583520 418068
rect 560 410316 583520 410716
rect 246 405140 583520 410316
rect 246 404740 583440 405140
rect 246 397660 583520 404740
rect 560 397260 583520 397660
rect 246 391948 583520 397260
rect 246 391548 583440 391948
rect 246 384604 583520 391548
rect 560 384204 583520 384604
rect 246 378620 583520 384204
rect 246 378220 583440 378620
rect 246 371548 583520 378220
rect 560 371148 583520 371548
rect 246 365292 583520 371148
rect 246 364892 583440 365292
rect 246 358628 583520 364892
rect 560 358228 583520 358628
rect 246 352100 583520 358228
rect 246 351700 583440 352100
rect 246 345572 583520 351700
rect 560 345172 583520 345572
rect 246 338772 583520 345172
rect 246 338372 583440 338772
rect 246 332516 583520 338372
rect 560 332116 583520 332516
rect 246 325444 583520 332116
rect 246 325044 583440 325444
rect 246 319460 583520 325044
rect 560 319060 583520 319460
rect 246 312252 583520 319060
rect 246 311852 583440 312252
rect 246 306404 583520 311852
rect 560 306004 583520 306404
rect 246 298924 583520 306004
rect 246 298524 583440 298924
rect 246 293348 583520 298524
rect 560 292948 583520 293348
rect 246 285596 583520 292948
rect 246 285196 583440 285596
rect 246 280292 583520 285196
rect 560 279892 583520 280292
rect 246 272404 583520 279892
rect 246 272004 583440 272404
rect 246 267372 583520 272004
rect 560 266972 583520 267372
rect 246 259076 583520 266972
rect 246 258676 583440 259076
rect 246 254316 583520 258676
rect 560 253916 583520 254316
rect 246 245748 583520 253916
rect 246 245348 583440 245748
rect 246 241260 583520 245348
rect 560 240860 583520 241260
rect 246 232556 583520 240860
rect 246 232156 583440 232556
rect 246 228204 583520 232156
rect 560 227804 583520 228204
rect 246 219228 583520 227804
rect 246 218828 583440 219228
rect 246 215148 583520 218828
rect 560 214748 583520 215148
rect 246 205900 583520 214748
rect 246 205500 583440 205900
rect 246 202092 583520 205500
rect 560 201692 583520 202092
rect 246 192708 583520 201692
rect 246 192308 583440 192708
rect 246 189036 583520 192308
rect 560 188636 583520 189036
rect 246 179380 583520 188636
rect 246 178980 583440 179380
rect 246 176116 583520 178980
rect 560 175716 583520 176116
rect 246 166052 583520 175716
rect 246 165652 583440 166052
rect 246 163060 583520 165652
rect 560 162660 583520 163060
rect 246 152860 583520 162660
rect 246 152460 583440 152860
rect 246 150004 583520 152460
rect 560 149604 583520 150004
rect 246 139532 583520 149604
rect 246 139132 583440 139532
rect 246 136948 583520 139132
rect 560 136548 583520 136948
rect 246 126204 583520 136548
rect 246 125804 583440 126204
rect 246 123892 583520 125804
rect 560 123492 583520 123892
rect 246 113012 583520 123492
rect 246 112612 583440 113012
rect 246 110836 583520 112612
rect 560 110436 583520 110836
rect 246 99684 583520 110436
rect 246 99284 583440 99684
rect 246 97780 583520 99284
rect 560 97380 583520 97780
rect 246 86356 583520 97380
rect 246 85956 583440 86356
rect 246 84860 583520 85956
rect 560 84460 583520 84860
rect 246 73164 583520 84460
rect 246 72764 583440 73164
rect 246 71804 583520 72764
rect 560 71404 583520 71804
rect 246 59836 583520 71404
rect 246 59436 583440 59836
rect 246 58748 583520 59436
rect 560 58348 583520 58748
rect 246 46508 583520 58348
rect 246 46108 583440 46508
rect 246 45692 583520 46108
rect 560 45292 583520 45692
rect 246 33316 583520 45292
rect 246 32916 583440 33316
rect 246 32636 583520 32916
rect 560 32236 583520 32636
rect 246 19988 583520 32236
rect 246 19588 583440 19988
rect 246 19580 583520 19588
rect 560 19347 583520 19580
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 -5734 9854 709670
rect 12954 -7654 13574 711590
rect 19794 -1894 20414 705830
rect 23514 -3814 24134 707750
rect 27234 -5734 27854 709670
rect 30954 -7654 31574 711590
rect 37794 -1894 38414 705830
rect 41514 -3814 42134 707750
rect 45234 -5734 45854 709670
rect 48954 -7654 49574 711590
rect 55794 -1894 56414 705830
rect 59514 625099 60134 707750
rect 63234 625099 63854 709670
rect 66954 625099 67574 711590
rect 73794 625099 74414 705830
rect 77514 625099 78134 707750
rect 81234 625099 81854 709670
rect 84954 625099 85574 711590
rect 91794 625099 92414 705830
rect 95514 625099 96134 707750
rect 99234 625099 99854 709670
rect 102954 625099 103574 711590
rect 109794 625099 110414 705830
rect 113514 625099 114134 707750
rect 117234 625099 117854 709670
rect 120954 625099 121574 711590
rect 59514 542000 60134 558000
rect 63234 542000 63854 558000
rect 66954 542000 67574 558000
rect 73794 542000 74414 558000
rect 77514 542000 78134 558000
rect 81234 542000 81854 558000
rect 84954 542000 85574 558000
rect 91794 542000 92414 558000
rect 95514 542000 96134 558000
rect 99234 542000 99854 558000
rect 102954 542000 103574 558000
rect 109794 542000 110414 558000
rect 113514 542000 114134 558000
rect 117234 542000 117854 558000
rect 120954 542000 121574 558000
rect 127794 542000 128414 705830
rect 131514 542000 132134 707750
rect 135234 542000 135854 709670
rect 138954 625099 139574 711590
rect 145794 625099 146414 705830
rect 149514 625099 150134 707750
rect 153234 625099 153854 709670
rect 156954 625099 157574 711590
rect 163794 625099 164414 705830
rect 167514 625099 168134 707750
rect 171234 625099 171854 709670
rect 174954 625099 175574 711590
rect 181794 625099 182414 705830
rect 185514 625099 186134 707750
rect 189234 625099 189854 709670
rect 192954 625099 193574 711590
rect 199794 625099 200414 705830
rect 138954 542000 139574 558000
rect 145794 542000 146414 558000
rect 149514 542000 150134 558000
rect 153234 542000 153854 558000
rect 156954 542000 157574 558000
rect 163794 542000 164414 558000
rect 167514 542000 168134 558000
rect 171234 542000 171854 558000
rect 174954 542000 175574 558000
rect 181794 542000 182414 558000
rect 185514 542000 186134 558000
rect 189234 542000 189854 558000
rect 192954 542000 193574 558000
rect 199794 542000 200414 558000
rect 203514 542000 204134 707750
rect 207234 542000 207854 709670
rect 210954 542000 211574 711590
rect 217794 625099 218414 705830
rect 221514 625099 222134 707750
rect 225234 625099 225854 709670
rect 228954 625099 229574 711590
rect 235794 625099 236414 705830
rect 239514 625099 240134 707750
rect 243234 625099 243854 709670
rect 246954 625099 247574 711590
rect 253794 625099 254414 705830
rect 257514 625099 258134 707750
rect 261234 625099 261854 709670
rect 264954 625099 265574 711590
rect 271794 625099 272414 705830
rect 275514 625099 276134 707750
rect 279234 625099 279854 709670
rect 282954 625099 283574 711590
rect 217794 542000 218414 558000
rect 221514 542000 222134 558000
rect 225234 542000 225854 558000
rect 228954 542000 229574 558000
rect 235794 542000 236414 558000
rect 239514 542000 240134 558000
rect 243234 542000 243854 558000
rect 246954 542000 247574 558000
rect 253794 542000 254414 558000
rect 257514 542000 258134 558000
rect 261234 542000 261854 558000
rect 264954 542000 265574 558000
rect 271794 542000 272414 558000
rect 275514 542000 276134 558000
rect 279234 542000 279854 558000
rect 282954 542000 283574 558000
rect 289794 542000 290414 705830
rect 293514 542000 294134 707750
rect 297234 542000 297854 709670
rect 300954 542000 301574 711590
rect 59514 460308 60134 478000
rect 63234 460308 63854 478000
rect 66954 460308 67574 478000
rect 73794 460308 74414 478000
rect 77514 460308 78134 478000
rect 81234 460308 81854 478000
rect 84954 460308 85574 478000
rect 91794 460308 92414 478000
rect 95514 460308 96134 478000
rect 99234 460308 99854 478000
rect 102954 460308 103574 478000
rect 109794 460308 110414 478000
rect 113514 460308 114134 478000
rect 117234 460308 117854 478000
rect 120954 460308 121574 478000
rect 127794 460308 128414 478000
rect 131514 460308 132134 478000
rect 135234 460308 135854 478000
rect 138954 460308 139574 478000
rect 145794 460308 146414 478000
rect 149514 460308 150134 478000
rect 153234 460308 153854 478000
rect 156954 460308 157574 478000
rect 163794 460308 164414 478000
rect 167514 460308 168134 478000
rect 171234 460308 171854 478000
rect 174954 460308 175574 478000
rect 181794 460308 182414 478000
rect 185514 460308 186134 478000
rect 189234 460308 189854 478000
rect 192954 460308 193574 478000
rect 59514 355308 60134 373000
rect 63234 355308 63854 373000
rect 66954 355308 67574 373000
rect 73794 355308 74414 373000
rect 77514 355308 78134 373000
rect 81234 355308 81854 373000
rect 84954 355308 85574 373000
rect 91794 355308 92414 373000
rect 95514 355308 96134 373000
rect 99234 355308 99854 373000
rect 102954 355308 103574 373000
rect 109794 355308 110414 373000
rect 113514 355308 114134 373000
rect 117234 355308 117854 373000
rect 120954 355308 121574 373000
rect 127794 355308 128414 373000
rect 131514 355308 132134 373000
rect 135234 355308 135854 373000
rect 138954 355308 139574 373000
rect 145794 355308 146414 373000
rect 149514 355308 150134 373000
rect 153234 355308 153854 373000
rect 156954 355308 157574 373000
rect 163794 355308 164414 373000
rect 167514 355308 168134 373000
rect 171234 355308 171854 373000
rect 174954 355308 175574 373000
rect 181794 355308 182414 373000
rect 185514 355308 186134 373000
rect 189234 355308 189854 373000
rect 192954 355308 193574 373000
rect 59514 250308 60134 268000
rect 63234 250308 63854 268000
rect 66954 250308 67574 268000
rect 73794 250308 74414 268000
rect 77514 250308 78134 268000
rect 81234 250308 81854 268000
rect 84954 250308 85574 268000
rect 91794 250308 92414 268000
rect 95514 250308 96134 268000
rect 99234 250308 99854 268000
rect 102954 250308 103574 268000
rect 109794 250308 110414 268000
rect 113514 250308 114134 268000
rect 117234 250308 117854 268000
rect 120954 250308 121574 268000
rect 127794 250308 128414 268000
rect 131514 250308 132134 268000
rect 135234 250308 135854 268000
rect 138954 250308 139574 268000
rect 145794 250308 146414 268000
rect 149514 250308 150134 268000
rect 153234 250308 153854 268000
rect 156954 250308 157574 268000
rect 163794 250308 164414 268000
rect 167514 250308 168134 268000
rect 171234 250308 171854 268000
rect 174954 250308 175574 268000
rect 181794 250308 182414 268000
rect 185514 250308 186134 268000
rect 189234 250308 189854 268000
rect 192954 250308 193574 268000
rect 59514 145308 60134 163000
rect 63234 145308 63854 163000
rect 66954 145308 67574 163000
rect 73794 145308 74414 163000
rect 77514 145308 78134 163000
rect 81234 145308 81854 163000
rect 84954 145308 85574 163000
rect 91794 145308 92414 163000
rect 95514 145308 96134 163000
rect 99234 145308 99854 163000
rect 102954 145308 103574 163000
rect 109794 145308 110414 163000
rect 113514 145308 114134 163000
rect 117234 145308 117854 163000
rect 120954 145308 121574 163000
rect 127794 145308 128414 163000
rect 131514 145308 132134 163000
rect 135234 145308 135854 163000
rect 138954 145308 139574 163000
rect 145794 145308 146414 163000
rect 149514 145308 150134 163000
rect 153234 145308 153854 163000
rect 156954 145308 157574 163000
rect 163794 145308 164414 163000
rect 167514 145308 168134 163000
rect 171234 145308 171854 163000
rect 174954 145308 175574 163000
rect 181794 145308 182414 163000
rect 185514 145308 186134 163000
rect 189234 145308 189854 163000
rect 192954 145308 193574 163000
rect 59514 -3814 60134 58000
rect 63234 -5734 63854 58000
rect 66954 -7654 67574 58000
rect 73794 -1894 74414 58000
rect 77514 -3814 78134 58000
rect 81234 -5734 81854 58000
rect 84954 -7654 85574 58000
rect 91794 -1894 92414 58000
rect 95514 -3814 96134 58000
rect 99234 -5734 99854 58000
rect 102954 -7654 103574 58000
rect 109794 -1894 110414 58000
rect 113514 -3814 114134 58000
rect 117234 -5734 117854 58000
rect 120954 -7654 121574 58000
rect 127794 -1894 128414 58000
rect 131514 -3814 132134 58000
rect 135234 -5734 135854 58000
rect 138954 -7654 139574 58000
rect 145794 -1894 146414 58000
rect 149514 -3814 150134 58000
rect 153234 -5734 153854 58000
rect 156954 -7654 157574 58000
rect 163794 -1894 164414 58000
rect 167514 -3814 168134 58000
rect 171234 -5734 171854 58000
rect 174954 -7654 175574 58000
rect 181794 -1894 182414 58000
rect 185514 -3814 186134 58000
rect 189234 -5734 189854 58000
rect 192954 -7654 193574 58000
rect 199794 -1894 200414 478000
rect 203514 -3814 204134 478000
rect 207234 -5734 207854 478000
rect 210954 -7654 211574 478000
rect 217794 460308 218414 478000
rect 221514 460308 222134 478000
rect 225234 460308 225854 478000
rect 228954 460308 229574 478000
rect 235794 460308 236414 478000
rect 239514 460308 240134 478000
rect 243234 460308 243854 478000
rect 246954 460308 247574 478000
rect 253794 460308 254414 478000
rect 257514 460308 258134 478000
rect 261234 460308 261854 478000
rect 264954 460308 265574 478000
rect 271794 460308 272414 478000
rect 275514 460308 276134 478000
rect 279234 460308 279854 478000
rect 282954 460308 283574 478000
rect 289794 460308 290414 478000
rect 293514 460308 294134 478000
rect 297234 460308 297854 478000
rect 300954 460308 301574 478000
rect 307794 460308 308414 705830
rect 311514 460308 312134 707750
rect 315234 460308 315854 709670
rect 318954 633033 319574 711590
rect 325794 633033 326414 705830
rect 329514 633033 330134 707750
rect 333234 633033 333854 709670
rect 336954 633033 337574 711590
rect 343794 633033 344414 705830
rect 347514 633033 348134 707750
rect 351234 633033 351854 709670
rect 354954 633033 355574 711590
rect 361794 633033 362414 705830
rect 365514 633033 366134 707750
rect 369234 633033 369854 709670
rect 372954 633033 373574 711590
rect 379794 633033 380414 705830
rect 383514 633033 384134 707750
rect 387234 633033 387854 709670
rect 390954 633033 391574 711590
rect 397794 633033 398414 705830
rect 401514 633033 402134 707750
rect 405234 633033 405854 709670
rect 408954 633033 409574 711590
rect 415794 633033 416414 705830
rect 419514 633033 420134 707750
rect 423234 633033 423854 709670
rect 426954 633033 427574 711590
rect 318954 460308 319574 518000
rect 325794 460308 326414 518000
rect 329514 460308 330134 518000
rect 333234 460308 333854 518000
rect 336954 460308 337574 518000
rect 343794 460308 344414 518000
rect 347514 460308 348134 518000
rect 351234 460308 351854 518000
rect 354954 460308 355574 518000
rect 217794 355308 218414 373000
rect 221514 355308 222134 373000
rect 225234 355308 225854 373000
rect 228954 355308 229574 373000
rect 235794 355308 236414 373000
rect 239514 355308 240134 373000
rect 243234 355308 243854 373000
rect 246954 355308 247574 373000
rect 253794 355308 254414 373000
rect 257514 355308 258134 373000
rect 261234 355308 261854 373000
rect 264954 355308 265574 373000
rect 271794 355308 272414 373000
rect 275514 355308 276134 373000
rect 279234 355308 279854 373000
rect 282954 355308 283574 373000
rect 289794 355308 290414 373000
rect 293514 355308 294134 373000
rect 297234 355308 297854 373000
rect 300954 355308 301574 373000
rect 307794 355308 308414 373000
rect 311514 355308 312134 373000
rect 315234 355308 315854 373000
rect 318954 355308 319574 373000
rect 325794 355308 326414 373000
rect 329514 355308 330134 373000
rect 333234 355308 333854 373000
rect 336954 355308 337574 373000
rect 343794 355308 344414 373000
rect 347514 355308 348134 373000
rect 351234 355308 351854 373000
rect 354954 355308 355574 373000
rect 217794 250308 218414 268000
rect 221514 250308 222134 268000
rect 225234 250308 225854 268000
rect 228954 250308 229574 268000
rect 235794 250308 236414 268000
rect 239514 250308 240134 268000
rect 243234 250308 243854 268000
rect 246954 250308 247574 268000
rect 253794 250308 254414 268000
rect 257514 250308 258134 268000
rect 261234 250308 261854 268000
rect 264954 250308 265574 268000
rect 271794 250308 272414 268000
rect 275514 250308 276134 268000
rect 279234 250308 279854 268000
rect 282954 250308 283574 268000
rect 289794 250308 290414 268000
rect 293514 250308 294134 268000
rect 297234 250308 297854 268000
rect 300954 250308 301574 268000
rect 307794 250308 308414 268000
rect 311514 250308 312134 268000
rect 315234 250308 315854 268000
rect 318954 250308 319574 268000
rect 325794 250308 326414 268000
rect 329514 250308 330134 268000
rect 333234 250308 333854 268000
rect 336954 250308 337574 268000
rect 343794 250308 344414 268000
rect 347514 250308 348134 268000
rect 351234 250308 351854 268000
rect 354954 250308 355574 268000
rect 217794 145308 218414 163000
rect 221514 145308 222134 163000
rect 225234 145308 225854 163000
rect 228954 145308 229574 163000
rect 235794 145308 236414 163000
rect 239514 145308 240134 163000
rect 243234 145308 243854 163000
rect 246954 145308 247574 163000
rect 253794 145308 254414 163000
rect 257514 145308 258134 163000
rect 261234 145308 261854 163000
rect 264954 145308 265574 163000
rect 271794 145308 272414 163000
rect 275514 145308 276134 163000
rect 279234 145308 279854 163000
rect 282954 145308 283574 163000
rect 289794 145308 290414 163000
rect 293514 145308 294134 163000
rect 297234 145308 297854 163000
rect 300954 145308 301574 163000
rect 307794 145308 308414 163000
rect 311514 145308 312134 163000
rect 315234 145308 315854 163000
rect 318954 145308 319574 163000
rect 325794 145308 326414 163000
rect 329514 145308 330134 163000
rect 333234 145308 333854 163000
rect 336954 145308 337574 163000
rect 343794 145308 344414 163000
rect 347514 145308 348134 163000
rect 351234 145308 351854 163000
rect 354954 145308 355574 163000
rect 217794 -1894 218414 58000
rect 221514 -3814 222134 58000
rect 225234 -5734 225854 58000
rect 228954 -7654 229574 58000
rect 235794 -1894 236414 58000
rect 239514 -3814 240134 58000
rect 243234 -5734 243854 58000
rect 246954 -7654 247574 58000
rect 253794 -1894 254414 58000
rect 257514 -3814 258134 58000
rect 261234 -5734 261854 58000
rect 264954 -7654 265574 58000
rect 271794 -1894 272414 58000
rect 275514 -3814 276134 58000
rect 279234 -5734 279854 58000
rect 282954 -7654 283574 58000
rect 289794 -1894 290414 58000
rect 293514 -3814 294134 58000
rect 297234 -5734 297854 58000
rect 300954 -7654 301574 58000
rect 307794 -1894 308414 58000
rect 311514 -3814 312134 58000
rect 315234 -5734 315854 58000
rect 318954 -7654 319574 58000
rect 325794 -1894 326414 58000
rect 329514 -3814 330134 58000
rect 333234 -5734 333854 58000
rect 336954 -7654 337574 58000
rect 343794 -1894 344414 58000
rect 347514 -3814 348134 58000
rect 351234 -5734 351854 58000
rect 354954 -7654 355574 58000
rect 361794 -1894 362414 518000
rect 365514 -3814 366134 518000
rect 369234 -5734 369854 518000
rect 372954 -7654 373574 518000
rect 379794 460308 380414 518000
rect 383514 460308 384134 518000
rect 387234 460308 387854 518000
rect 390954 460308 391574 518000
rect 397794 460308 398414 518000
rect 401514 460308 402134 518000
rect 405234 460308 405854 518000
rect 408954 460308 409574 518000
rect 415794 460308 416414 518000
rect 419514 460308 420134 518000
rect 423234 460308 423854 518000
rect 426954 460308 427574 518000
rect 433794 460308 434414 705830
rect 437514 460308 438134 707750
rect 441234 460308 441854 709670
rect 444954 460308 445574 711590
rect 451794 460308 452414 705830
rect 455514 460308 456134 707750
rect 459234 622000 459854 709670
rect 462954 622000 463574 711590
rect 469794 622000 470414 705830
rect 473514 622000 474134 707750
rect 477234 622000 477854 709670
rect 480954 622000 481574 711590
rect 487794 622000 488414 705830
rect 491514 622000 492134 707750
rect 495234 622000 495854 709670
rect 498954 622000 499574 711590
rect 505794 622000 506414 705830
rect 509514 622000 510134 707750
rect 459234 460308 459854 568000
rect 462954 460308 463574 568000
rect 469794 460308 470414 568000
rect 473514 460308 474134 568000
rect 477234 460308 477854 568000
rect 480954 460308 481574 568000
rect 487794 460308 488414 568000
rect 491514 460308 492134 568000
rect 495234 460308 495854 568000
rect 498954 460308 499574 568000
rect 505794 460308 506414 568000
rect 509514 460308 510134 568000
rect 513234 460308 513854 709670
rect 516954 460308 517574 711590
rect 379794 355308 380414 373000
rect 383514 355308 384134 373000
rect 387234 355308 387854 373000
rect 390954 355308 391574 373000
rect 397794 355308 398414 373000
rect 401514 355308 402134 373000
rect 405234 355308 405854 373000
rect 408954 355308 409574 373000
rect 415794 355308 416414 373000
rect 419514 355308 420134 373000
rect 423234 355308 423854 373000
rect 426954 355308 427574 373000
rect 433794 355308 434414 373000
rect 437514 355308 438134 373000
rect 441234 355308 441854 373000
rect 444954 355308 445574 373000
rect 451794 355308 452414 373000
rect 455514 355308 456134 373000
rect 459234 355308 459854 373000
rect 462954 355308 463574 373000
rect 469794 355308 470414 373000
rect 473514 355308 474134 373000
rect 477234 355308 477854 373000
rect 480954 355308 481574 373000
rect 487794 355308 488414 373000
rect 491514 355308 492134 373000
rect 495234 355308 495854 373000
rect 498954 355308 499574 373000
rect 505794 355308 506414 373000
rect 509514 355308 510134 373000
rect 513234 355308 513854 373000
rect 516954 355308 517574 373000
rect 379794 250308 380414 268000
rect 383514 250308 384134 268000
rect 387234 250308 387854 268000
rect 390954 250308 391574 268000
rect 397794 250308 398414 268000
rect 401514 250308 402134 268000
rect 405234 250308 405854 268000
rect 408954 250308 409574 268000
rect 415794 250308 416414 268000
rect 419514 250308 420134 268000
rect 423234 250308 423854 268000
rect 426954 250308 427574 268000
rect 433794 250308 434414 268000
rect 437514 250308 438134 268000
rect 441234 250308 441854 268000
rect 444954 250308 445574 268000
rect 451794 250308 452414 268000
rect 455514 250308 456134 268000
rect 459234 250308 459854 268000
rect 462954 250308 463574 268000
rect 469794 250308 470414 268000
rect 473514 250308 474134 268000
rect 477234 250308 477854 268000
rect 480954 250308 481574 268000
rect 487794 250308 488414 268000
rect 491514 250308 492134 268000
rect 495234 250308 495854 268000
rect 498954 250308 499574 268000
rect 505794 250308 506414 268000
rect 509514 250308 510134 268000
rect 513234 250308 513854 268000
rect 516954 250308 517574 268000
rect 379794 145308 380414 163000
rect 383514 145308 384134 163000
rect 387234 145308 387854 163000
rect 390954 145308 391574 163000
rect 397794 145308 398414 163000
rect 401514 145308 402134 163000
rect 405234 145308 405854 163000
rect 408954 145308 409574 163000
rect 415794 145308 416414 163000
rect 419514 145308 420134 163000
rect 423234 145308 423854 163000
rect 426954 145308 427574 163000
rect 433794 145308 434414 163000
rect 437514 145308 438134 163000
rect 441234 145308 441854 163000
rect 444954 145308 445574 163000
rect 451794 145308 452414 163000
rect 455514 145308 456134 163000
rect 459234 145308 459854 163000
rect 462954 145308 463574 163000
rect 469794 145308 470414 163000
rect 473514 145308 474134 163000
rect 477234 145308 477854 163000
rect 480954 145308 481574 163000
rect 487794 145308 488414 163000
rect 491514 145308 492134 163000
rect 495234 145308 495854 163000
rect 498954 145308 499574 163000
rect 505794 145308 506414 163000
rect 509514 145308 510134 163000
rect 513234 145308 513854 163000
rect 516954 145308 517574 163000
rect 379794 -1894 380414 58000
rect 383514 -3814 384134 58000
rect 387234 -5734 387854 58000
rect 390954 -7654 391574 58000
rect 397794 -1894 398414 58000
rect 401514 -3814 402134 58000
rect 405234 -5734 405854 58000
rect 408954 -7654 409574 58000
rect 415794 -1894 416414 58000
rect 419514 -3814 420134 58000
rect 423234 -5734 423854 58000
rect 426954 -7654 427574 58000
rect 433794 -1894 434414 58000
rect 437514 -3814 438134 58000
rect 441234 -5734 441854 58000
rect 444954 -7654 445574 58000
rect 451794 -1894 452414 58000
rect 455514 -3814 456134 58000
rect 459234 -5734 459854 58000
rect 462954 -7654 463574 58000
rect 469794 -1894 470414 58000
rect 473514 -3814 474134 58000
rect 477234 -5734 477854 58000
rect 480954 -7654 481574 58000
rect 487794 -1894 488414 58000
rect 491514 -3814 492134 58000
rect 495234 -5734 495854 58000
rect 498954 -7654 499574 58000
rect 505794 -1894 506414 58000
rect 509514 -3814 510134 58000
rect 513234 -5734 513854 58000
rect 516954 -7654 517574 58000
rect 523794 -1894 524414 705830
rect 527514 -3814 528134 707750
rect 531234 -5734 531854 709670
rect 534954 -7654 535574 711590
rect 541794 -1894 542414 705830
rect 545514 -3814 546134 707750
rect 549234 -5734 549854 709670
rect 552954 -7654 553574 711590
rect 559794 -1894 560414 705830
rect 563514 -3814 564134 707750
rect 567234 -5734 567854 709670
rect 570954 -7654 571574 711590
rect 577794 -1894 578414 705830
rect 581514 -3814 582134 707750
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 44955 54707 45154 630869
rect 45934 54707 48874 630869
rect 49654 54707 55714 630869
rect 56494 625019 59434 630869
rect 60214 625019 63154 630869
rect 63934 625019 66874 630869
rect 67654 625019 73714 630869
rect 74494 625019 77434 630869
rect 78214 625019 81154 630869
rect 81934 625019 84874 630869
rect 85654 625019 91714 630869
rect 92494 625019 95434 630869
rect 96214 625019 99154 630869
rect 99934 625019 102874 630869
rect 103654 625019 109714 630869
rect 110494 625019 113434 630869
rect 114214 625019 117154 630869
rect 117934 625019 120874 630869
rect 121654 625019 127714 630869
rect 56494 558080 127714 625019
rect 56494 541920 59434 558080
rect 60214 541920 63154 558080
rect 63934 541920 66874 558080
rect 67654 541920 73714 558080
rect 74494 541920 77434 558080
rect 78214 541920 81154 558080
rect 81934 541920 84874 558080
rect 85654 541920 91714 558080
rect 92494 541920 95434 558080
rect 96214 541920 99154 558080
rect 99934 541920 102874 558080
rect 103654 541920 109714 558080
rect 110494 541920 113434 558080
rect 114214 541920 117154 558080
rect 117934 541920 120874 558080
rect 121654 541920 127714 558080
rect 128494 541920 131434 630869
rect 132214 541920 135154 630869
rect 135934 625019 138874 630869
rect 139654 625019 145714 630869
rect 146494 625019 149434 630869
rect 150214 625019 153154 630869
rect 153934 625019 156874 630869
rect 157654 625019 163714 630869
rect 164494 625019 167434 630869
rect 168214 625019 171154 630869
rect 171934 625019 174874 630869
rect 175654 625019 181714 630869
rect 182494 625019 185434 630869
rect 186214 625019 189154 630869
rect 189934 625019 192874 630869
rect 193654 625019 199714 630869
rect 200494 625019 203434 630869
rect 135934 558080 203434 625019
rect 135934 541920 138874 558080
rect 139654 541920 145714 558080
rect 146494 541920 149434 558080
rect 150214 541920 153154 558080
rect 153934 541920 156874 558080
rect 157654 541920 163714 558080
rect 164494 541920 167434 558080
rect 168214 541920 171154 558080
rect 171934 541920 174874 558080
rect 175654 541920 181714 558080
rect 182494 541920 185434 558080
rect 186214 541920 189154 558080
rect 189934 541920 192874 558080
rect 193654 541920 199714 558080
rect 200494 541920 203434 558080
rect 204214 541920 207154 630869
rect 207934 541920 210874 630869
rect 211654 625019 217714 630869
rect 218494 625019 221434 630869
rect 222214 625019 225154 630869
rect 225934 625019 228874 630869
rect 229654 625019 235714 630869
rect 236494 625019 239434 630869
rect 240214 625019 243154 630869
rect 243934 625019 246874 630869
rect 247654 625019 253714 630869
rect 254494 625019 257434 630869
rect 258214 625019 261154 630869
rect 261934 625019 264874 630869
rect 265654 625019 271714 630869
rect 272494 625019 275434 630869
rect 276214 625019 279154 630869
rect 279934 625019 282874 630869
rect 283654 625019 289714 630869
rect 211654 558080 289714 625019
rect 211654 541920 217714 558080
rect 218494 541920 221434 558080
rect 222214 541920 225154 558080
rect 225934 541920 228874 558080
rect 229654 541920 235714 558080
rect 236494 541920 239434 558080
rect 240214 541920 243154 558080
rect 243934 541920 246874 558080
rect 247654 541920 253714 558080
rect 254494 541920 257434 558080
rect 258214 541920 261154 558080
rect 261934 541920 264874 558080
rect 265654 541920 271714 558080
rect 272494 541920 275434 558080
rect 276214 541920 279154 558080
rect 279934 541920 282874 558080
rect 283654 541920 289714 558080
rect 290494 541920 293434 630869
rect 294214 541920 297154 630869
rect 297934 541920 300874 630869
rect 301654 541920 307714 630869
rect 56494 478080 307714 541920
rect 56494 460228 59434 478080
rect 60214 460228 63154 478080
rect 63934 460228 66874 478080
rect 67654 460228 73714 478080
rect 74494 460228 77434 478080
rect 78214 460228 81154 478080
rect 81934 460228 84874 478080
rect 85654 460228 91714 478080
rect 92494 460228 95434 478080
rect 96214 460228 99154 478080
rect 99934 460228 102874 478080
rect 103654 460228 109714 478080
rect 110494 460228 113434 478080
rect 114214 460228 117154 478080
rect 117934 460228 120874 478080
rect 121654 460228 127714 478080
rect 128494 460228 131434 478080
rect 132214 460228 135154 478080
rect 135934 460228 138874 478080
rect 139654 460228 145714 478080
rect 146494 460228 149434 478080
rect 150214 460228 153154 478080
rect 153934 460228 156874 478080
rect 157654 460228 163714 478080
rect 164494 460228 167434 478080
rect 168214 460228 171154 478080
rect 171934 460228 174874 478080
rect 175654 460228 181714 478080
rect 182494 460228 185434 478080
rect 186214 460228 189154 478080
rect 189934 460228 192874 478080
rect 193654 460228 199714 478080
rect 56494 373080 199714 460228
rect 56494 355228 59434 373080
rect 60214 355228 63154 373080
rect 63934 355228 66874 373080
rect 67654 355228 73714 373080
rect 74494 355228 77434 373080
rect 78214 355228 81154 373080
rect 81934 355228 84874 373080
rect 85654 355228 91714 373080
rect 92494 355228 95434 373080
rect 96214 355228 99154 373080
rect 99934 355228 102874 373080
rect 103654 355228 109714 373080
rect 110494 355228 113434 373080
rect 114214 355228 117154 373080
rect 117934 355228 120874 373080
rect 121654 355228 127714 373080
rect 128494 355228 131434 373080
rect 132214 355228 135154 373080
rect 135934 355228 138874 373080
rect 139654 355228 145714 373080
rect 146494 355228 149434 373080
rect 150214 355228 153154 373080
rect 153934 355228 156874 373080
rect 157654 355228 163714 373080
rect 164494 355228 167434 373080
rect 168214 355228 171154 373080
rect 171934 355228 174874 373080
rect 175654 355228 181714 373080
rect 182494 355228 185434 373080
rect 186214 355228 189154 373080
rect 189934 355228 192874 373080
rect 193654 355228 199714 373080
rect 56494 268080 199714 355228
rect 56494 250228 59434 268080
rect 60214 250228 63154 268080
rect 63934 250228 66874 268080
rect 67654 250228 73714 268080
rect 74494 250228 77434 268080
rect 78214 250228 81154 268080
rect 81934 250228 84874 268080
rect 85654 250228 91714 268080
rect 92494 250228 95434 268080
rect 96214 250228 99154 268080
rect 99934 250228 102874 268080
rect 103654 250228 109714 268080
rect 110494 250228 113434 268080
rect 114214 250228 117154 268080
rect 117934 250228 120874 268080
rect 121654 250228 127714 268080
rect 128494 250228 131434 268080
rect 132214 250228 135154 268080
rect 135934 250228 138874 268080
rect 139654 250228 145714 268080
rect 146494 250228 149434 268080
rect 150214 250228 153154 268080
rect 153934 250228 156874 268080
rect 157654 250228 163714 268080
rect 164494 250228 167434 268080
rect 168214 250228 171154 268080
rect 171934 250228 174874 268080
rect 175654 250228 181714 268080
rect 182494 250228 185434 268080
rect 186214 250228 189154 268080
rect 189934 250228 192874 268080
rect 193654 250228 199714 268080
rect 56494 163080 199714 250228
rect 56494 145228 59434 163080
rect 60214 145228 63154 163080
rect 63934 145228 66874 163080
rect 67654 145228 73714 163080
rect 74494 145228 77434 163080
rect 78214 145228 81154 163080
rect 81934 145228 84874 163080
rect 85654 145228 91714 163080
rect 92494 145228 95434 163080
rect 96214 145228 99154 163080
rect 99934 145228 102874 163080
rect 103654 145228 109714 163080
rect 110494 145228 113434 163080
rect 114214 145228 117154 163080
rect 117934 145228 120874 163080
rect 121654 145228 127714 163080
rect 128494 145228 131434 163080
rect 132214 145228 135154 163080
rect 135934 145228 138874 163080
rect 139654 145228 145714 163080
rect 146494 145228 149434 163080
rect 150214 145228 153154 163080
rect 153934 145228 156874 163080
rect 157654 145228 163714 163080
rect 164494 145228 167434 163080
rect 168214 145228 171154 163080
rect 171934 145228 174874 163080
rect 175654 145228 181714 163080
rect 182494 145228 185434 163080
rect 186214 145228 189154 163080
rect 189934 145228 192874 163080
rect 193654 145228 199714 163080
rect 56494 58080 199714 145228
rect 56494 54707 59434 58080
rect 60214 54707 63154 58080
rect 63934 54707 66874 58080
rect 67654 54707 73714 58080
rect 74494 54707 77434 58080
rect 78214 54707 81154 58080
rect 81934 54707 84874 58080
rect 85654 54707 91714 58080
rect 92494 54707 95434 58080
rect 96214 54707 99154 58080
rect 99934 54707 102874 58080
rect 103654 54707 109714 58080
rect 110494 54707 113434 58080
rect 114214 54707 117154 58080
rect 117934 54707 120874 58080
rect 121654 54707 127714 58080
rect 128494 54707 131434 58080
rect 132214 54707 135154 58080
rect 135934 54707 138874 58080
rect 139654 54707 145714 58080
rect 146494 54707 149434 58080
rect 150214 54707 153154 58080
rect 153934 54707 156874 58080
rect 157654 54707 163714 58080
rect 164494 54707 167434 58080
rect 168214 54707 171154 58080
rect 171934 54707 174874 58080
rect 175654 54707 181714 58080
rect 182494 54707 185434 58080
rect 186214 54707 189154 58080
rect 189934 54707 192874 58080
rect 193654 54707 199714 58080
rect 200494 54707 203434 478080
rect 204214 54707 207154 478080
rect 207934 54707 210874 478080
rect 211654 460228 217714 478080
rect 218494 460228 221434 478080
rect 222214 460228 225154 478080
rect 225934 460228 228874 478080
rect 229654 460228 235714 478080
rect 236494 460228 239434 478080
rect 240214 460228 243154 478080
rect 243934 460228 246874 478080
rect 247654 460228 253714 478080
rect 254494 460228 257434 478080
rect 258214 460228 261154 478080
rect 261934 460228 264874 478080
rect 265654 460228 271714 478080
rect 272494 460228 275434 478080
rect 276214 460228 279154 478080
rect 279934 460228 282874 478080
rect 283654 460228 289714 478080
rect 290494 460228 293434 478080
rect 294214 460228 297154 478080
rect 297934 460228 300874 478080
rect 301654 460228 307714 478080
rect 308494 460228 311434 630869
rect 312214 460228 315154 630869
rect 315934 518080 433714 630869
rect 315934 460228 318874 518080
rect 319654 460228 325714 518080
rect 326494 460228 329434 518080
rect 330214 460228 333154 518080
rect 333934 460228 336874 518080
rect 337654 460228 343714 518080
rect 344494 460228 347434 518080
rect 348214 460228 351154 518080
rect 351934 460228 354874 518080
rect 355654 460228 361714 518080
rect 211654 373080 361714 460228
rect 211654 355228 217714 373080
rect 218494 355228 221434 373080
rect 222214 355228 225154 373080
rect 225934 355228 228874 373080
rect 229654 355228 235714 373080
rect 236494 355228 239434 373080
rect 240214 355228 243154 373080
rect 243934 355228 246874 373080
rect 247654 355228 253714 373080
rect 254494 355228 257434 373080
rect 258214 355228 261154 373080
rect 261934 355228 264874 373080
rect 265654 355228 271714 373080
rect 272494 355228 275434 373080
rect 276214 355228 279154 373080
rect 279934 355228 282874 373080
rect 283654 355228 289714 373080
rect 290494 355228 293434 373080
rect 294214 355228 297154 373080
rect 297934 355228 300874 373080
rect 301654 355228 307714 373080
rect 308494 355228 311434 373080
rect 312214 355228 315154 373080
rect 315934 355228 318874 373080
rect 319654 355228 325714 373080
rect 326494 355228 329434 373080
rect 330214 355228 333154 373080
rect 333934 355228 336874 373080
rect 337654 355228 343714 373080
rect 344494 355228 347434 373080
rect 348214 355228 351154 373080
rect 351934 355228 354874 373080
rect 355654 355228 361714 373080
rect 211654 268080 361714 355228
rect 211654 250228 217714 268080
rect 218494 250228 221434 268080
rect 222214 250228 225154 268080
rect 225934 250228 228874 268080
rect 229654 250228 235714 268080
rect 236494 250228 239434 268080
rect 240214 250228 243154 268080
rect 243934 250228 246874 268080
rect 247654 250228 253714 268080
rect 254494 250228 257434 268080
rect 258214 250228 261154 268080
rect 261934 250228 264874 268080
rect 265654 250228 271714 268080
rect 272494 250228 275434 268080
rect 276214 250228 279154 268080
rect 279934 250228 282874 268080
rect 283654 250228 289714 268080
rect 290494 250228 293434 268080
rect 294214 250228 297154 268080
rect 297934 250228 300874 268080
rect 301654 250228 307714 268080
rect 308494 250228 311434 268080
rect 312214 250228 315154 268080
rect 315934 250228 318874 268080
rect 319654 250228 325714 268080
rect 326494 250228 329434 268080
rect 330214 250228 333154 268080
rect 333934 250228 336874 268080
rect 337654 250228 343714 268080
rect 344494 250228 347434 268080
rect 348214 250228 351154 268080
rect 351934 250228 354874 268080
rect 355654 250228 361714 268080
rect 211654 163080 361714 250228
rect 211654 145228 217714 163080
rect 218494 145228 221434 163080
rect 222214 145228 225154 163080
rect 225934 145228 228874 163080
rect 229654 145228 235714 163080
rect 236494 145228 239434 163080
rect 240214 145228 243154 163080
rect 243934 145228 246874 163080
rect 247654 145228 253714 163080
rect 254494 145228 257434 163080
rect 258214 145228 261154 163080
rect 261934 145228 264874 163080
rect 265654 145228 271714 163080
rect 272494 145228 275434 163080
rect 276214 145228 279154 163080
rect 279934 145228 282874 163080
rect 283654 145228 289714 163080
rect 290494 145228 293434 163080
rect 294214 145228 297154 163080
rect 297934 145228 300874 163080
rect 301654 145228 307714 163080
rect 308494 145228 311434 163080
rect 312214 145228 315154 163080
rect 315934 145228 318874 163080
rect 319654 145228 325714 163080
rect 326494 145228 329434 163080
rect 330214 145228 333154 163080
rect 333934 145228 336874 163080
rect 337654 145228 343714 163080
rect 344494 145228 347434 163080
rect 348214 145228 351154 163080
rect 351934 145228 354874 163080
rect 355654 145228 361714 163080
rect 211654 58080 361714 145228
rect 211654 54707 217714 58080
rect 218494 54707 221434 58080
rect 222214 54707 225154 58080
rect 225934 54707 228874 58080
rect 229654 54707 235714 58080
rect 236494 54707 239434 58080
rect 240214 54707 243154 58080
rect 243934 54707 246874 58080
rect 247654 54707 253714 58080
rect 254494 54707 257434 58080
rect 258214 54707 261154 58080
rect 261934 54707 264874 58080
rect 265654 54707 271714 58080
rect 272494 54707 275434 58080
rect 276214 54707 279154 58080
rect 279934 54707 282874 58080
rect 283654 54707 289714 58080
rect 290494 54707 293434 58080
rect 294214 54707 297154 58080
rect 297934 54707 300874 58080
rect 301654 54707 307714 58080
rect 308494 54707 311434 58080
rect 312214 54707 315154 58080
rect 315934 54707 318874 58080
rect 319654 54707 325714 58080
rect 326494 54707 329434 58080
rect 330214 54707 333154 58080
rect 333934 54707 336874 58080
rect 337654 54707 343714 58080
rect 344494 54707 347434 58080
rect 348214 54707 351154 58080
rect 351934 54707 354874 58080
rect 355654 54707 361714 58080
rect 362494 54707 365434 518080
rect 366214 54707 369154 518080
rect 369934 54707 372874 518080
rect 373654 460228 379714 518080
rect 380494 460228 383434 518080
rect 384214 460228 387154 518080
rect 387934 460228 390874 518080
rect 391654 460228 397714 518080
rect 398494 460228 401434 518080
rect 402214 460228 405154 518080
rect 405934 460228 408874 518080
rect 409654 460228 415714 518080
rect 416494 460228 419434 518080
rect 420214 460228 423154 518080
rect 423934 460228 426874 518080
rect 427654 460228 433714 518080
rect 434494 460228 437434 630869
rect 438214 460228 441154 630869
rect 441934 460228 444874 630869
rect 445654 460228 451714 630869
rect 452494 460228 455434 630869
rect 456214 621920 459154 630869
rect 459934 621920 462874 630869
rect 463654 621920 469714 630869
rect 470494 621920 473434 630869
rect 474214 621920 477154 630869
rect 477934 621920 480874 630869
rect 481654 621920 487714 630869
rect 488494 621920 491434 630869
rect 492214 621920 495154 630869
rect 495934 621920 498874 630869
rect 499654 621920 505714 630869
rect 506494 621920 509434 630869
rect 510214 621920 513154 630869
rect 456214 568080 513154 621920
rect 456214 460228 459154 568080
rect 459934 460228 462874 568080
rect 463654 460228 469714 568080
rect 470494 460228 473434 568080
rect 474214 460228 477154 568080
rect 477934 460228 480874 568080
rect 481654 460228 487714 568080
rect 488494 460228 491434 568080
rect 492214 460228 495154 568080
rect 495934 460228 498874 568080
rect 499654 460228 505714 568080
rect 506494 460228 509434 568080
rect 510214 460228 513154 568080
rect 513934 460228 516496 630869
rect 373654 373080 516496 460228
rect 373654 355228 379714 373080
rect 380494 355228 383434 373080
rect 384214 355228 387154 373080
rect 387934 355228 390874 373080
rect 391654 355228 397714 373080
rect 398494 355228 401434 373080
rect 402214 355228 405154 373080
rect 405934 355228 408874 373080
rect 409654 355228 415714 373080
rect 416494 355228 419434 373080
rect 420214 355228 423154 373080
rect 423934 355228 426874 373080
rect 427654 355228 433714 373080
rect 434494 355228 437434 373080
rect 438214 355228 441154 373080
rect 441934 355228 444874 373080
rect 445654 355228 451714 373080
rect 452494 355228 455434 373080
rect 456214 355228 459154 373080
rect 459934 355228 462874 373080
rect 463654 355228 469714 373080
rect 470494 355228 473434 373080
rect 474214 355228 477154 373080
rect 477934 355228 480874 373080
rect 481654 355228 487714 373080
rect 488494 355228 491434 373080
rect 492214 355228 495154 373080
rect 495934 355228 498874 373080
rect 499654 355228 505714 373080
rect 506494 355228 509434 373080
rect 510214 355228 513154 373080
rect 513934 355228 516496 373080
rect 373654 268080 516496 355228
rect 373654 250228 379714 268080
rect 380494 250228 383434 268080
rect 384214 250228 387154 268080
rect 387934 250228 390874 268080
rect 391654 250228 397714 268080
rect 398494 250228 401434 268080
rect 402214 250228 405154 268080
rect 405934 250228 408874 268080
rect 409654 250228 415714 268080
rect 416494 250228 419434 268080
rect 420214 250228 423154 268080
rect 423934 250228 426874 268080
rect 427654 250228 433714 268080
rect 434494 250228 437434 268080
rect 438214 250228 441154 268080
rect 441934 250228 444874 268080
rect 445654 250228 451714 268080
rect 452494 250228 455434 268080
rect 456214 250228 459154 268080
rect 459934 250228 462874 268080
rect 463654 250228 469714 268080
rect 470494 250228 473434 268080
rect 474214 250228 477154 268080
rect 477934 250228 480874 268080
rect 481654 250228 487714 268080
rect 488494 250228 491434 268080
rect 492214 250228 495154 268080
rect 495934 250228 498874 268080
rect 499654 250228 505714 268080
rect 506494 250228 509434 268080
rect 510214 250228 513154 268080
rect 513934 250228 516496 268080
rect 373654 163080 516496 250228
rect 373654 145228 379714 163080
rect 380494 145228 383434 163080
rect 384214 145228 387154 163080
rect 387934 145228 390874 163080
rect 391654 145228 397714 163080
rect 398494 145228 401434 163080
rect 402214 145228 405154 163080
rect 405934 145228 408874 163080
rect 409654 145228 415714 163080
rect 416494 145228 419434 163080
rect 420214 145228 423154 163080
rect 423934 145228 426874 163080
rect 427654 145228 433714 163080
rect 434494 145228 437434 163080
rect 438214 145228 441154 163080
rect 441934 145228 444874 163080
rect 445654 145228 451714 163080
rect 452494 145228 455434 163080
rect 456214 145228 459154 163080
rect 459934 145228 462874 163080
rect 463654 145228 469714 163080
rect 470494 145228 473434 163080
rect 474214 145228 477154 163080
rect 477934 145228 480874 163080
rect 481654 145228 487714 163080
rect 488494 145228 491434 163080
rect 492214 145228 495154 163080
rect 495934 145228 498874 163080
rect 499654 145228 505714 163080
rect 506494 145228 509434 163080
rect 510214 145228 513154 163080
rect 513934 145228 516496 163080
rect 373654 58080 516496 145228
rect 373654 54707 379714 58080
rect 380494 54707 383434 58080
rect 384214 54707 387154 58080
rect 387934 54707 390874 58080
rect 391654 54707 397714 58080
rect 398494 54707 401434 58080
rect 402214 54707 405154 58080
rect 405934 54707 408874 58080
rect 409654 54707 415714 58080
rect 416494 54707 419434 58080
rect 420214 54707 423154 58080
rect 423934 54707 426874 58080
rect 427654 54707 433714 58080
rect 434494 54707 437434 58080
rect 438214 54707 441154 58080
rect 441934 54707 444874 58080
rect 445654 54707 451714 58080
rect 452494 54707 455434 58080
rect 456214 54707 459154 58080
rect 459934 54707 462874 58080
rect 463654 54707 469714 58080
rect 470494 54707 473434 58080
rect 474214 54707 477154 58080
rect 477934 54707 480874 58080
rect 481654 54707 487714 58080
rect 488494 54707 491434 58080
rect 492214 54707 495154 58080
rect 495934 54707 498874 58080
rect 499654 54707 505714 58080
rect 506494 54707 509434 58080
rect 510214 54707 513154 58080
rect 513934 54707 516496 58080
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -6806 694306 590730 694926
rect -4886 690586 588810 691206
rect -2966 686866 586890 687486
rect -8726 680026 592650 680646
rect -6806 676306 590730 676926
rect -4886 672586 588810 673206
rect -2966 668866 586890 669486
rect -8726 662026 592650 662646
rect -6806 658306 590730 658926
rect -4886 654586 588810 655206
rect -2966 650866 586890 651486
rect -8726 644026 592650 644646
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -2966 632866 586890 633486
rect -8726 626026 592650 626646
rect -6806 622306 590730 622926
rect -4886 618586 588810 619206
rect -2966 614866 586890 615486
rect -8726 608026 592650 608646
rect -6806 604306 590730 604926
rect -4886 600586 588810 601206
rect -2966 596866 586890 597486
rect -8726 590026 592650 590646
rect -6806 586306 590730 586926
rect -4886 582586 588810 583206
rect -2966 578866 586890 579486
rect -8726 572026 592650 572646
rect -6806 568306 590730 568926
rect -4886 564586 588810 565206
rect -2966 560866 586890 561486
rect -8726 554026 592650 554646
rect 66954 553086 283574 553706
rect -6806 550306 590730 550926
rect 63234 549366 279854 549986
rect 59514 547526 276134 548146
rect -4886 546586 588810 547206
rect 91794 543806 272414 544426
rect -2966 542866 586890 543486
rect -8726 536026 592650 536646
rect -6806 532306 590730 532926
rect -4886 528586 588810 529206
rect -2966 524866 586890 525486
rect -8726 518026 592650 518646
rect -6806 514306 590730 514926
rect -4886 510586 588810 511206
rect -2966 506866 586890 507486
rect -8726 500026 592650 500646
rect -6806 496306 590730 496926
rect -4886 492586 588810 493206
rect -2966 488866 586890 489486
rect -8726 482026 592650 482646
rect -6806 478306 590730 478926
rect -4886 474586 588810 475206
rect 59514 473646 276134 474266
rect -2966 470866 586890 471486
rect 91794 470110 272414 470546
rect 63234 469490 279854 470110
rect 81234 468550 297854 469170
rect 84954 464966 301574 465586
rect -8726 464026 592650 464646
rect -6806 460306 590730 460926
rect -4886 456586 588810 457206
rect -2966 452866 586890 453486
rect -8726 446026 592650 446646
rect -6806 442306 590730 442926
rect -4886 438586 588810 439206
rect -2966 434866 586890 435486
rect -8726 428026 592650 428646
rect -6806 424306 590730 424926
rect -4886 420586 588810 421206
rect -2966 416866 586890 417486
rect -8726 410026 592650 410646
rect -6806 406306 590730 406926
rect -4886 402586 588810 403206
rect -2966 398866 586890 399486
rect -8726 392026 592650 392646
rect -6806 388306 590730 388926
rect -4886 384586 588810 385206
rect -2966 380866 586890 381486
rect -8726 374026 592650 374646
rect -6806 370306 590730 370926
rect 63234 369366 495854 369986
rect -4886 366586 588810 367206
rect 59514 365646 492134 366266
rect 91794 363806 488414 364426
rect -2966 362866 586890 363486
rect 84954 356966 517574 357586
rect -8726 356026 592650 356646
rect -6806 352306 590730 352926
rect -4886 348586 588810 349206
rect -2966 344866 586890 345486
rect -8726 338026 592650 338646
rect -6806 334306 590730 334926
rect -4886 330586 588810 331206
rect -2966 326866 586890 327486
rect -8726 320026 592650 320646
rect -6806 316306 590730 316926
rect -4886 312586 588810 313206
rect -2966 308866 586890 309486
rect -8726 302026 592650 302646
rect -6806 298306 590730 298926
rect -4886 294586 588810 295206
rect -2966 290866 586890 291486
rect -8726 284026 592650 284646
rect -6806 280306 590730 280926
rect -4886 276586 588810 277206
rect -2966 272866 586890 273486
rect -8726 266026 592650 266646
rect 66954 265086 499574 265706
rect -6806 262306 590730 262926
rect 63234 261366 495854 261986
rect 59514 259526 492134 260146
rect -4886 258586 588810 259206
rect 91794 255806 488414 256426
rect -2966 254866 586890 255486
rect -8726 248026 592650 248646
rect -6806 244306 590730 244926
rect -4886 240586 588810 241206
rect -2966 236866 586890 237486
rect -8726 230026 592650 230646
rect -6806 226306 590730 226926
rect -4886 222586 588810 223206
rect -2966 218866 586890 219486
rect -8726 212026 592650 212646
rect -6806 208306 590730 208926
rect -4886 204586 588810 205206
rect -2966 200866 586890 201486
rect -8726 194026 592650 194646
rect -6806 190306 590730 190926
rect -4886 186586 588810 187206
rect -2966 182866 586890 183486
rect -8726 176026 592650 176646
rect -6806 172306 590730 172926
rect -4886 168586 588810 169206
rect -2966 164866 586890 165486
rect -8726 158026 592650 158646
rect 66954 157086 499574 157706
rect -6806 154306 590730 154926
rect 63234 153366 495854 153986
rect 59514 151526 492134 152146
rect -4886 150586 588810 151206
rect 91794 147806 488414 148426
rect -2966 146866 586890 147486
rect -8726 140026 592650 140646
rect -6806 136306 590730 136926
rect -4886 132586 588810 133206
rect -2966 128866 586890 129486
rect -8726 122026 592650 122646
rect -6806 118306 590730 118926
rect -4886 114586 588810 115206
rect -2966 110866 586890 111486
rect -8726 104026 592650 104646
rect -6806 100306 590730 100926
rect -4886 96586 588810 97206
rect -2966 92866 586890 93486
rect -8726 86026 592650 86646
rect -6806 82306 590730 82926
rect -4886 78586 588810 79206
rect -2966 74866 586890 75486
rect -8726 68026 592650 68646
rect -6806 64306 590730 64926
rect -4886 60586 588810 61206
rect -2966 56866 586890 57486
rect -8726 50026 592650 50646
rect -6806 46306 590730 46926
rect -4886 42586 588810 43206
rect -2966 38866 586890 39486
rect -8726 32026 592650 32646
rect -6806 28306 590730 28926
rect -4886 24586 588810 25206
rect -2966 20866 586890 21486
rect -8726 14026 592650 14646
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 145308 74414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 145308 110414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 145308 146414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 145308 182414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 145308 218414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 145308 254414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 145308 290414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 145308 326414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 145308 398414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 145308 434414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 145308 470414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 145308 506414 163000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 250308 74414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 250308 110414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 250308 146414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 250308 182414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 250308 218414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 250308 254414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 250308 290414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 250308 326414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 250308 398414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 250308 434414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 250308 470414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 250308 506414 268000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 355308 74414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 355308 110414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 355308 146414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 355308 182414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 355308 218414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 355308 254414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 355308 290414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 355308 326414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 355308 398414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 355308 434414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 355308 470414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 355308 506414 373000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 460308 74414 478000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 460308 110414 478000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 460308 146414 478000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 460308 182414 478000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 460308 218414 478000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 460308 254414 478000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 460308 290414 478000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 460308 326414 518000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 -1894 362414 518000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 460308 398414 518000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 542000 74414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 542000 110414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 542000 146414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 542000 182414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 542000 218414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 542000 254414 558000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 460308 470414 568000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 460308 506414 568000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 625099 74414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 625099 110414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 625099 146414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 625099 182414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 625099 218414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 625099 254414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 542000 290414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 633033 326414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 633033 362414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 633033 398414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 460308 434414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 622000 470414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 622000 506414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 533 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 145308 78134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 145308 114134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 145308 150134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 145308 186134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 145308 222134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 145308 258134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 145308 294134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 145308 330134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 401514 145308 402134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 437514 145308 438134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 473514 145308 474134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 145308 510134 163000 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 250308 78134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 250308 114134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 250308 150134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 250308 186134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 250308 222134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 250308 258134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 250308 294134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 250308 330134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 401514 250308 402134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 437514 250308 438134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 473514 250308 474134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 250308 510134 268000 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 355308 78134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 355308 114134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 355308 150134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 355308 186134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 355308 222134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 355308 258134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 355308 294134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 355308 330134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 401514 355308 402134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 437514 355308 438134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 473514 355308 474134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 355308 510134 373000 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 460308 78134 478000 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 460308 114134 478000 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 460308 150134 478000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 460308 186134 478000 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 460308 222134 478000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 460308 258134 478000 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 460308 294134 478000 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 460308 330134 518000 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 -3814 366134 518000 6 vccd2
port 533 nsew power input
rlabel metal4 s 401514 460308 402134 518000 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 542000 78134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 542000 114134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 542000 150134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 542000 186134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 542000 222134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 542000 258134 558000 6 vccd2
port 533 nsew power input
rlabel metal4 s 473514 460308 474134 568000 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 460308 510134 568000 6 vccd2
port 533 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 625099 78134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 625099 114134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 625099 150134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 625099 186134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 625099 222134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 625099 258134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 542000 294134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 633033 330134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 633033 366134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 401514 633033 402134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 437514 460308 438134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 473514 622000 474134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 622000 510134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 533 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 534 nsew power input
rlabel metal5 s 81234 468550 297854 469170 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 534 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 145308 81854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 145308 117854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 145308 153854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 145308 189854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 145308 225854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 145308 261854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 145308 297854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 145308 333854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 405234 145308 405854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 441234 145308 441854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 477234 145308 477854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 145308 513854 163000 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 250308 81854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 250308 117854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 250308 153854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 250308 189854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 250308 225854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 250308 261854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 250308 297854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 250308 333854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 405234 250308 405854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 441234 250308 441854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 477234 250308 477854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 250308 513854 268000 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 355308 81854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 355308 117854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 355308 153854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 355308 189854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 355308 225854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 355308 261854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 355308 297854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 355308 333854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 405234 355308 405854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 441234 355308 441854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 477234 355308 477854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 355308 513854 373000 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 460308 81854 478000 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 460308 117854 478000 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 460308 153854 478000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 460308 189854 478000 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 460308 225854 478000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 460308 261854 478000 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 460308 297854 478000 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 460308 333854 518000 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 -5734 369854 518000 6 vdda1
port 534 nsew power input
rlabel metal4 s 405234 460308 405854 518000 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 542000 81854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 542000 117854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 542000 153854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 542000 189854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 542000 225854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 542000 261854 558000 6 vdda1
port 534 nsew power input
rlabel metal4 s 477234 460308 477854 568000 6 vdda1
port 534 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 625099 81854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 625099 117854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 625099 153854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 625099 189854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 625099 225854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 625099 261854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 542000 297854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 633033 333854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 633033 369854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 405234 633033 405854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 441234 460308 441854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 477234 622000 477854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 460308 513854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 534 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 535 nsew power input
rlabel metal5 s 84954 356966 517574 357586 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 535 nsew power input
rlabel metal5 s 84954 464966 301574 465586 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 535 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 145308 85574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 145308 121574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 145308 157574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 145308 193574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 145308 229574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 145308 265574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 145308 301574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 145308 337574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 408954 145308 409574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 444954 145308 445574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 480954 145308 481574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 145308 517574 163000 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 250308 85574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 250308 121574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 250308 157574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 250308 193574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 250308 229574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 250308 265574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 250308 301574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 250308 337574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 408954 250308 409574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 444954 250308 445574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 480954 250308 481574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 250308 517574 268000 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 355308 85574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 355308 121574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 355308 157574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 355308 193574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 355308 229574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 355308 265574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 355308 301574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 355308 337574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 408954 355308 409574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 444954 355308 445574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 480954 355308 481574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 355308 517574 373000 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 460308 85574 478000 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 460308 121574 478000 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 460308 157574 478000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 460308 193574 478000 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 460308 229574 478000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 460308 265574 478000 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 460308 301574 478000 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 460308 337574 518000 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 -7654 373574 518000 6 vdda2
port 535 nsew power input
rlabel metal4 s 408954 460308 409574 518000 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 542000 85574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 542000 121574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 542000 157574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 542000 193574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 542000 229574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 542000 265574 558000 6 vdda2
port 535 nsew power input
rlabel metal4 s 480954 460308 481574 568000 6 vdda2
port 535 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 625099 85574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 625099 121574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 625099 157574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 625099 193574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 625099 229574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 625099 265574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 542000 301574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 633033 337574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 633033 373574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 408954 633033 409574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 444954 460308 445574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 480954 622000 481574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 460308 517574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 535 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 536 nsew ground input
rlabel metal5 s 63234 153366 495854 153986 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 536 nsew ground input
rlabel metal5 s 63234 261366 495854 261986 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 536 nsew ground input
rlabel metal5 s 63234 369366 495854 369986 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 536 nsew ground input
rlabel metal5 s 63234 469490 279854 470110 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 536 nsew ground input
rlabel metal5 s 63234 549366 279854 549986 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 145308 63854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 145308 99854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 145308 135854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 145308 171854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 145308 243854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 145308 279854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 315234 145308 315854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 145308 351854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 145308 387854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423234 145308 423854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 145308 459854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495234 145308 495854 163000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 250308 63854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 250308 99854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 250308 135854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 250308 171854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 250308 243854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 250308 279854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 315234 250308 315854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 250308 351854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 250308 387854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423234 250308 423854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 250308 459854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495234 250308 495854 268000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 355308 63854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 355308 99854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 355308 135854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 355308 171854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 355308 243854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 355308 279854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 315234 355308 315854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 355308 351854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 355308 387854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423234 355308 423854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 355308 459854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495234 355308 495854 373000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 460308 63854 478000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 460308 99854 478000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 460308 135854 478000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 460308 171854 478000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 207234 -5734 207854 478000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 460308 243854 478000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 460308 279854 478000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 460308 351854 518000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 460308 387854 518000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423234 460308 423854 518000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 542000 63854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 542000 99854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 542000 171854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 542000 243854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 542000 279854 558000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 460308 459854 568000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495234 460308 495854 568000 6 vssa1
port 536 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 625099 63854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 625099 99854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 542000 135854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 625099 171854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 207234 542000 207854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 625099 243854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 625099 279854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 315234 460308 315854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 633033 351854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 633033 387854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423234 633033 423854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 622000 459854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495234 622000 495854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 537 nsew ground input
rlabel metal5 s 66954 157086 499574 157706 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 537 nsew ground input
rlabel metal5 s 66954 265086 499574 265706 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 537 nsew ground input
rlabel metal5 s 66954 553086 283574 553706 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 145308 67574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 145308 103574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 145308 139574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 145308 175574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 145308 247574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 145308 283574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 145308 319574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 145308 355574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 145308 391574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 426954 145308 427574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 145308 463574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 498954 145308 499574 163000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 250308 67574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 250308 103574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 250308 139574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 250308 175574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 250308 247574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 250308 283574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 250308 319574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 250308 355574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 250308 391574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 426954 250308 427574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 250308 463574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 498954 250308 499574 268000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 355308 67574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 355308 103574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 355308 139574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 355308 175574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 355308 247574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 355308 283574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 355308 319574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 355308 355574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 355308 391574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 426954 355308 427574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 355308 463574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 498954 355308 499574 373000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 460308 67574 478000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 460308 103574 478000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 460308 139574 478000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 460308 175574 478000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 210954 -7654 211574 478000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 460308 247574 478000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 460308 283574 478000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 460308 319574 518000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 460308 355574 518000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 460308 391574 518000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 426954 460308 427574 518000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 542000 67574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 542000 103574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 542000 139574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 542000 175574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 542000 247574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 542000 283574 558000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 460308 463574 568000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 498954 460308 499574 568000 6 vssa2
port 537 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 625099 67574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 625099 103574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 625099 139574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 625099 175574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 210954 542000 211574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 625099 247574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 625099 283574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 633033 319574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 633033 355574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 633033 391574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 426954 633033 427574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 622000 463574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 498954 622000 499574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 538 nsew ground input
rlabel metal5 s 91794 147806 488414 148426 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 538 nsew ground input
rlabel metal5 s 91794 255806 488414 256426 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 538 nsew ground input
rlabel metal5 s 91794 363806 488414 364426 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 538 nsew ground input
rlabel metal5 s 91794 469926 272414 470546 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 538 nsew ground input
rlabel metal5 s 91794 543806 272414 544426 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 145308 92414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 145308 128414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 145308 164414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 145308 236414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 145308 272414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 307794 145308 308414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 145308 344414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 145308 380414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 415794 145308 416414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 145308 452414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 487794 145308 488414 163000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 250308 92414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 250308 128414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 250308 164414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 250308 236414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 250308 272414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 307794 250308 308414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 250308 344414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 250308 380414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 415794 250308 416414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 250308 452414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 487794 250308 488414 268000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 355308 92414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 355308 128414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 355308 164414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 355308 236414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 355308 272414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 307794 355308 308414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 355308 344414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 355308 380414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 415794 355308 416414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 355308 452414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 487794 355308 488414 373000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 460308 92414 478000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 460308 128414 478000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 460308 164414 478000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 199794 -1894 200414 478000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 460308 236414 478000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 460308 272414 478000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 460308 344414 518000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 460308 380414 518000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 415794 460308 416414 518000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 542000 92414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 542000 164414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 199794 542000 200414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 542000 236414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 542000 272414 558000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 487794 460308 488414 568000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 625099 92414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 542000 128414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 625099 164414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 199794 625099 200414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 625099 236414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 625099 272414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 307794 460308 308414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 633033 344414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 633033 380414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 415794 633033 416414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 460308 452414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 487794 622000 488414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 539 nsew ground input
rlabel metal5 s 59514 151526 492134 152146 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 539 nsew ground input
rlabel metal5 s 59514 259526 492134 260146 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 539 nsew ground input
rlabel metal5 s 59514 365646 492134 366266 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 539 nsew ground input
rlabel metal5 s 59514 473646 276134 474266 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 539 nsew ground input
rlabel metal5 s 59514 547526 276134 548146 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 145308 60134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 145308 96134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 145308 132134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 145308 168134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 145308 240134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 145308 276134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 311514 145308 312134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 145308 348134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 145308 384134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 419514 145308 420134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 145308 456134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491514 145308 492134 163000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 250308 60134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 250308 96134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 250308 132134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 250308 168134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 250308 240134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 250308 276134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 311514 250308 312134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 250308 348134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 250308 384134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 419514 250308 420134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 250308 456134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491514 250308 492134 268000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 355308 60134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 355308 96134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 355308 132134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 355308 168134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 355308 240134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 355308 276134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 311514 355308 312134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 355308 348134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 355308 384134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 419514 355308 420134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 355308 456134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491514 355308 492134 373000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 460308 60134 478000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 460308 96134 478000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 460308 132134 478000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 460308 168134 478000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 203514 -3814 204134 478000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 460308 240134 478000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 460308 276134 478000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 460308 348134 518000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 460308 384134 518000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 419514 460308 420134 518000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 542000 60134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 542000 96134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 542000 168134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 542000 240134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 542000 276134 558000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491514 460308 492134 568000 6 vssd2
port 539 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 625099 60134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 625099 96134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 542000 132134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 625099 168134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 203514 542000 204134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 625099 240134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 625099 276134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 311514 460308 312134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 633033 348134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 633033 384134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 419514 633033 420134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 460308 456134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491514 622000 492134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 97543972
string GDS_FILE /home/burak/asic_tools/caravel_vscpu3x/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 94134178
<< end >>

