VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO main_controller
  CLASS BLOCK ;
  FOREIGN main_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 735.000 ;
  PIN agent_1_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 445.440 600.000 446.040 ;
    END
  END agent_1_mem_ctrl_addr[0]
  PIN agent_1_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 472.640 600.000 473.240 ;
    END
  END agent_1_mem_ctrl_addr[10]
  PIN agent_1_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 475.360 600.000 475.960 ;
    END
  END agent_1_mem_ctrl_addr[11]
  PIN agent_1_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 478.080 600.000 478.680 ;
    END
  END agent_1_mem_ctrl_addr[12]
  PIN agent_1_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 480.800 600.000 481.400 ;
    END
  END agent_1_mem_ctrl_addr[13]
  PIN agent_1_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 448.160 600.000 448.760 ;
    END
  END agent_1_mem_ctrl_addr[1]
  PIN agent_1_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 450.880 600.000 451.480 ;
    END
  END agent_1_mem_ctrl_addr[2]
  PIN agent_1_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 453.600 600.000 454.200 ;
    END
  END agent_1_mem_ctrl_addr[3]
  PIN agent_1_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 456.320 600.000 456.920 ;
    END
  END agent_1_mem_ctrl_addr[4]
  PIN agent_1_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 459.040 600.000 459.640 ;
    END
  END agent_1_mem_ctrl_addr[5]
  PIN agent_1_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 461.760 600.000 462.360 ;
    END
  END agent_1_mem_ctrl_addr[6]
  PIN agent_1_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 464.480 600.000 465.080 ;
    END
  END agent_1_mem_ctrl_addr[7]
  PIN agent_1_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 467.200 600.000 467.800 ;
    END
  END agent_1_mem_ctrl_addr[8]
  PIN agent_1_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 469.920 600.000 470.520 ;
    END
  END agent_1_mem_ctrl_addr[9]
  PIN agent_1_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 483.520 600.000 484.120 ;
    END
  END agent_1_mem_ctrl_in[0]
  PIN agent_1_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 511.400 600.000 512.000 ;
    END
  END agent_1_mem_ctrl_in[10]
  PIN agent_1_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 514.120 600.000 514.720 ;
    END
  END agent_1_mem_ctrl_in[11]
  PIN agent_1_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 516.840 600.000 517.440 ;
    END
  END agent_1_mem_ctrl_in[12]
  PIN agent_1_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 519.560 600.000 520.160 ;
    END
  END agent_1_mem_ctrl_in[13]
  PIN agent_1_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 522.280 600.000 522.880 ;
    END
  END agent_1_mem_ctrl_in[14]
  PIN agent_1_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 525.000 600.000 525.600 ;
    END
  END agent_1_mem_ctrl_in[15]
  PIN agent_1_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 527.720 600.000 528.320 ;
    END
  END agent_1_mem_ctrl_in[16]
  PIN agent_1_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 530.440 600.000 531.040 ;
    END
  END agent_1_mem_ctrl_in[17]
  PIN agent_1_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 533.160 600.000 533.760 ;
    END
  END agent_1_mem_ctrl_in[18]
  PIN agent_1_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 535.880 600.000 536.480 ;
    END
  END agent_1_mem_ctrl_in[19]
  PIN agent_1_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 486.240 600.000 486.840 ;
    END
  END agent_1_mem_ctrl_in[1]
  PIN agent_1_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 538.600 600.000 539.200 ;
    END
  END agent_1_mem_ctrl_in[20]
  PIN agent_1_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 541.320 600.000 541.920 ;
    END
  END agent_1_mem_ctrl_in[21]
  PIN agent_1_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 544.040 600.000 544.640 ;
    END
  END agent_1_mem_ctrl_in[22]
  PIN agent_1_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 546.760 600.000 547.360 ;
    END
  END agent_1_mem_ctrl_in[23]
  PIN agent_1_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 549.480 600.000 550.080 ;
    END
  END agent_1_mem_ctrl_in[24]
  PIN agent_1_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 552.200 600.000 552.800 ;
    END
  END agent_1_mem_ctrl_in[25]
  PIN agent_1_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 554.920 600.000 555.520 ;
    END
  END agent_1_mem_ctrl_in[26]
  PIN agent_1_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 557.640 600.000 558.240 ;
    END
  END agent_1_mem_ctrl_in[27]
  PIN agent_1_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 560.360 600.000 560.960 ;
    END
  END agent_1_mem_ctrl_in[28]
  PIN agent_1_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 563.080 600.000 563.680 ;
    END
  END agent_1_mem_ctrl_in[29]
  PIN agent_1_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 488.960 600.000 489.560 ;
    END
  END agent_1_mem_ctrl_in[2]
  PIN agent_1_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 565.800 600.000 566.400 ;
    END
  END agent_1_mem_ctrl_in[30]
  PIN agent_1_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 568.520 600.000 569.120 ;
    END
  END agent_1_mem_ctrl_in[31]
  PIN agent_1_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 492.360 600.000 492.960 ;
    END
  END agent_1_mem_ctrl_in[3]
  PIN agent_1_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 495.080 600.000 495.680 ;
    END
  END agent_1_mem_ctrl_in[4]
  PIN agent_1_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 497.800 600.000 498.400 ;
    END
  END agent_1_mem_ctrl_in[5]
  PIN agent_1_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 500.520 600.000 501.120 ;
    END
  END agent_1_mem_ctrl_in[6]
  PIN agent_1_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 503.240 600.000 503.840 ;
    END
  END agent_1_mem_ctrl_in[7]
  PIN agent_1_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 505.960 600.000 506.560 ;
    END
  END agent_1_mem_ctrl_in[8]
  PIN agent_1_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 508.680 600.000 509.280 ;
    END
  END agent_1_mem_ctrl_in[9]
  PIN agent_1_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 571.240 600.000 571.840 ;
    END
  END agent_1_mem_ctrl_out[0]
  PIN agent_1_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 599.120 600.000 599.720 ;
    END
  END agent_1_mem_ctrl_out[10]
  PIN agent_1_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 601.840 600.000 602.440 ;
    END
  END agent_1_mem_ctrl_out[11]
  PIN agent_1_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 604.560 600.000 605.160 ;
    END
  END agent_1_mem_ctrl_out[12]
  PIN agent_1_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 607.280 600.000 607.880 ;
    END
  END agent_1_mem_ctrl_out[13]
  PIN agent_1_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 610.000 600.000 610.600 ;
    END
  END agent_1_mem_ctrl_out[14]
  PIN agent_1_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 612.720 600.000 613.320 ;
    END
  END agent_1_mem_ctrl_out[15]
  PIN agent_1_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 615.440 600.000 616.040 ;
    END
  END agent_1_mem_ctrl_out[16]
  PIN agent_1_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 618.160 600.000 618.760 ;
    END
  END agent_1_mem_ctrl_out[17]
  PIN agent_1_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 620.880 600.000 621.480 ;
    END
  END agent_1_mem_ctrl_out[18]
  PIN agent_1_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 623.600 600.000 624.200 ;
    END
  END agent_1_mem_ctrl_out[19]
  PIN agent_1_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 574.640 600.000 575.240 ;
    END
  END agent_1_mem_ctrl_out[1]
  PIN agent_1_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 626.320 600.000 626.920 ;
    END
  END agent_1_mem_ctrl_out[20]
  PIN agent_1_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 629.040 600.000 629.640 ;
    END
  END agent_1_mem_ctrl_out[21]
  PIN agent_1_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 631.760 600.000 632.360 ;
    END
  END agent_1_mem_ctrl_out[22]
  PIN agent_1_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 634.480 600.000 635.080 ;
    END
  END agent_1_mem_ctrl_out[23]
  PIN agent_1_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 637.200 600.000 637.800 ;
    END
  END agent_1_mem_ctrl_out[24]
  PIN agent_1_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 639.920 600.000 640.520 ;
    END
  END agent_1_mem_ctrl_out[25]
  PIN agent_1_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 642.640 600.000 643.240 ;
    END
  END agent_1_mem_ctrl_out[26]
  PIN agent_1_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 645.360 600.000 645.960 ;
    END
  END agent_1_mem_ctrl_out[27]
  PIN agent_1_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 648.080 600.000 648.680 ;
    END
  END agent_1_mem_ctrl_out[28]
  PIN agent_1_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 650.800 600.000 651.400 ;
    END
  END agent_1_mem_ctrl_out[29]
  PIN agent_1_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 577.360 600.000 577.960 ;
    END
  END agent_1_mem_ctrl_out[2]
  PIN agent_1_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 653.520 600.000 654.120 ;
    END
  END agent_1_mem_ctrl_out[30]
  PIN agent_1_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 656.920 600.000 657.520 ;
    END
  END agent_1_mem_ctrl_out[31]
  PIN agent_1_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 580.080 600.000 580.680 ;
    END
  END agent_1_mem_ctrl_out[3]
  PIN agent_1_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 582.800 600.000 583.400 ;
    END
  END agent_1_mem_ctrl_out[4]
  PIN agent_1_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 585.520 600.000 586.120 ;
    END
  END agent_1_mem_ctrl_out[5]
  PIN agent_1_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 588.240 600.000 588.840 ;
    END
  END agent_1_mem_ctrl_out[6]
  PIN agent_1_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 590.960 600.000 591.560 ;
    END
  END agent_1_mem_ctrl_out[7]
  PIN agent_1_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 593.680 600.000 594.280 ;
    END
  END agent_1_mem_ctrl_out[8]
  PIN agent_1_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 596.400 600.000 597.000 ;
    END
  END agent_1_mem_ctrl_out[9]
  PIN agent_1_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 659.640 600.000 660.240 ;
    END
  END agent_1_mem_ctrl_req
  PIN agent_1_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 662.360 600.000 662.960 ;
    END
  END agent_1_mem_ctrl_vld
  PIN agent_1_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 665.080 600.000 665.680 ;
    END
  END agent_1_mem_ctrl_we
  PIN agent_1_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END agent_1_sram0_csb0
  PIN agent_1_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END agent_1_sram0_dout0[0]
  PIN agent_1_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END agent_1_sram0_dout0[10]
  PIN agent_1_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END agent_1_sram0_dout0[11]
  PIN agent_1_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END agent_1_sram0_dout0[12]
  PIN agent_1_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END agent_1_sram0_dout0[13]
  PIN agent_1_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END agent_1_sram0_dout0[14]
  PIN agent_1_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END agent_1_sram0_dout0[15]
  PIN agent_1_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END agent_1_sram0_dout0[16]
  PIN agent_1_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END agent_1_sram0_dout0[17]
  PIN agent_1_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END agent_1_sram0_dout0[18]
  PIN agent_1_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END agent_1_sram0_dout0[19]
  PIN agent_1_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END agent_1_sram0_dout0[1]
  PIN agent_1_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END agent_1_sram0_dout0[20]
  PIN agent_1_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END agent_1_sram0_dout0[21]
  PIN agent_1_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END agent_1_sram0_dout0[22]
  PIN agent_1_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END agent_1_sram0_dout0[23]
  PIN agent_1_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END agent_1_sram0_dout0[24]
  PIN agent_1_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END agent_1_sram0_dout0[25]
  PIN agent_1_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END agent_1_sram0_dout0[26]
  PIN agent_1_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END agent_1_sram0_dout0[27]
  PIN agent_1_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END agent_1_sram0_dout0[28]
  PIN agent_1_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END agent_1_sram0_dout0[29]
  PIN agent_1_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END agent_1_sram0_dout0[2]
  PIN agent_1_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END agent_1_sram0_dout0[30]
  PIN agent_1_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END agent_1_sram0_dout0[31]
  PIN agent_1_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END agent_1_sram0_dout0[3]
  PIN agent_1_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END agent_1_sram0_dout0[4]
  PIN agent_1_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END agent_1_sram0_dout0[5]
  PIN agent_1_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END agent_1_sram0_dout0[6]
  PIN agent_1_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END agent_1_sram0_dout0[7]
  PIN agent_1_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END agent_1_sram0_dout0[8]
  PIN agent_1_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END agent_1_sram0_dout0[9]
  PIN agent_1_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END agent_1_sram0_web0
  PIN agent_1_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END agent_1_sram1_csb0
  PIN agent_1_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END agent_1_sram1_dout0[0]
  PIN agent_1_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END agent_1_sram1_dout0[10]
  PIN agent_1_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END agent_1_sram1_dout0[11]
  PIN agent_1_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END agent_1_sram1_dout0[12]
  PIN agent_1_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END agent_1_sram1_dout0[13]
  PIN agent_1_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END agent_1_sram1_dout0[14]
  PIN agent_1_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END agent_1_sram1_dout0[15]
  PIN agent_1_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END agent_1_sram1_dout0[16]
  PIN agent_1_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END agent_1_sram1_dout0[17]
  PIN agent_1_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END agent_1_sram1_dout0[18]
  PIN agent_1_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END agent_1_sram1_dout0[19]
  PIN agent_1_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END agent_1_sram1_dout0[1]
  PIN agent_1_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END agent_1_sram1_dout0[20]
  PIN agent_1_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END agent_1_sram1_dout0[21]
  PIN agent_1_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END agent_1_sram1_dout0[22]
  PIN agent_1_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END agent_1_sram1_dout0[23]
  PIN agent_1_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END agent_1_sram1_dout0[24]
  PIN agent_1_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END agent_1_sram1_dout0[25]
  PIN agent_1_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END agent_1_sram1_dout0[26]
  PIN agent_1_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END agent_1_sram1_dout0[27]
  PIN agent_1_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END agent_1_sram1_dout0[28]
  PIN agent_1_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END agent_1_sram1_dout0[29]
  PIN agent_1_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END agent_1_sram1_dout0[2]
  PIN agent_1_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END agent_1_sram1_dout0[30]
  PIN agent_1_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END agent_1_sram1_dout0[31]
  PIN agent_1_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END agent_1_sram1_dout0[3]
  PIN agent_1_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END agent_1_sram1_dout0[4]
  PIN agent_1_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END agent_1_sram1_dout0[5]
  PIN agent_1_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END agent_1_sram1_dout0[6]
  PIN agent_1_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END agent_1_sram1_dout0[7]
  PIN agent_1_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END agent_1_sram1_dout0[8]
  PIN agent_1_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END agent_1_sram1_dout0[9]
  PIN agent_1_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END agent_1_sram1_web0
  PIN agent_1_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END agent_1_sram2_csb0
  PIN agent_1_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 498.480 4.000 499.080 ;
    END
  END agent_1_sram2_dout0[0]
  PIN agent_1_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END agent_1_sram2_dout0[10]
  PIN agent_1_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END agent_1_sram2_dout0[11]
  PIN agent_1_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END agent_1_sram2_dout0[12]
  PIN agent_1_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END agent_1_sram2_dout0[13]
  PIN agent_1_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END agent_1_sram2_dout0[14]
  PIN agent_1_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END agent_1_sram2_dout0[15]
  PIN agent_1_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END agent_1_sram2_dout0[16]
  PIN agent_1_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END agent_1_sram2_dout0[17]
  PIN agent_1_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END agent_1_sram2_dout0[18]
  PIN agent_1_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END agent_1_sram2_dout0[19]
  PIN agent_1_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END agent_1_sram2_dout0[1]
  PIN agent_1_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END agent_1_sram2_dout0[20]
  PIN agent_1_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END agent_1_sram2_dout0[21]
  PIN agent_1_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END agent_1_sram2_dout0[22]
  PIN agent_1_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END agent_1_sram2_dout0[23]
  PIN agent_1_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END agent_1_sram2_dout0[24]
  PIN agent_1_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END agent_1_sram2_dout0[25]
  PIN agent_1_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END agent_1_sram2_dout0[26]
  PIN agent_1_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END agent_1_sram2_dout0[27]
  PIN agent_1_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END agent_1_sram2_dout0[28]
  PIN agent_1_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END agent_1_sram2_dout0[29]
  PIN agent_1_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END agent_1_sram2_dout0[2]
  PIN agent_1_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END agent_1_sram2_dout0[30]
  PIN agent_1_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END agent_1_sram2_dout0[31]
  PIN agent_1_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END agent_1_sram2_dout0[3]
  PIN agent_1_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END agent_1_sram2_dout0[4]
  PIN agent_1_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END agent_1_sram2_dout0[5]
  PIN agent_1_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END agent_1_sram2_dout0[6]
  PIN agent_1_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END agent_1_sram2_dout0[7]
  PIN agent_1_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END agent_1_sram2_dout0[8]
  PIN agent_1_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END agent_1_sram2_dout0[9]
  PIN agent_1_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END agent_1_sram2_web0
  PIN agent_1_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END agent_1_sram_comm_addr0[0]
  PIN agent_1_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END agent_1_sram_comm_addr0[1]
  PIN agent_1_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END agent_1_sram_comm_addr0[2]
  PIN agent_1_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.080 4.000 614.680 ;
    END
  END agent_1_sram_comm_addr0[3]
  PIN agent_1_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END agent_1_sram_comm_addr0[4]
  PIN agent_1_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.880 4.000 621.480 ;
    END
  END agent_1_sram_comm_addr0[5]
  PIN agent_1_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END agent_1_sram_comm_addr0[6]
  PIN agent_1_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END agent_1_sram_comm_addr0[7]
  PIN agent_1_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END agent_1_sram_comm_addr0[8]
  PIN agent_1_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END agent_1_sram_comm_din0[0]
  PIN agent_1_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.760 4.000 666.360 ;
    END
  END agent_1_sram_comm_din0[10]
  PIN agent_1_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END agent_1_sram_comm_din0[11]
  PIN agent_1_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END agent_1_sram_comm_din0[12]
  PIN agent_1_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.280 4.000 675.880 ;
    END
  END agent_1_sram_comm_din0[13]
  PIN agent_1_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END agent_1_sram_comm_din0[14]
  PIN agent_1_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END agent_1_sram_comm_din0[15]
  PIN agent_1_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END agent_1_sram_comm_din0[16]
  PIN agent_1_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END agent_1_sram_comm_din0[17]
  PIN agent_1_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END agent_1_sram_comm_din0[18]
  PIN agent_1_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 694.320 4.000 694.920 ;
    END
  END agent_1_sram_comm_din0[19]
  PIN agent_1_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END agent_1_sram_comm_din0[1]
  PIN agent_1_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END agent_1_sram_comm_din0[20]
  PIN agent_1_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.120 4.000 701.720 ;
    END
  END agent_1_sram_comm_din0[21]
  PIN agent_1_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END agent_1_sram_comm_din0[22]
  PIN agent_1_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END agent_1_sram_comm_din0[23]
  PIN agent_1_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END agent_1_sram_comm_din0[24]
  PIN agent_1_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 713.360 4.000 713.960 ;
    END
  END agent_1_sram_comm_din0[25]
  PIN agent_1_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END agent_1_sram_comm_din0[26]
  PIN agent_1_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END agent_1_sram_comm_din0[27]
  PIN agent_1_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 723.560 4.000 724.160 ;
    END
  END agent_1_sram_comm_din0[28]
  PIN agent_1_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END agent_1_sram_comm_din0[29]
  PIN agent_1_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END agent_1_sram_comm_din0[2]
  PIN agent_1_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END agent_1_sram_comm_din0[30]
  PIN agent_1_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END agent_1_sram_comm_din0[31]
  PIN agent_1_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END agent_1_sram_comm_din0[3]
  PIN agent_1_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END agent_1_sram_comm_din0[4]
  PIN agent_1_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END agent_1_sram_comm_din0[5]
  PIN agent_1_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END agent_1_sram_comm_din0[6]
  PIN agent_1_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END agent_1_sram_comm_din0[7]
  PIN agent_1_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 4.000 659.560 ;
    END
  END agent_1_sram_comm_din0[8]
  PIN agent_1_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END agent_1_sram_comm_din0[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END clk
  PIN cm_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 1.400 600.000 2.000 ;
    END
  END cm_mem_ctrl_addr[0]
  PIN cm_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 28.600 600.000 29.200 ;
    END
  END cm_mem_ctrl_addr[10]
  PIN cm_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 31.320 600.000 31.920 ;
    END
  END cm_mem_ctrl_addr[11]
  PIN cm_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 34.040 600.000 34.640 ;
    END
  END cm_mem_ctrl_addr[12]
  PIN cm_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 36.760 600.000 37.360 ;
    END
  END cm_mem_ctrl_addr[13]
  PIN cm_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 4.120 600.000 4.720 ;
    END
  END cm_mem_ctrl_addr[1]
  PIN cm_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 6.840 600.000 7.440 ;
    END
  END cm_mem_ctrl_addr[2]
  PIN cm_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 9.560 600.000 10.160 ;
    END
  END cm_mem_ctrl_addr[3]
  PIN cm_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 12.280 600.000 12.880 ;
    END
  END cm_mem_ctrl_addr[4]
  PIN cm_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 15.000 600.000 15.600 ;
    END
  END cm_mem_ctrl_addr[5]
  PIN cm_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 17.720 600.000 18.320 ;
    END
  END cm_mem_ctrl_addr[6]
  PIN cm_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 20.440 600.000 21.040 ;
    END
  END cm_mem_ctrl_addr[7]
  PIN cm_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 23.160 600.000 23.760 ;
    END
  END cm_mem_ctrl_addr[8]
  PIN cm_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 25.880 600.000 26.480 ;
    END
  END cm_mem_ctrl_addr[9]
  PIN cm_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 39.480 600.000 40.080 ;
    END
  END cm_mem_ctrl_in[0]
  PIN cm_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 66.680 600.000 67.280 ;
    END
  END cm_mem_ctrl_in[10]
  PIN cm_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 69.400 600.000 70.000 ;
    END
  END cm_mem_ctrl_in[11]
  PIN cm_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 72.120 600.000 72.720 ;
    END
  END cm_mem_ctrl_in[12]
  PIN cm_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 74.840 600.000 75.440 ;
    END
  END cm_mem_ctrl_in[13]
  PIN cm_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 77.560 600.000 78.160 ;
    END
  END cm_mem_ctrl_in[14]
  PIN cm_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 80.280 600.000 80.880 ;
    END
  END cm_mem_ctrl_in[15]
  PIN cm_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 83.680 600.000 84.280 ;
    END
  END cm_mem_ctrl_in[16]
  PIN cm_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 86.400 600.000 87.000 ;
    END
  END cm_mem_ctrl_in[17]
  PIN cm_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 89.120 600.000 89.720 ;
    END
  END cm_mem_ctrl_in[18]
  PIN cm_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 91.840 600.000 92.440 ;
    END
  END cm_mem_ctrl_in[19]
  PIN cm_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 42.200 600.000 42.800 ;
    END
  END cm_mem_ctrl_in[1]
  PIN cm_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 94.560 600.000 95.160 ;
    END
  END cm_mem_ctrl_in[20]
  PIN cm_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 97.280 600.000 97.880 ;
    END
  END cm_mem_ctrl_in[21]
  PIN cm_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 100.000 600.000 100.600 ;
    END
  END cm_mem_ctrl_in[22]
  PIN cm_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 102.720 600.000 103.320 ;
    END
  END cm_mem_ctrl_in[23]
  PIN cm_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 105.440 600.000 106.040 ;
    END
  END cm_mem_ctrl_in[24]
  PIN cm_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 108.160 600.000 108.760 ;
    END
  END cm_mem_ctrl_in[25]
  PIN cm_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 110.880 600.000 111.480 ;
    END
  END cm_mem_ctrl_in[26]
  PIN cm_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 113.600 600.000 114.200 ;
    END
  END cm_mem_ctrl_in[27]
  PIN cm_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 116.320 600.000 116.920 ;
    END
  END cm_mem_ctrl_in[28]
  PIN cm_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 119.040 600.000 119.640 ;
    END
  END cm_mem_ctrl_in[29]
  PIN cm_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 44.920 600.000 45.520 ;
    END
  END cm_mem_ctrl_in[2]
  PIN cm_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 121.760 600.000 122.360 ;
    END
  END cm_mem_ctrl_in[30]
  PIN cm_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 124.480 600.000 125.080 ;
    END
  END cm_mem_ctrl_in[31]
  PIN cm_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 47.640 600.000 48.240 ;
    END
  END cm_mem_ctrl_in[3]
  PIN cm_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 50.360 600.000 50.960 ;
    END
  END cm_mem_ctrl_in[4]
  PIN cm_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 53.080 600.000 53.680 ;
    END
  END cm_mem_ctrl_in[5]
  PIN cm_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 55.800 600.000 56.400 ;
    END
  END cm_mem_ctrl_in[6]
  PIN cm_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 58.520 600.000 59.120 ;
    END
  END cm_mem_ctrl_in[7]
  PIN cm_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 61.240 600.000 61.840 ;
    END
  END cm_mem_ctrl_in[8]
  PIN cm_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 63.960 600.000 64.560 ;
    END
  END cm_mem_ctrl_in[9]
  PIN cm_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 127.200 600.000 127.800 ;
    END
  END cm_mem_ctrl_out[0]
  PIN cm_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 154.400 600.000 155.000 ;
    END
  END cm_mem_ctrl_out[10]
  PIN cm_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 157.120 600.000 157.720 ;
    END
  END cm_mem_ctrl_out[11]
  PIN cm_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 159.840 600.000 160.440 ;
    END
  END cm_mem_ctrl_out[12]
  PIN cm_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 162.560 600.000 163.160 ;
    END
  END cm_mem_ctrl_out[13]
  PIN cm_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 165.960 600.000 166.560 ;
    END
  END cm_mem_ctrl_out[14]
  PIN cm_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 168.680 600.000 169.280 ;
    END
  END cm_mem_ctrl_out[15]
  PIN cm_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 171.400 600.000 172.000 ;
    END
  END cm_mem_ctrl_out[16]
  PIN cm_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 174.120 600.000 174.720 ;
    END
  END cm_mem_ctrl_out[17]
  PIN cm_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 176.840 600.000 177.440 ;
    END
  END cm_mem_ctrl_out[18]
  PIN cm_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 179.560 600.000 180.160 ;
    END
  END cm_mem_ctrl_out[19]
  PIN cm_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 129.920 600.000 130.520 ;
    END
  END cm_mem_ctrl_out[1]
  PIN cm_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 182.280 600.000 182.880 ;
    END
  END cm_mem_ctrl_out[20]
  PIN cm_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 185.000 600.000 185.600 ;
    END
  END cm_mem_ctrl_out[21]
  PIN cm_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 187.720 600.000 188.320 ;
    END
  END cm_mem_ctrl_out[22]
  PIN cm_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 190.440 600.000 191.040 ;
    END
  END cm_mem_ctrl_out[23]
  PIN cm_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 193.160 600.000 193.760 ;
    END
  END cm_mem_ctrl_out[24]
  PIN cm_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 195.880 600.000 196.480 ;
    END
  END cm_mem_ctrl_out[25]
  PIN cm_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 198.600 600.000 199.200 ;
    END
  END cm_mem_ctrl_out[26]
  PIN cm_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 201.320 600.000 201.920 ;
    END
  END cm_mem_ctrl_out[27]
  PIN cm_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 204.040 600.000 204.640 ;
    END
  END cm_mem_ctrl_out[28]
  PIN cm_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 206.760 600.000 207.360 ;
    END
  END cm_mem_ctrl_out[29]
  PIN cm_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 132.640 600.000 133.240 ;
    END
  END cm_mem_ctrl_out[2]
  PIN cm_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 209.480 600.000 210.080 ;
    END
  END cm_mem_ctrl_out[30]
  PIN cm_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 212.200 600.000 212.800 ;
    END
  END cm_mem_ctrl_out[31]
  PIN cm_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 135.360 600.000 135.960 ;
    END
  END cm_mem_ctrl_out[3]
  PIN cm_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 138.080 600.000 138.680 ;
    END
  END cm_mem_ctrl_out[4]
  PIN cm_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 140.800 600.000 141.400 ;
    END
  END cm_mem_ctrl_out[5]
  PIN cm_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 143.520 600.000 144.120 ;
    END
  END cm_mem_ctrl_out[6]
  PIN cm_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 146.240 600.000 146.840 ;
    END
  END cm_mem_ctrl_out[7]
  PIN cm_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 148.960 600.000 149.560 ;
    END
  END cm_mem_ctrl_out[8]
  PIN cm_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 151.680 600.000 152.280 ;
    END
  END cm_mem_ctrl_out[9]
  PIN cm_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 214.920 600.000 215.520 ;
    END
  END cm_mem_ctrl_req
  PIN cm_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 217.640 600.000 218.240 ;
    END
  END cm_mem_ctrl_vld
  PIN cm_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 220.360 600.000 220.960 ;
    END
  END cm_mem_ctrl_we
  PIN cm_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END cm_sram0_csb0
  PIN cm_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END cm_sram0_dout0[0]
  PIN cm_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END cm_sram0_dout0[10]
  PIN cm_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END cm_sram0_dout0[11]
  PIN cm_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END cm_sram0_dout0[12]
  PIN cm_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END cm_sram0_dout0[13]
  PIN cm_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END cm_sram0_dout0[14]
  PIN cm_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END cm_sram0_dout0[15]
  PIN cm_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END cm_sram0_dout0[16]
  PIN cm_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END cm_sram0_dout0[17]
  PIN cm_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END cm_sram0_dout0[18]
  PIN cm_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END cm_sram0_dout0[19]
  PIN cm_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END cm_sram0_dout0[1]
  PIN cm_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END cm_sram0_dout0[20]
  PIN cm_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END cm_sram0_dout0[21]
  PIN cm_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END cm_sram0_dout0[22]
  PIN cm_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END cm_sram0_dout0[23]
  PIN cm_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END cm_sram0_dout0[24]
  PIN cm_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END cm_sram0_dout0[25]
  PIN cm_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END cm_sram0_dout0[26]
  PIN cm_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END cm_sram0_dout0[27]
  PIN cm_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END cm_sram0_dout0[28]
  PIN cm_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END cm_sram0_dout0[29]
  PIN cm_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END cm_sram0_dout0[2]
  PIN cm_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END cm_sram0_dout0[30]
  PIN cm_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END cm_sram0_dout0[31]
  PIN cm_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END cm_sram0_dout0[3]
  PIN cm_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END cm_sram0_dout0[4]
  PIN cm_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END cm_sram0_dout0[5]
  PIN cm_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END cm_sram0_dout0[6]
  PIN cm_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END cm_sram0_dout0[7]
  PIN cm_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END cm_sram0_dout0[8]
  PIN cm_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END cm_sram0_dout0[9]
  PIN cm_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END cm_sram0_web0
  PIN cm_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END cm_sram1_csb0
  PIN cm_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END cm_sram1_dout0[0]
  PIN cm_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END cm_sram1_dout0[10]
  PIN cm_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END cm_sram1_dout0[11]
  PIN cm_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END cm_sram1_dout0[12]
  PIN cm_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END cm_sram1_dout0[13]
  PIN cm_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END cm_sram1_dout0[14]
  PIN cm_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END cm_sram1_dout0[15]
  PIN cm_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END cm_sram1_dout0[16]
  PIN cm_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END cm_sram1_dout0[17]
  PIN cm_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END cm_sram1_dout0[18]
  PIN cm_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END cm_sram1_dout0[19]
  PIN cm_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END cm_sram1_dout0[1]
  PIN cm_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END cm_sram1_dout0[20]
  PIN cm_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END cm_sram1_dout0[21]
  PIN cm_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END cm_sram1_dout0[22]
  PIN cm_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END cm_sram1_dout0[23]
  PIN cm_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END cm_sram1_dout0[24]
  PIN cm_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END cm_sram1_dout0[25]
  PIN cm_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END cm_sram1_dout0[26]
  PIN cm_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END cm_sram1_dout0[27]
  PIN cm_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END cm_sram1_dout0[28]
  PIN cm_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END cm_sram1_dout0[29]
  PIN cm_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END cm_sram1_dout0[2]
  PIN cm_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END cm_sram1_dout0[30]
  PIN cm_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END cm_sram1_dout0[31]
  PIN cm_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END cm_sram1_dout0[3]
  PIN cm_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END cm_sram1_dout0[4]
  PIN cm_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END cm_sram1_dout0[5]
  PIN cm_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END cm_sram1_dout0[6]
  PIN cm_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END cm_sram1_dout0[7]
  PIN cm_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END cm_sram1_dout0[8]
  PIN cm_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END cm_sram1_dout0[9]
  PIN cm_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END cm_sram1_web0
  PIN cm_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END cm_sram2_csb0
  PIN cm_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END cm_sram2_dout0[0]
  PIN cm_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END cm_sram2_dout0[10]
  PIN cm_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END cm_sram2_dout0[11]
  PIN cm_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END cm_sram2_dout0[12]
  PIN cm_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END cm_sram2_dout0[13]
  PIN cm_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END cm_sram2_dout0[14]
  PIN cm_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END cm_sram2_dout0[15]
  PIN cm_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END cm_sram2_dout0[16]
  PIN cm_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END cm_sram2_dout0[17]
  PIN cm_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END cm_sram2_dout0[18]
  PIN cm_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END cm_sram2_dout0[19]
  PIN cm_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END cm_sram2_dout0[1]
  PIN cm_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END cm_sram2_dout0[20]
  PIN cm_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END cm_sram2_dout0[21]
  PIN cm_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END cm_sram2_dout0[22]
  PIN cm_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END cm_sram2_dout0[23]
  PIN cm_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END cm_sram2_dout0[24]
  PIN cm_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END cm_sram2_dout0[25]
  PIN cm_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END cm_sram2_dout0[26]
  PIN cm_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END cm_sram2_dout0[27]
  PIN cm_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END cm_sram2_dout0[28]
  PIN cm_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END cm_sram2_dout0[29]
  PIN cm_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END cm_sram2_dout0[2]
  PIN cm_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END cm_sram2_dout0[30]
  PIN cm_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END cm_sram2_dout0[31]
  PIN cm_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END cm_sram2_dout0[3]
  PIN cm_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END cm_sram2_dout0[4]
  PIN cm_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END cm_sram2_dout0[5]
  PIN cm_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END cm_sram2_dout0[6]
  PIN cm_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END cm_sram2_dout0[7]
  PIN cm_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END cm_sram2_dout0[8]
  PIN cm_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END cm_sram2_dout0[9]
  PIN cm_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END cm_sram2_web0
  PIN cm_sram3_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END cm_sram3_csb0
  PIN cm_sram3_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END cm_sram3_dout0[0]
  PIN cm_sram3_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END cm_sram3_dout0[10]
  PIN cm_sram3_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END cm_sram3_dout0[11]
  PIN cm_sram3_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END cm_sram3_dout0[12]
  PIN cm_sram3_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END cm_sram3_dout0[13]
  PIN cm_sram3_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END cm_sram3_dout0[14]
  PIN cm_sram3_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END cm_sram3_dout0[15]
  PIN cm_sram3_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END cm_sram3_dout0[16]
  PIN cm_sram3_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END cm_sram3_dout0[17]
  PIN cm_sram3_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END cm_sram3_dout0[18]
  PIN cm_sram3_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END cm_sram3_dout0[19]
  PIN cm_sram3_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END cm_sram3_dout0[1]
  PIN cm_sram3_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END cm_sram3_dout0[20]
  PIN cm_sram3_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END cm_sram3_dout0[21]
  PIN cm_sram3_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END cm_sram3_dout0[22]
  PIN cm_sram3_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END cm_sram3_dout0[23]
  PIN cm_sram3_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END cm_sram3_dout0[24]
  PIN cm_sram3_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END cm_sram3_dout0[25]
  PIN cm_sram3_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END cm_sram3_dout0[26]
  PIN cm_sram3_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END cm_sram3_dout0[27]
  PIN cm_sram3_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END cm_sram3_dout0[28]
  PIN cm_sram3_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END cm_sram3_dout0[29]
  PIN cm_sram3_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END cm_sram3_dout0[2]
  PIN cm_sram3_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END cm_sram3_dout0[30]
  PIN cm_sram3_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END cm_sram3_dout0[31]
  PIN cm_sram3_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END cm_sram3_dout0[3]
  PIN cm_sram3_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END cm_sram3_dout0[4]
  PIN cm_sram3_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END cm_sram3_dout0[5]
  PIN cm_sram3_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END cm_sram3_dout0[6]
  PIN cm_sram3_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END cm_sram3_dout0[7]
  PIN cm_sram3_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END cm_sram3_dout0[8]
  PIN cm_sram3_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END cm_sram3_dout0[9]
  PIN cm_sram3_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END cm_sram3_web0
  PIN cm_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END cm_sram_comm_addr0[0]
  PIN cm_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END cm_sram_comm_addr0[1]
  PIN cm_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END cm_sram_comm_addr0[2]
  PIN cm_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END cm_sram_comm_addr0[3]
  PIN cm_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END cm_sram_comm_addr0[4]
  PIN cm_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END cm_sram_comm_addr0[5]
  PIN cm_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 4.000 ;
    END
  END cm_sram_comm_addr0[6]
  PIN cm_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END cm_sram_comm_addr0[7]
  PIN cm_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END cm_sram_comm_addr0[8]
  PIN cm_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END cm_sram_comm_din0[0]
  PIN cm_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END cm_sram_comm_din0[10]
  PIN cm_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END cm_sram_comm_din0[11]
  PIN cm_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END cm_sram_comm_din0[12]
  PIN cm_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END cm_sram_comm_din0[13]
  PIN cm_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END cm_sram_comm_din0[14]
  PIN cm_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END cm_sram_comm_din0[15]
  PIN cm_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END cm_sram_comm_din0[16]
  PIN cm_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END cm_sram_comm_din0[17]
  PIN cm_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END cm_sram_comm_din0[18]
  PIN cm_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END cm_sram_comm_din0[19]
  PIN cm_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END cm_sram_comm_din0[1]
  PIN cm_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END cm_sram_comm_din0[20]
  PIN cm_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END cm_sram_comm_din0[21]
  PIN cm_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END cm_sram_comm_din0[22]
  PIN cm_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END cm_sram_comm_din0[23]
  PIN cm_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END cm_sram_comm_din0[24]
  PIN cm_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END cm_sram_comm_din0[25]
  PIN cm_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END cm_sram_comm_din0[26]
  PIN cm_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END cm_sram_comm_din0[27]
  PIN cm_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END cm_sram_comm_din0[28]
  PIN cm_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END cm_sram_comm_din0[29]
  PIN cm_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END cm_sram_comm_din0[2]
  PIN cm_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END cm_sram_comm_din0[30]
  PIN cm_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END cm_sram_comm_din0[31]
  PIN cm_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END cm_sram_comm_din0[3]
  PIN cm_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END cm_sram_comm_din0[4]
  PIN cm_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END cm_sram_comm_din0[5]
  PIN cm_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END cm_sram_comm_din0[6]
  PIN cm_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END cm_sram_comm_din0[7]
  PIN cm_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END cm_sram_comm_din0[8]
  PIN cm_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END cm_sram_comm_din0[9]
  PIN ct_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 223.080 600.000 223.680 ;
    END
  END ct_mem_ctrl_addr[0]
  PIN ct_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 250.960 600.000 251.560 ;
    END
  END ct_mem_ctrl_addr[10]
  PIN ct_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 253.680 600.000 254.280 ;
    END
  END ct_mem_ctrl_addr[11]
  PIN ct_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 256.400 600.000 257.000 ;
    END
  END ct_mem_ctrl_addr[12]
  PIN ct_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 259.120 600.000 259.720 ;
    END
  END ct_mem_ctrl_addr[13]
  PIN ct_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 225.800 600.000 226.400 ;
    END
  END ct_mem_ctrl_addr[1]
  PIN ct_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 228.520 600.000 229.120 ;
    END
  END ct_mem_ctrl_addr[2]
  PIN ct_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 231.240 600.000 231.840 ;
    END
  END ct_mem_ctrl_addr[3]
  PIN ct_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 233.960 600.000 234.560 ;
    END
  END ct_mem_ctrl_addr[4]
  PIN ct_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 236.680 600.000 237.280 ;
    END
  END ct_mem_ctrl_addr[5]
  PIN ct_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 239.400 600.000 240.000 ;
    END
  END ct_mem_ctrl_addr[6]
  PIN ct_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 242.120 600.000 242.720 ;
    END
  END ct_mem_ctrl_addr[7]
  PIN ct_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 244.840 600.000 245.440 ;
    END
  END ct_mem_ctrl_addr[8]
  PIN ct_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 248.240 600.000 248.840 ;
    END
  END ct_mem_ctrl_addr[9]
  PIN ct_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 261.840 600.000 262.440 ;
    END
  END ct_mem_ctrl_in[0]
  PIN ct_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 289.040 600.000 289.640 ;
    END
  END ct_mem_ctrl_in[10]
  PIN ct_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 291.760 600.000 292.360 ;
    END
  END ct_mem_ctrl_in[11]
  PIN ct_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 294.480 600.000 295.080 ;
    END
  END ct_mem_ctrl_in[12]
  PIN ct_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 297.200 600.000 297.800 ;
    END
  END ct_mem_ctrl_in[13]
  PIN ct_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 299.920 600.000 300.520 ;
    END
  END ct_mem_ctrl_in[14]
  PIN ct_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 302.640 600.000 303.240 ;
    END
  END ct_mem_ctrl_in[15]
  PIN ct_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 305.360 600.000 305.960 ;
    END
  END ct_mem_ctrl_in[16]
  PIN ct_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 308.080 600.000 308.680 ;
    END
  END ct_mem_ctrl_in[17]
  PIN ct_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 310.800 600.000 311.400 ;
    END
  END ct_mem_ctrl_in[18]
  PIN ct_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 313.520 600.000 314.120 ;
    END
  END ct_mem_ctrl_in[19]
  PIN ct_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 264.560 600.000 265.160 ;
    END
  END ct_mem_ctrl_in[1]
  PIN ct_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 316.240 600.000 316.840 ;
    END
  END ct_mem_ctrl_in[20]
  PIN ct_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 318.960 600.000 319.560 ;
    END
  END ct_mem_ctrl_in[21]
  PIN ct_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 321.680 600.000 322.280 ;
    END
  END ct_mem_ctrl_in[22]
  PIN ct_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 324.400 600.000 325.000 ;
    END
  END ct_mem_ctrl_in[23]
  PIN ct_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 327.120 600.000 327.720 ;
    END
  END ct_mem_ctrl_in[24]
  PIN ct_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 330.520 600.000 331.120 ;
    END
  END ct_mem_ctrl_in[25]
  PIN ct_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 333.240 600.000 333.840 ;
    END
  END ct_mem_ctrl_in[26]
  PIN ct_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 335.960 600.000 336.560 ;
    END
  END ct_mem_ctrl_in[27]
  PIN ct_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 338.680 600.000 339.280 ;
    END
  END ct_mem_ctrl_in[28]
  PIN ct_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 341.400 600.000 342.000 ;
    END
  END ct_mem_ctrl_in[29]
  PIN ct_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 267.280 600.000 267.880 ;
    END
  END ct_mem_ctrl_in[2]
  PIN ct_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 344.120 600.000 344.720 ;
    END
  END ct_mem_ctrl_in[30]
  PIN ct_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 346.840 600.000 347.440 ;
    END
  END ct_mem_ctrl_in[31]
  PIN ct_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 270.000 600.000 270.600 ;
    END
  END ct_mem_ctrl_in[3]
  PIN ct_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 272.720 600.000 273.320 ;
    END
  END ct_mem_ctrl_in[4]
  PIN ct_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 275.440 600.000 276.040 ;
    END
  END ct_mem_ctrl_in[5]
  PIN ct_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 278.160 600.000 278.760 ;
    END
  END ct_mem_ctrl_in[6]
  PIN ct_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 280.880 600.000 281.480 ;
    END
  END ct_mem_ctrl_in[7]
  PIN ct_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 283.600 600.000 284.200 ;
    END
  END ct_mem_ctrl_in[8]
  PIN ct_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 286.320 600.000 286.920 ;
    END
  END ct_mem_ctrl_in[9]
  PIN ct_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 349.560 600.000 350.160 ;
    END
  END ct_mem_ctrl_out[0]
  PIN ct_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 376.760 600.000 377.360 ;
    END
  END ct_mem_ctrl_out[10]
  PIN ct_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 379.480 600.000 380.080 ;
    END
  END ct_mem_ctrl_out[11]
  PIN ct_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 382.200 600.000 382.800 ;
    END
  END ct_mem_ctrl_out[12]
  PIN ct_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 384.920 600.000 385.520 ;
    END
  END ct_mem_ctrl_out[13]
  PIN ct_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 387.640 600.000 388.240 ;
    END
  END ct_mem_ctrl_out[14]
  PIN ct_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 390.360 600.000 390.960 ;
    END
  END ct_mem_ctrl_out[15]
  PIN ct_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 393.080 600.000 393.680 ;
    END
  END ct_mem_ctrl_out[16]
  PIN ct_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 395.800 600.000 396.400 ;
    END
  END ct_mem_ctrl_out[17]
  PIN ct_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 398.520 600.000 399.120 ;
    END
  END ct_mem_ctrl_out[18]
  PIN ct_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 401.240 600.000 401.840 ;
    END
  END ct_mem_ctrl_out[19]
  PIN ct_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 352.280 600.000 352.880 ;
    END
  END ct_mem_ctrl_out[1]
  PIN ct_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 403.960 600.000 404.560 ;
    END
  END ct_mem_ctrl_out[20]
  PIN ct_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 406.680 600.000 407.280 ;
    END
  END ct_mem_ctrl_out[21]
  PIN ct_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 410.080 600.000 410.680 ;
    END
  END ct_mem_ctrl_out[22]
  PIN ct_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 412.800 600.000 413.400 ;
    END
  END ct_mem_ctrl_out[23]
  PIN ct_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 415.520 600.000 416.120 ;
    END
  END ct_mem_ctrl_out[24]
  PIN ct_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 418.240 600.000 418.840 ;
    END
  END ct_mem_ctrl_out[25]
  PIN ct_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 420.960 600.000 421.560 ;
    END
  END ct_mem_ctrl_out[26]
  PIN ct_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 423.680 600.000 424.280 ;
    END
  END ct_mem_ctrl_out[27]
  PIN ct_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 426.400 600.000 427.000 ;
    END
  END ct_mem_ctrl_out[28]
  PIN ct_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 429.120 600.000 429.720 ;
    END
  END ct_mem_ctrl_out[29]
  PIN ct_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 355.000 600.000 355.600 ;
    END
  END ct_mem_ctrl_out[2]
  PIN ct_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 431.840 600.000 432.440 ;
    END
  END ct_mem_ctrl_out[30]
  PIN ct_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 434.560 600.000 435.160 ;
    END
  END ct_mem_ctrl_out[31]
  PIN ct_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 357.720 600.000 358.320 ;
    END
  END ct_mem_ctrl_out[3]
  PIN ct_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 360.440 600.000 361.040 ;
    END
  END ct_mem_ctrl_out[4]
  PIN ct_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 363.160 600.000 363.760 ;
    END
  END ct_mem_ctrl_out[5]
  PIN ct_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 365.880 600.000 366.480 ;
    END
  END ct_mem_ctrl_out[6]
  PIN ct_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 368.600 600.000 369.200 ;
    END
  END ct_mem_ctrl_out[7]
  PIN ct_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 371.320 600.000 371.920 ;
    END
  END ct_mem_ctrl_out[8]
  PIN ct_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 374.040 600.000 374.640 ;
    END
  END ct_mem_ctrl_out[9]
  PIN ct_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 437.280 600.000 437.880 ;
    END
  END ct_mem_ctrl_req
  PIN ct_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 440.000 600.000 440.600 ;
    END
  END ct_mem_ctrl_vld
  PIN ct_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 442.720 600.000 443.320 ;
    END
  END ct_mem_ctrl_we
  PIN ct_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 731.000 1.750 735.000 ;
    END
  END ct_sram0_csb0
  PIN ct_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 731.000 4.510 735.000 ;
    END
  END ct_sram0_dout0[0]
  PIN ct_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 731.000 32.570 735.000 ;
    END
  END ct_sram0_dout0[10]
  PIN ct_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 731.000 35.790 735.000 ;
    END
  END ct_sram0_dout0[11]
  PIN ct_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 731.000 38.550 735.000 ;
    END
  END ct_sram0_dout0[12]
  PIN ct_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 731.000 41.310 735.000 ;
    END
  END ct_sram0_dout0[13]
  PIN ct_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 731.000 44.070 735.000 ;
    END
  END ct_sram0_dout0[14]
  PIN ct_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 731.000 46.830 735.000 ;
    END
  END ct_sram0_dout0[15]
  PIN ct_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 731.000 50.050 735.000 ;
    END
  END ct_sram0_dout0[16]
  PIN ct_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 731.000 52.810 735.000 ;
    END
  END ct_sram0_dout0[17]
  PIN ct_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 731.000 55.570 735.000 ;
    END
  END ct_sram0_dout0[18]
  PIN ct_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 731.000 58.330 735.000 ;
    END
  END ct_sram0_dout0[19]
  PIN ct_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 731.000 7.270 735.000 ;
    END
  END ct_sram0_dout0[1]
  PIN ct_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 731.000 61.090 735.000 ;
    END
  END ct_sram0_dout0[20]
  PIN ct_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 731.000 63.850 735.000 ;
    END
  END ct_sram0_dout0[21]
  PIN ct_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 731.000 67.070 735.000 ;
    END
  END ct_sram0_dout0[22]
  PIN ct_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 731.000 69.830 735.000 ;
    END
  END ct_sram0_dout0[23]
  PIN ct_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 731.000 72.590 735.000 ;
    END
  END ct_sram0_dout0[24]
  PIN ct_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 731.000 75.350 735.000 ;
    END
  END ct_sram0_dout0[25]
  PIN ct_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 731.000 78.110 735.000 ;
    END
  END ct_sram0_dout0[26]
  PIN ct_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 731.000 81.330 735.000 ;
    END
  END ct_sram0_dout0[27]
  PIN ct_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 731.000 84.090 735.000 ;
    END
  END ct_sram0_dout0[28]
  PIN ct_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 731.000 86.850 735.000 ;
    END
  END ct_sram0_dout0[29]
  PIN ct_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 731.000 10.030 735.000 ;
    END
  END ct_sram0_dout0[2]
  PIN ct_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 731.000 89.610 735.000 ;
    END
  END ct_sram0_dout0[30]
  PIN ct_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 731.000 92.370 735.000 ;
    END
  END ct_sram0_dout0[31]
  PIN ct_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 731.000 12.790 735.000 ;
    END
  END ct_sram0_dout0[3]
  PIN ct_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 731.000 15.550 735.000 ;
    END
  END ct_sram0_dout0[4]
  PIN ct_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 731.000 18.770 735.000 ;
    END
  END ct_sram0_dout0[5]
  PIN ct_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 731.000 21.530 735.000 ;
    END
  END ct_sram0_dout0[6]
  PIN ct_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 731.000 24.290 735.000 ;
    END
  END ct_sram0_dout0[7]
  PIN ct_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 731.000 27.050 735.000 ;
    END
  END ct_sram0_dout0[8]
  PIN ct_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 731.000 29.810 735.000 ;
    END
  END ct_sram0_dout0[9]
  PIN ct_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 731.000 95.130 735.000 ;
    END
  END ct_sram0_web0
  PIN ct_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 731.000 98.350 735.000 ;
    END
  END ct_sram1_csb0
  PIN ct_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 731.000 101.110 735.000 ;
    END
  END ct_sram1_dout0[0]
  PIN ct_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 731.000 129.630 735.000 ;
    END
  END ct_sram1_dout0[10]
  PIN ct_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 731.000 132.390 735.000 ;
    END
  END ct_sram1_dout0[11]
  PIN ct_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 731.000 135.150 735.000 ;
    END
  END ct_sram1_dout0[12]
  PIN ct_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 731.000 137.910 735.000 ;
    END
  END ct_sram1_dout0[13]
  PIN ct_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 731.000 140.670 735.000 ;
    END
  END ct_sram1_dout0[14]
  PIN ct_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 731.000 143.890 735.000 ;
    END
  END ct_sram1_dout0[15]
  PIN ct_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 731.000 146.650 735.000 ;
    END
  END ct_sram1_dout0[16]
  PIN ct_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 731.000 149.410 735.000 ;
    END
  END ct_sram1_dout0[17]
  PIN ct_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 731.000 152.170 735.000 ;
    END
  END ct_sram1_dout0[18]
  PIN ct_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 731.000 154.930 735.000 ;
    END
  END ct_sram1_dout0[19]
  PIN ct_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 731.000 103.870 735.000 ;
    END
  END ct_sram1_dout0[1]
  PIN ct_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 731.000 157.690 735.000 ;
    END
  END ct_sram1_dout0[20]
  PIN ct_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 731.000 160.910 735.000 ;
    END
  END ct_sram1_dout0[21]
  PIN ct_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 731.000 163.670 735.000 ;
    END
  END ct_sram1_dout0[22]
  PIN ct_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 731.000 166.430 735.000 ;
    END
  END ct_sram1_dout0[23]
  PIN ct_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 731.000 169.190 735.000 ;
    END
  END ct_sram1_dout0[24]
  PIN ct_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 731.000 171.950 735.000 ;
    END
  END ct_sram1_dout0[25]
  PIN ct_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 731.000 174.710 735.000 ;
    END
  END ct_sram1_dout0[26]
  PIN ct_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 731.000 177.930 735.000 ;
    END
  END ct_sram1_dout0[27]
  PIN ct_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 731.000 180.690 735.000 ;
    END
  END ct_sram1_dout0[28]
  PIN ct_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 731.000 183.450 735.000 ;
    END
  END ct_sram1_dout0[29]
  PIN ct_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 731.000 106.630 735.000 ;
    END
  END ct_sram1_dout0[2]
  PIN ct_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 731.000 186.210 735.000 ;
    END
  END ct_sram1_dout0[30]
  PIN ct_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 731.000 188.970 735.000 ;
    END
  END ct_sram1_dout0[31]
  PIN ct_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 731.000 109.390 735.000 ;
    END
  END ct_sram1_dout0[3]
  PIN ct_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 731.000 112.610 735.000 ;
    END
  END ct_sram1_dout0[4]
  PIN ct_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 731.000 115.370 735.000 ;
    END
  END ct_sram1_dout0[5]
  PIN ct_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 731.000 118.130 735.000 ;
    END
  END ct_sram1_dout0[6]
  PIN ct_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 731.000 120.890 735.000 ;
    END
  END ct_sram1_dout0[7]
  PIN ct_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 731.000 123.650 735.000 ;
    END
  END ct_sram1_dout0[8]
  PIN ct_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 731.000 126.410 735.000 ;
    END
  END ct_sram1_dout0[9]
  PIN ct_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 731.000 192.190 735.000 ;
    END
  END ct_sram1_web0
  PIN ct_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 731.000 194.950 735.000 ;
    END
  END ct_sram2_csb0
  PIN ct_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 731.000 197.710 735.000 ;
    END
  END ct_sram2_dout0[0]
  PIN ct_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 731.000 226.230 735.000 ;
    END
  END ct_sram2_dout0[10]
  PIN ct_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 731.000 228.990 735.000 ;
    END
  END ct_sram2_dout0[11]
  PIN ct_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 731.000 231.750 735.000 ;
    END
  END ct_sram2_dout0[12]
  PIN ct_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 731.000 234.510 735.000 ;
    END
  END ct_sram2_dout0[13]
  PIN ct_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 731.000 237.270 735.000 ;
    END
  END ct_sram2_dout0[14]
  PIN ct_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 731.000 240.490 735.000 ;
    END
  END ct_sram2_dout0[15]
  PIN ct_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 731.000 243.250 735.000 ;
    END
  END ct_sram2_dout0[16]
  PIN ct_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 731.000 246.010 735.000 ;
    END
  END ct_sram2_dout0[17]
  PIN ct_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 731.000 248.770 735.000 ;
    END
  END ct_sram2_dout0[18]
  PIN ct_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 731.000 251.530 735.000 ;
    END
  END ct_sram2_dout0[19]
  PIN ct_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 731.000 200.470 735.000 ;
    END
  END ct_sram2_dout0[1]
  PIN ct_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 731.000 254.750 735.000 ;
    END
  END ct_sram2_dout0[20]
  PIN ct_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 731.000 257.510 735.000 ;
    END
  END ct_sram2_dout0[21]
  PIN ct_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 731.000 260.270 735.000 ;
    END
  END ct_sram2_dout0[22]
  PIN ct_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 731.000 263.030 735.000 ;
    END
  END ct_sram2_dout0[23]
  PIN ct_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 731.000 265.790 735.000 ;
    END
  END ct_sram2_dout0[24]
  PIN ct_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 731.000 268.550 735.000 ;
    END
  END ct_sram2_dout0[25]
  PIN ct_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 731.000 271.770 735.000 ;
    END
  END ct_sram2_dout0[26]
  PIN ct_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 731.000 274.530 735.000 ;
    END
  END ct_sram2_dout0[27]
  PIN ct_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 731.000 277.290 735.000 ;
    END
  END ct_sram2_dout0[28]
  PIN ct_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 731.000 280.050 735.000 ;
    END
  END ct_sram2_dout0[29]
  PIN ct_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 731.000 203.230 735.000 ;
    END
  END ct_sram2_dout0[2]
  PIN ct_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 731.000 282.810 735.000 ;
    END
  END ct_sram2_dout0[30]
  PIN ct_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 731.000 286.030 735.000 ;
    END
  END ct_sram2_dout0[31]
  PIN ct_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 731.000 205.990 735.000 ;
    END
  END ct_sram2_dout0[3]
  PIN ct_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 731.000 209.210 735.000 ;
    END
  END ct_sram2_dout0[4]
  PIN ct_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 731.000 211.970 735.000 ;
    END
  END ct_sram2_dout0[5]
  PIN ct_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 731.000 214.730 735.000 ;
    END
  END ct_sram2_dout0[6]
  PIN ct_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 731.000 217.490 735.000 ;
    END
  END ct_sram2_dout0[7]
  PIN ct_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 731.000 220.250 735.000 ;
    END
  END ct_sram2_dout0[8]
  PIN ct_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 731.000 223.470 735.000 ;
    END
  END ct_sram2_dout0[9]
  PIN ct_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 731.000 288.790 735.000 ;
    END
  END ct_sram2_web0
  PIN ct_sram3_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 731.000 291.550 735.000 ;
    END
  END ct_sram3_csb0
  PIN ct_sram3_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 731.000 294.310 735.000 ;
    END
  END ct_sram3_dout0[0]
  PIN ct_sram3_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 731.000 322.830 735.000 ;
    END
  END ct_sram3_dout0[10]
  PIN ct_sram3_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 731.000 325.590 735.000 ;
    END
  END ct_sram3_dout0[11]
  PIN ct_sram3_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 731.000 328.350 735.000 ;
    END
  END ct_sram3_dout0[12]
  PIN ct_sram3_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 731.000 331.110 735.000 ;
    END
  END ct_sram3_dout0[13]
  PIN ct_sram3_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 731.000 334.330 735.000 ;
    END
  END ct_sram3_dout0[14]
  PIN ct_sram3_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 731.000 337.090 735.000 ;
    END
  END ct_sram3_dout0[15]
  PIN ct_sram3_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 731.000 339.850 735.000 ;
    END
  END ct_sram3_dout0[16]
  PIN ct_sram3_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 731.000 342.610 735.000 ;
    END
  END ct_sram3_dout0[17]
  PIN ct_sram3_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 731.000 345.370 735.000 ;
    END
  END ct_sram3_dout0[18]
  PIN ct_sram3_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 731.000 348.130 735.000 ;
    END
  END ct_sram3_dout0[19]
  PIN ct_sram3_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 731.000 297.070 735.000 ;
    END
  END ct_sram3_dout0[1]
  PIN ct_sram3_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 731.000 351.350 735.000 ;
    END
  END ct_sram3_dout0[20]
  PIN ct_sram3_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 731.000 354.110 735.000 ;
    END
  END ct_sram3_dout0[21]
  PIN ct_sram3_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 731.000 356.870 735.000 ;
    END
  END ct_sram3_dout0[22]
  PIN ct_sram3_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 731.000 359.630 735.000 ;
    END
  END ct_sram3_dout0[23]
  PIN ct_sram3_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 731.000 362.390 735.000 ;
    END
  END ct_sram3_dout0[24]
  PIN ct_sram3_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 731.000 365.610 735.000 ;
    END
  END ct_sram3_dout0[25]
  PIN ct_sram3_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 731.000 368.370 735.000 ;
    END
  END ct_sram3_dout0[26]
  PIN ct_sram3_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 731.000 371.130 735.000 ;
    END
  END ct_sram3_dout0[27]
  PIN ct_sram3_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 731.000 373.890 735.000 ;
    END
  END ct_sram3_dout0[28]
  PIN ct_sram3_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 731.000 376.650 735.000 ;
    END
  END ct_sram3_dout0[29]
  PIN ct_sram3_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 731.000 299.830 735.000 ;
    END
  END ct_sram3_dout0[2]
  PIN ct_sram3_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 731.000 379.410 735.000 ;
    END
  END ct_sram3_dout0[30]
  PIN ct_sram3_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 731.000 382.630 735.000 ;
    END
  END ct_sram3_dout0[31]
  PIN ct_sram3_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 731.000 303.050 735.000 ;
    END
  END ct_sram3_dout0[3]
  PIN ct_sram3_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 731.000 305.810 735.000 ;
    END
  END ct_sram3_dout0[4]
  PIN ct_sram3_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 731.000 308.570 735.000 ;
    END
  END ct_sram3_dout0[5]
  PIN ct_sram3_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 731.000 311.330 735.000 ;
    END
  END ct_sram3_dout0[6]
  PIN ct_sram3_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 731.000 314.090 735.000 ;
    END
  END ct_sram3_dout0[7]
  PIN ct_sram3_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 731.000 316.850 735.000 ;
    END
  END ct_sram3_dout0[8]
  PIN ct_sram3_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 731.000 320.070 735.000 ;
    END
  END ct_sram3_dout0[9]
  PIN ct_sram3_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 731.000 385.390 735.000 ;
    END
  END ct_sram3_web0
  PIN ct_sram4_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 731.000 388.150 735.000 ;
    END
  END ct_sram4_csb0
  PIN ct_sram4_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 731.000 390.910 735.000 ;
    END
  END ct_sram4_dout0[0]
  PIN ct_sram4_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 731.000 419.430 735.000 ;
    END
  END ct_sram4_dout0[10]
  PIN ct_sram4_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 731.000 422.190 735.000 ;
    END
  END ct_sram4_dout0[11]
  PIN ct_sram4_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 731.000 424.950 735.000 ;
    END
  END ct_sram4_dout0[12]
  PIN ct_sram4_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 731.000 428.170 735.000 ;
    END
  END ct_sram4_dout0[13]
  PIN ct_sram4_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 731.000 430.930 735.000 ;
    END
  END ct_sram4_dout0[14]
  PIN ct_sram4_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 731.000 433.690 735.000 ;
    END
  END ct_sram4_dout0[15]
  PIN ct_sram4_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 731.000 436.450 735.000 ;
    END
  END ct_sram4_dout0[16]
  PIN ct_sram4_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 731.000 439.210 735.000 ;
    END
  END ct_sram4_dout0[17]
  PIN ct_sram4_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 731.000 441.970 735.000 ;
    END
  END ct_sram4_dout0[18]
  PIN ct_sram4_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 731.000 445.190 735.000 ;
    END
  END ct_sram4_dout0[19]
  PIN ct_sram4_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 731.000 393.670 735.000 ;
    END
  END ct_sram4_dout0[1]
  PIN ct_sram4_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 731.000 447.950 735.000 ;
    END
  END ct_sram4_dout0[20]
  PIN ct_sram4_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 731.000 450.710 735.000 ;
    END
  END ct_sram4_dout0[21]
  PIN ct_sram4_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 731.000 453.470 735.000 ;
    END
  END ct_sram4_dout0[22]
  PIN ct_sram4_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 731.000 456.230 735.000 ;
    END
  END ct_sram4_dout0[23]
  PIN ct_sram4_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 731.000 458.990 735.000 ;
    END
  END ct_sram4_dout0[24]
  PIN ct_sram4_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 731.000 462.210 735.000 ;
    END
  END ct_sram4_dout0[25]
  PIN ct_sram4_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 731.000 464.970 735.000 ;
    END
  END ct_sram4_dout0[26]
  PIN ct_sram4_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 731.000 467.730 735.000 ;
    END
  END ct_sram4_dout0[27]
  PIN ct_sram4_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 731.000 470.490 735.000 ;
    END
  END ct_sram4_dout0[28]
  PIN ct_sram4_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 731.000 473.250 735.000 ;
    END
  END ct_sram4_dout0[29]
  PIN ct_sram4_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 731.000 396.890 735.000 ;
    END
  END ct_sram4_dout0[2]
  PIN ct_sram4_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 731.000 476.470 735.000 ;
    END
  END ct_sram4_dout0[30]
  PIN ct_sram4_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 731.000 479.230 735.000 ;
    END
  END ct_sram4_dout0[31]
  PIN ct_sram4_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 731.000 399.650 735.000 ;
    END
  END ct_sram4_dout0[3]
  PIN ct_sram4_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 731.000 402.410 735.000 ;
    END
  END ct_sram4_dout0[4]
  PIN ct_sram4_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 731.000 405.170 735.000 ;
    END
  END ct_sram4_dout0[5]
  PIN ct_sram4_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 731.000 407.930 735.000 ;
    END
  END ct_sram4_dout0[6]
  PIN ct_sram4_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 731.000 410.690 735.000 ;
    END
  END ct_sram4_dout0[7]
  PIN ct_sram4_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 731.000 413.910 735.000 ;
    END
  END ct_sram4_dout0[8]
  PIN ct_sram4_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 731.000 416.670 735.000 ;
    END
  END ct_sram4_dout0[9]
  PIN ct_sram4_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 731.000 481.990 735.000 ;
    END
  END ct_sram4_web0
  PIN ct_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 731.000 484.750 735.000 ;
    END
  END ct_sram_comm_addr0[0]
  PIN ct_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 731.000 487.510 735.000 ;
    END
  END ct_sram_comm_addr0[1]
  PIN ct_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 731.000 490.270 735.000 ;
    END
  END ct_sram_comm_addr0[2]
  PIN ct_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 731.000 493.490 735.000 ;
    END
  END ct_sram_comm_addr0[3]
  PIN ct_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 731.000 496.250 735.000 ;
    END
  END ct_sram_comm_addr0[4]
  PIN ct_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 731.000 499.010 735.000 ;
    END
  END ct_sram_comm_addr0[5]
  PIN ct_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 731.000 501.770 735.000 ;
    END
  END ct_sram_comm_addr0[6]
  PIN ct_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 731.000 504.530 735.000 ;
    END
  END ct_sram_comm_addr0[7]
  PIN ct_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 731.000 507.750 735.000 ;
    END
  END ct_sram_comm_addr0[8]
  PIN ct_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 731.000 510.510 735.000 ;
    END
  END ct_sram_comm_din0[0]
  PIN ct_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 731.000 539.030 735.000 ;
    END
  END ct_sram_comm_din0[10]
  PIN ct_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 731.000 541.790 735.000 ;
    END
  END ct_sram_comm_din0[11]
  PIN ct_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 731.000 544.550 735.000 ;
    END
  END ct_sram_comm_din0[12]
  PIN ct_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 731.000 547.310 735.000 ;
    END
  END ct_sram_comm_din0[13]
  PIN ct_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 731.000 550.070 735.000 ;
    END
  END ct_sram_comm_din0[14]
  PIN ct_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 731.000 552.830 735.000 ;
    END
  END ct_sram_comm_din0[15]
  PIN ct_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 731.000 556.050 735.000 ;
    END
  END ct_sram_comm_din0[16]
  PIN ct_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 731.000 558.810 735.000 ;
    END
  END ct_sram_comm_din0[17]
  PIN ct_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 731.000 561.570 735.000 ;
    END
  END ct_sram_comm_din0[18]
  PIN ct_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 731.000 564.330 735.000 ;
    END
  END ct_sram_comm_din0[19]
  PIN ct_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 731.000 513.270 735.000 ;
    END
  END ct_sram_comm_din0[1]
  PIN ct_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 731.000 567.090 735.000 ;
    END
  END ct_sram_comm_din0[20]
  PIN ct_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 731.000 570.310 735.000 ;
    END
  END ct_sram_comm_din0[21]
  PIN ct_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 731.000 573.070 735.000 ;
    END
  END ct_sram_comm_din0[22]
  PIN ct_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 731.000 575.830 735.000 ;
    END
  END ct_sram_comm_din0[23]
  PIN ct_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 731.000 578.590 735.000 ;
    END
  END ct_sram_comm_din0[24]
  PIN ct_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 731.000 581.350 735.000 ;
    END
  END ct_sram_comm_din0[25]
  PIN ct_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 731.000 584.110 735.000 ;
    END
  END ct_sram_comm_din0[26]
  PIN ct_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 731.000 587.330 735.000 ;
    END
  END ct_sram_comm_din0[27]
  PIN ct_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 731.000 590.090 735.000 ;
    END
  END ct_sram_comm_din0[28]
  PIN ct_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 731.000 592.850 735.000 ;
    END
  END ct_sram_comm_din0[29]
  PIN ct_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 731.000 516.030 735.000 ;
    END
  END ct_sram_comm_din0[2]
  PIN ct_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 731.000 595.610 735.000 ;
    END
  END ct_sram_comm_din0[30]
  PIN ct_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 731.000 598.370 735.000 ;
    END
  END ct_sram_comm_din0[31]
  PIN ct_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 731.000 518.790 735.000 ;
    END
  END ct_sram_comm_din0[3]
  PIN ct_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 731.000 521.550 735.000 ;
    END
  END ct_sram_comm_din0[4]
  PIN ct_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 731.000 524.770 735.000 ;
    END
  END ct_sram_comm_din0[5]
  PIN ct_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 731.000 527.530 735.000 ;
    END
  END ct_sram_comm_din0[6]
  PIN ct_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 731.000 530.290 735.000 ;
    END
  END ct_sram_comm_din0[7]
  PIN ct_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 731.000 533.050 735.000 ;
    END
  END ct_sram_comm_din0[8]
  PIN ct_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 731.000 535.810 735.000 ;
    END
  END ct_sram_comm_din0[9]
  PIN main_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END main_mem_addr[0]
  PIN main_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END main_mem_addr[1]
  PIN main_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END main_mem_addr[2]
  PIN main_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END main_mem_addr[3]
  PIN main_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END main_mem_addr[4]
  PIN main_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END main_mem_addr[5]
  PIN main_mem_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END main_mem_in[0]
  PIN main_mem_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END main_mem_in[10]
  PIN main_mem_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END main_mem_in[11]
  PIN main_mem_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END main_mem_in[12]
  PIN main_mem_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END main_mem_in[13]
  PIN main_mem_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END main_mem_in[14]
  PIN main_mem_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END main_mem_in[15]
  PIN main_mem_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END main_mem_in[16]
  PIN main_mem_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END main_mem_in[17]
  PIN main_mem_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END main_mem_in[18]
  PIN main_mem_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END main_mem_in[19]
  PIN main_mem_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END main_mem_in[1]
  PIN main_mem_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END main_mem_in[20]
  PIN main_mem_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END main_mem_in[21]
  PIN main_mem_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END main_mem_in[22]
  PIN main_mem_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END main_mem_in[23]
  PIN main_mem_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END main_mem_in[24]
  PIN main_mem_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END main_mem_in[25]
  PIN main_mem_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END main_mem_in[26]
  PIN main_mem_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END main_mem_in[27]
  PIN main_mem_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END main_mem_in[28]
  PIN main_mem_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END main_mem_in[29]
  PIN main_mem_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END main_mem_in[2]
  PIN main_mem_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END main_mem_in[30]
  PIN main_mem_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END main_mem_in[31]
  PIN main_mem_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END main_mem_in[3]
  PIN main_mem_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END main_mem_in[4]
  PIN main_mem_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END main_mem_in[5]
  PIN main_mem_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END main_mem_in[6]
  PIN main_mem_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END main_mem_in[7]
  PIN main_mem_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END main_mem_in[8]
  PIN main_mem_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END main_mem_in[9]
  PIN main_mem_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END main_mem_out[0]
  PIN main_mem_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END main_mem_out[10]
  PIN main_mem_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END main_mem_out[11]
  PIN main_mem_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END main_mem_out[12]
  PIN main_mem_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END main_mem_out[13]
  PIN main_mem_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END main_mem_out[14]
  PIN main_mem_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END main_mem_out[15]
  PIN main_mem_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END main_mem_out[16]
  PIN main_mem_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END main_mem_out[17]
  PIN main_mem_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END main_mem_out[18]
  PIN main_mem_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END main_mem_out[19]
  PIN main_mem_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END main_mem_out[1]
  PIN main_mem_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END main_mem_out[20]
  PIN main_mem_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END main_mem_out[21]
  PIN main_mem_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END main_mem_out[22]
  PIN main_mem_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END main_mem_out[23]
  PIN main_mem_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END main_mem_out[24]
  PIN main_mem_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END main_mem_out[25]
  PIN main_mem_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END main_mem_out[26]
  PIN main_mem_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END main_mem_out[27]
  PIN main_mem_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END main_mem_out[28]
  PIN main_mem_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END main_mem_out[29]
  PIN main_mem_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END main_mem_out[2]
  PIN main_mem_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END main_mem_out[30]
  PIN main_mem_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END main_mem_out[31]
  PIN main_mem_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END main_mem_out[3]
  PIN main_mem_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END main_mem_out[4]
  PIN main_mem_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END main_mem_out[5]
  PIN main_mem_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END main_mem_out[6]
  PIN main_mem_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END main_mem_out[7]
  PIN main_mem_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END main_mem_out[8]
  PIN main_mem_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END main_mem_out[9]
  PIN main_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END main_mem_we
  PIN program_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 673.240 600.000 673.840 ;
    END
  END program_sel[0]
  PIN program_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 675.960 600.000 676.560 ;
    END
  END program_sel[1]
  PIN r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 714.040 600.000 714.640 ;
    END
  END r_data[0]
  PIN r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 716.760 600.000 717.360 ;
    END
  END r_data[1]
  PIN r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 719.480 600.000 720.080 ;
    END
  END r_data[2]
  PIN r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 722.200 600.000 722.800 ;
    END
  END r_data[3]
  PIN r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 724.920 600.000 725.520 ;
    END
  END r_data[4]
  PIN r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 727.640 600.000 728.240 ;
    END
  END r_data[5]
  PIN r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 730.360 600.000 730.960 ;
    END
  END r_data[6]
  PIN r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 733.080 600.000 733.680 ;
    END
  END r_data[7]
  PIN rd_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 681.400 600.000 682.000 ;
    END
  END rd_uart
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 667.800 600.000 668.400 ;
    END
  END rst
  PIN rst_asserted
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 670.520 600.000 671.120 ;
    END
  END rst_asserted
  PIN rx_empty
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 711.320 600.000 711.920 ;
    END
  END rx_empty
  PIN rx_fifo_flush_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 678.680 600.000 679.280 ;
    END
  END rx_fifo_flush_enable
  PIN sram_const_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END sram_const_addr1[0]
  PIN sram_const_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END sram_const_addr1[1]
  PIN sram_const_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END sram_const_addr1[2]
  PIN sram_const_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END sram_const_addr1[3]
  PIN sram_const_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END sram_const_addr1[4]
  PIN sram_const_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END sram_const_addr1[5]
  PIN sram_const_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END sram_const_addr1[6]
  PIN sram_const_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END sram_const_addr1[7]
  PIN sram_const_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END sram_const_addr1[8]
  PIN sram_const_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END sram_const_csb1
  PIN sram_const_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END sram_const_wmask0[0]
  PIN sram_const_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END sram_const_wmask0[1]
  PIN sram_const_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END sram_const_wmask0[2]
  PIN sram_const_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END sram_const_wmask0[3]
  PIN tx_full
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 708.600 600.000 709.200 ;
    END
  END tx_full
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 723.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 723.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 723.760 ;
    END
  END vssd1
  PIN w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 686.840 600.000 687.440 ;
    END
  END w_data[0]
  PIN w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 689.560 600.000 690.160 ;
    END
  END w_data[1]
  PIN w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 692.280 600.000 692.880 ;
    END
  END w_data[2]
  PIN w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 695.000 600.000 695.600 ;
    END
  END w_data[3]
  PIN w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 697.720 600.000 698.320 ;
    END
  END w_data[4]
  PIN w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 700.440 600.000 701.040 ;
    END
  END w_data[5]
  PIN w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 703.160 600.000 703.760 ;
    END
  END w_data[6]
  PIN w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 705.880 600.000 706.480 ;
    END
  END w_data[7]
  PIN wr_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 684.120 600.000 684.720 ;
    END
  END wr_uart
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 723.605 ;
      LAYER met1 ;
        RECT 1.450 5.480 599.770 725.520 ;
      LAYER met2 ;
        RECT 2.030 730.720 3.950 733.565 ;
        RECT 4.790 730.720 6.710 733.565 ;
        RECT 7.550 730.720 9.470 733.565 ;
        RECT 10.310 730.720 12.230 733.565 ;
        RECT 13.070 730.720 14.990 733.565 ;
        RECT 15.830 730.720 18.210 733.565 ;
        RECT 19.050 730.720 20.970 733.565 ;
        RECT 21.810 730.720 23.730 733.565 ;
        RECT 24.570 730.720 26.490 733.565 ;
        RECT 27.330 730.720 29.250 733.565 ;
        RECT 30.090 730.720 32.010 733.565 ;
        RECT 32.850 730.720 35.230 733.565 ;
        RECT 36.070 730.720 37.990 733.565 ;
        RECT 38.830 730.720 40.750 733.565 ;
        RECT 41.590 730.720 43.510 733.565 ;
        RECT 44.350 730.720 46.270 733.565 ;
        RECT 47.110 730.720 49.490 733.565 ;
        RECT 50.330 730.720 52.250 733.565 ;
        RECT 53.090 730.720 55.010 733.565 ;
        RECT 55.850 730.720 57.770 733.565 ;
        RECT 58.610 730.720 60.530 733.565 ;
        RECT 61.370 730.720 63.290 733.565 ;
        RECT 64.130 730.720 66.510 733.565 ;
        RECT 67.350 730.720 69.270 733.565 ;
        RECT 70.110 730.720 72.030 733.565 ;
        RECT 72.870 730.720 74.790 733.565 ;
        RECT 75.630 730.720 77.550 733.565 ;
        RECT 78.390 730.720 80.770 733.565 ;
        RECT 81.610 730.720 83.530 733.565 ;
        RECT 84.370 730.720 86.290 733.565 ;
        RECT 87.130 730.720 89.050 733.565 ;
        RECT 89.890 730.720 91.810 733.565 ;
        RECT 92.650 730.720 94.570 733.565 ;
        RECT 95.410 730.720 97.790 733.565 ;
        RECT 98.630 730.720 100.550 733.565 ;
        RECT 101.390 730.720 103.310 733.565 ;
        RECT 104.150 730.720 106.070 733.565 ;
        RECT 106.910 730.720 108.830 733.565 ;
        RECT 109.670 730.720 112.050 733.565 ;
        RECT 112.890 730.720 114.810 733.565 ;
        RECT 115.650 730.720 117.570 733.565 ;
        RECT 118.410 730.720 120.330 733.565 ;
        RECT 121.170 730.720 123.090 733.565 ;
        RECT 123.930 730.720 125.850 733.565 ;
        RECT 126.690 730.720 129.070 733.565 ;
        RECT 129.910 730.720 131.830 733.565 ;
        RECT 132.670 730.720 134.590 733.565 ;
        RECT 135.430 730.720 137.350 733.565 ;
        RECT 138.190 730.720 140.110 733.565 ;
        RECT 140.950 730.720 143.330 733.565 ;
        RECT 144.170 730.720 146.090 733.565 ;
        RECT 146.930 730.720 148.850 733.565 ;
        RECT 149.690 730.720 151.610 733.565 ;
        RECT 152.450 730.720 154.370 733.565 ;
        RECT 155.210 730.720 157.130 733.565 ;
        RECT 157.970 730.720 160.350 733.565 ;
        RECT 161.190 730.720 163.110 733.565 ;
        RECT 163.950 730.720 165.870 733.565 ;
        RECT 166.710 730.720 168.630 733.565 ;
        RECT 169.470 730.720 171.390 733.565 ;
        RECT 172.230 730.720 174.150 733.565 ;
        RECT 174.990 730.720 177.370 733.565 ;
        RECT 178.210 730.720 180.130 733.565 ;
        RECT 180.970 730.720 182.890 733.565 ;
        RECT 183.730 730.720 185.650 733.565 ;
        RECT 186.490 730.720 188.410 733.565 ;
        RECT 189.250 730.720 191.630 733.565 ;
        RECT 192.470 730.720 194.390 733.565 ;
        RECT 195.230 730.720 197.150 733.565 ;
        RECT 197.990 730.720 199.910 733.565 ;
        RECT 200.750 730.720 202.670 733.565 ;
        RECT 203.510 730.720 205.430 733.565 ;
        RECT 206.270 730.720 208.650 733.565 ;
        RECT 209.490 730.720 211.410 733.565 ;
        RECT 212.250 730.720 214.170 733.565 ;
        RECT 215.010 730.720 216.930 733.565 ;
        RECT 217.770 730.720 219.690 733.565 ;
        RECT 220.530 730.720 222.910 733.565 ;
        RECT 223.750 730.720 225.670 733.565 ;
        RECT 226.510 730.720 228.430 733.565 ;
        RECT 229.270 730.720 231.190 733.565 ;
        RECT 232.030 730.720 233.950 733.565 ;
        RECT 234.790 730.720 236.710 733.565 ;
        RECT 237.550 730.720 239.930 733.565 ;
        RECT 240.770 730.720 242.690 733.565 ;
        RECT 243.530 730.720 245.450 733.565 ;
        RECT 246.290 730.720 248.210 733.565 ;
        RECT 249.050 730.720 250.970 733.565 ;
        RECT 251.810 730.720 254.190 733.565 ;
        RECT 255.030 730.720 256.950 733.565 ;
        RECT 257.790 730.720 259.710 733.565 ;
        RECT 260.550 730.720 262.470 733.565 ;
        RECT 263.310 730.720 265.230 733.565 ;
        RECT 266.070 730.720 267.990 733.565 ;
        RECT 268.830 730.720 271.210 733.565 ;
        RECT 272.050 730.720 273.970 733.565 ;
        RECT 274.810 730.720 276.730 733.565 ;
        RECT 277.570 730.720 279.490 733.565 ;
        RECT 280.330 730.720 282.250 733.565 ;
        RECT 283.090 730.720 285.470 733.565 ;
        RECT 286.310 730.720 288.230 733.565 ;
        RECT 289.070 730.720 290.990 733.565 ;
        RECT 291.830 730.720 293.750 733.565 ;
        RECT 294.590 730.720 296.510 733.565 ;
        RECT 297.350 730.720 299.270 733.565 ;
        RECT 300.110 730.720 302.490 733.565 ;
        RECT 303.330 730.720 305.250 733.565 ;
        RECT 306.090 730.720 308.010 733.565 ;
        RECT 308.850 730.720 310.770 733.565 ;
        RECT 311.610 730.720 313.530 733.565 ;
        RECT 314.370 730.720 316.290 733.565 ;
        RECT 317.130 730.720 319.510 733.565 ;
        RECT 320.350 730.720 322.270 733.565 ;
        RECT 323.110 730.720 325.030 733.565 ;
        RECT 325.870 730.720 327.790 733.565 ;
        RECT 328.630 730.720 330.550 733.565 ;
        RECT 331.390 730.720 333.770 733.565 ;
        RECT 334.610 730.720 336.530 733.565 ;
        RECT 337.370 730.720 339.290 733.565 ;
        RECT 340.130 730.720 342.050 733.565 ;
        RECT 342.890 730.720 344.810 733.565 ;
        RECT 345.650 730.720 347.570 733.565 ;
        RECT 348.410 730.720 350.790 733.565 ;
        RECT 351.630 730.720 353.550 733.565 ;
        RECT 354.390 730.720 356.310 733.565 ;
        RECT 357.150 730.720 359.070 733.565 ;
        RECT 359.910 730.720 361.830 733.565 ;
        RECT 362.670 730.720 365.050 733.565 ;
        RECT 365.890 730.720 367.810 733.565 ;
        RECT 368.650 730.720 370.570 733.565 ;
        RECT 371.410 730.720 373.330 733.565 ;
        RECT 374.170 730.720 376.090 733.565 ;
        RECT 376.930 730.720 378.850 733.565 ;
        RECT 379.690 730.720 382.070 733.565 ;
        RECT 382.910 730.720 384.830 733.565 ;
        RECT 385.670 730.720 387.590 733.565 ;
        RECT 388.430 730.720 390.350 733.565 ;
        RECT 391.190 730.720 393.110 733.565 ;
        RECT 393.950 730.720 396.330 733.565 ;
        RECT 397.170 730.720 399.090 733.565 ;
        RECT 399.930 730.720 401.850 733.565 ;
        RECT 402.690 730.720 404.610 733.565 ;
        RECT 405.450 730.720 407.370 733.565 ;
        RECT 408.210 730.720 410.130 733.565 ;
        RECT 410.970 730.720 413.350 733.565 ;
        RECT 414.190 730.720 416.110 733.565 ;
        RECT 416.950 730.720 418.870 733.565 ;
        RECT 419.710 730.720 421.630 733.565 ;
        RECT 422.470 730.720 424.390 733.565 ;
        RECT 425.230 730.720 427.610 733.565 ;
        RECT 428.450 730.720 430.370 733.565 ;
        RECT 431.210 730.720 433.130 733.565 ;
        RECT 433.970 730.720 435.890 733.565 ;
        RECT 436.730 730.720 438.650 733.565 ;
        RECT 439.490 730.720 441.410 733.565 ;
        RECT 442.250 730.720 444.630 733.565 ;
        RECT 445.470 730.720 447.390 733.565 ;
        RECT 448.230 730.720 450.150 733.565 ;
        RECT 450.990 730.720 452.910 733.565 ;
        RECT 453.750 730.720 455.670 733.565 ;
        RECT 456.510 730.720 458.430 733.565 ;
        RECT 459.270 730.720 461.650 733.565 ;
        RECT 462.490 730.720 464.410 733.565 ;
        RECT 465.250 730.720 467.170 733.565 ;
        RECT 468.010 730.720 469.930 733.565 ;
        RECT 470.770 730.720 472.690 733.565 ;
        RECT 473.530 730.720 475.910 733.565 ;
        RECT 476.750 730.720 478.670 733.565 ;
        RECT 479.510 730.720 481.430 733.565 ;
        RECT 482.270 730.720 484.190 733.565 ;
        RECT 485.030 730.720 486.950 733.565 ;
        RECT 487.790 730.720 489.710 733.565 ;
        RECT 490.550 730.720 492.930 733.565 ;
        RECT 493.770 730.720 495.690 733.565 ;
        RECT 496.530 730.720 498.450 733.565 ;
        RECT 499.290 730.720 501.210 733.565 ;
        RECT 502.050 730.720 503.970 733.565 ;
        RECT 504.810 730.720 507.190 733.565 ;
        RECT 508.030 730.720 509.950 733.565 ;
        RECT 510.790 730.720 512.710 733.565 ;
        RECT 513.550 730.720 515.470 733.565 ;
        RECT 516.310 730.720 518.230 733.565 ;
        RECT 519.070 730.720 520.990 733.565 ;
        RECT 521.830 730.720 524.210 733.565 ;
        RECT 525.050 730.720 526.970 733.565 ;
        RECT 527.810 730.720 529.730 733.565 ;
        RECT 530.570 730.720 532.490 733.565 ;
        RECT 533.330 730.720 535.250 733.565 ;
        RECT 536.090 730.720 538.470 733.565 ;
        RECT 539.310 730.720 541.230 733.565 ;
        RECT 542.070 730.720 543.990 733.565 ;
        RECT 544.830 730.720 546.750 733.565 ;
        RECT 547.590 730.720 549.510 733.565 ;
        RECT 550.350 730.720 552.270 733.565 ;
        RECT 553.110 730.720 555.490 733.565 ;
        RECT 556.330 730.720 558.250 733.565 ;
        RECT 559.090 730.720 561.010 733.565 ;
        RECT 561.850 730.720 563.770 733.565 ;
        RECT 564.610 730.720 566.530 733.565 ;
        RECT 567.370 730.720 569.750 733.565 ;
        RECT 570.590 730.720 572.510 733.565 ;
        RECT 573.350 730.720 575.270 733.565 ;
        RECT 576.110 730.720 578.030 733.565 ;
        RECT 578.870 730.720 580.790 733.565 ;
        RECT 581.630 730.720 583.550 733.565 ;
        RECT 584.390 730.720 586.770 733.565 ;
        RECT 587.610 730.720 589.530 733.565 ;
        RECT 590.370 730.720 592.290 733.565 ;
        RECT 593.130 730.720 595.050 733.565 ;
        RECT 595.890 730.720 597.810 733.565 ;
        RECT 598.650 730.720 599.740 733.565 ;
        RECT 1.480 4.280 599.740 730.720 ;
        RECT 2.030 1.515 4.410 4.280 ;
        RECT 5.250 1.515 7.630 4.280 ;
        RECT 8.470 1.515 11.310 4.280 ;
        RECT 12.150 1.515 14.530 4.280 ;
        RECT 15.370 1.515 17.750 4.280 ;
        RECT 18.590 1.515 21.430 4.280 ;
        RECT 22.270 1.515 24.650 4.280 ;
        RECT 25.490 1.515 27.870 4.280 ;
        RECT 28.710 1.515 31.550 4.280 ;
        RECT 32.390 1.515 34.770 4.280 ;
        RECT 35.610 1.515 38.450 4.280 ;
        RECT 39.290 1.515 41.670 4.280 ;
        RECT 42.510 1.515 44.890 4.280 ;
        RECT 45.730 1.515 48.570 4.280 ;
        RECT 49.410 1.515 51.790 4.280 ;
        RECT 52.630 1.515 55.010 4.280 ;
        RECT 55.850 1.515 58.690 4.280 ;
        RECT 59.530 1.515 61.910 4.280 ;
        RECT 62.750 1.515 65.130 4.280 ;
        RECT 65.970 1.515 68.810 4.280 ;
        RECT 69.650 1.515 72.030 4.280 ;
        RECT 72.870 1.515 75.710 4.280 ;
        RECT 76.550 1.515 78.930 4.280 ;
        RECT 79.770 1.515 82.150 4.280 ;
        RECT 82.990 1.515 85.830 4.280 ;
        RECT 86.670 1.515 89.050 4.280 ;
        RECT 89.890 1.515 92.270 4.280 ;
        RECT 93.110 1.515 95.950 4.280 ;
        RECT 96.790 1.515 99.170 4.280 ;
        RECT 100.010 1.515 102.850 4.280 ;
        RECT 103.690 1.515 106.070 4.280 ;
        RECT 106.910 1.515 109.290 4.280 ;
        RECT 110.130 1.515 112.970 4.280 ;
        RECT 113.810 1.515 116.190 4.280 ;
        RECT 117.030 1.515 119.410 4.280 ;
        RECT 120.250 1.515 123.090 4.280 ;
        RECT 123.930 1.515 126.310 4.280 ;
        RECT 127.150 1.515 129.530 4.280 ;
        RECT 130.370 1.515 133.210 4.280 ;
        RECT 134.050 1.515 136.430 4.280 ;
        RECT 137.270 1.515 140.110 4.280 ;
        RECT 140.950 1.515 143.330 4.280 ;
        RECT 144.170 1.515 146.550 4.280 ;
        RECT 147.390 1.515 150.230 4.280 ;
        RECT 151.070 1.515 153.450 4.280 ;
        RECT 154.290 1.515 156.670 4.280 ;
        RECT 157.510 1.515 160.350 4.280 ;
        RECT 161.190 1.515 163.570 4.280 ;
        RECT 164.410 1.515 166.790 4.280 ;
        RECT 167.630 1.515 170.470 4.280 ;
        RECT 171.310 1.515 173.690 4.280 ;
        RECT 174.530 1.515 177.370 4.280 ;
        RECT 178.210 1.515 180.590 4.280 ;
        RECT 181.430 1.515 183.810 4.280 ;
        RECT 184.650 1.515 187.490 4.280 ;
        RECT 188.330 1.515 190.710 4.280 ;
        RECT 191.550 1.515 193.930 4.280 ;
        RECT 194.770 1.515 197.610 4.280 ;
        RECT 198.450 1.515 200.830 4.280 ;
        RECT 201.670 1.515 204.510 4.280 ;
        RECT 205.350 1.515 207.730 4.280 ;
        RECT 208.570 1.515 210.950 4.280 ;
        RECT 211.790 1.515 214.630 4.280 ;
        RECT 215.470 1.515 217.850 4.280 ;
        RECT 218.690 1.515 221.070 4.280 ;
        RECT 221.910 1.515 224.750 4.280 ;
        RECT 225.590 1.515 227.970 4.280 ;
        RECT 228.810 1.515 231.190 4.280 ;
        RECT 232.030 1.515 234.870 4.280 ;
        RECT 235.710 1.515 238.090 4.280 ;
        RECT 238.930 1.515 241.770 4.280 ;
        RECT 242.610 1.515 244.990 4.280 ;
        RECT 245.830 1.515 248.210 4.280 ;
        RECT 249.050 1.515 251.890 4.280 ;
        RECT 252.730 1.515 255.110 4.280 ;
        RECT 255.950 1.515 258.330 4.280 ;
        RECT 259.170 1.515 262.010 4.280 ;
        RECT 262.850 1.515 265.230 4.280 ;
        RECT 266.070 1.515 268.910 4.280 ;
        RECT 269.750 1.515 272.130 4.280 ;
        RECT 272.970 1.515 275.350 4.280 ;
        RECT 276.190 1.515 279.030 4.280 ;
        RECT 279.870 1.515 282.250 4.280 ;
        RECT 283.090 1.515 285.470 4.280 ;
        RECT 286.310 1.515 289.150 4.280 ;
        RECT 289.990 1.515 292.370 4.280 ;
        RECT 293.210 1.515 295.590 4.280 ;
        RECT 296.430 1.515 299.270 4.280 ;
        RECT 300.110 1.515 302.490 4.280 ;
        RECT 303.330 1.515 306.170 4.280 ;
        RECT 307.010 1.515 309.390 4.280 ;
        RECT 310.230 1.515 312.610 4.280 ;
        RECT 313.450 1.515 316.290 4.280 ;
        RECT 317.130 1.515 319.510 4.280 ;
        RECT 320.350 1.515 322.730 4.280 ;
        RECT 323.570 1.515 326.410 4.280 ;
        RECT 327.250 1.515 329.630 4.280 ;
        RECT 330.470 1.515 332.850 4.280 ;
        RECT 333.690 1.515 336.530 4.280 ;
        RECT 337.370 1.515 339.750 4.280 ;
        RECT 340.590 1.515 343.430 4.280 ;
        RECT 344.270 1.515 346.650 4.280 ;
        RECT 347.490 1.515 349.870 4.280 ;
        RECT 350.710 1.515 353.550 4.280 ;
        RECT 354.390 1.515 356.770 4.280 ;
        RECT 357.610 1.515 359.990 4.280 ;
        RECT 360.830 1.515 363.670 4.280 ;
        RECT 364.510 1.515 366.890 4.280 ;
        RECT 367.730 1.515 370.570 4.280 ;
        RECT 371.410 1.515 373.790 4.280 ;
        RECT 374.630 1.515 377.010 4.280 ;
        RECT 377.850 1.515 380.690 4.280 ;
        RECT 381.530 1.515 383.910 4.280 ;
        RECT 384.750 1.515 387.130 4.280 ;
        RECT 387.970 1.515 390.810 4.280 ;
        RECT 391.650 1.515 394.030 4.280 ;
        RECT 394.870 1.515 397.250 4.280 ;
        RECT 398.090 1.515 400.930 4.280 ;
        RECT 401.770 1.515 404.150 4.280 ;
        RECT 404.990 1.515 407.830 4.280 ;
        RECT 408.670 1.515 411.050 4.280 ;
        RECT 411.890 1.515 414.270 4.280 ;
        RECT 415.110 1.515 417.950 4.280 ;
        RECT 418.790 1.515 421.170 4.280 ;
        RECT 422.010 1.515 424.390 4.280 ;
        RECT 425.230 1.515 428.070 4.280 ;
        RECT 428.910 1.515 431.290 4.280 ;
        RECT 432.130 1.515 434.970 4.280 ;
        RECT 435.810 1.515 438.190 4.280 ;
        RECT 439.030 1.515 441.410 4.280 ;
        RECT 442.250 1.515 445.090 4.280 ;
        RECT 445.930 1.515 448.310 4.280 ;
        RECT 449.150 1.515 451.530 4.280 ;
        RECT 452.370 1.515 455.210 4.280 ;
        RECT 456.050 1.515 458.430 4.280 ;
        RECT 459.270 1.515 461.650 4.280 ;
        RECT 462.490 1.515 465.330 4.280 ;
        RECT 466.170 1.515 468.550 4.280 ;
        RECT 469.390 1.515 472.230 4.280 ;
        RECT 473.070 1.515 475.450 4.280 ;
        RECT 476.290 1.515 478.670 4.280 ;
        RECT 479.510 1.515 482.350 4.280 ;
        RECT 483.190 1.515 485.570 4.280 ;
        RECT 486.410 1.515 488.790 4.280 ;
        RECT 489.630 1.515 492.470 4.280 ;
        RECT 493.310 1.515 495.690 4.280 ;
        RECT 496.530 1.515 498.910 4.280 ;
        RECT 499.750 1.515 502.590 4.280 ;
        RECT 503.430 1.515 505.810 4.280 ;
        RECT 506.650 1.515 509.490 4.280 ;
        RECT 510.330 1.515 512.710 4.280 ;
        RECT 513.550 1.515 515.930 4.280 ;
        RECT 516.770 1.515 519.610 4.280 ;
        RECT 520.450 1.515 522.830 4.280 ;
        RECT 523.670 1.515 526.050 4.280 ;
        RECT 526.890 1.515 529.730 4.280 ;
        RECT 530.570 1.515 532.950 4.280 ;
        RECT 533.790 1.515 536.630 4.280 ;
        RECT 537.470 1.515 539.850 4.280 ;
        RECT 540.690 1.515 543.070 4.280 ;
        RECT 543.910 1.515 546.750 4.280 ;
        RECT 547.590 1.515 549.970 4.280 ;
        RECT 550.810 1.515 553.190 4.280 ;
        RECT 554.030 1.515 556.870 4.280 ;
        RECT 557.710 1.515 560.090 4.280 ;
        RECT 560.930 1.515 563.310 4.280 ;
        RECT 564.150 1.515 566.990 4.280 ;
        RECT 567.830 1.515 570.210 4.280 ;
        RECT 571.050 1.515 573.890 4.280 ;
        RECT 574.730 1.515 577.110 4.280 ;
        RECT 577.950 1.515 580.330 4.280 ;
        RECT 581.170 1.515 584.010 4.280 ;
        RECT 584.850 1.515 587.230 4.280 ;
        RECT 588.070 1.515 590.450 4.280 ;
        RECT 591.290 1.515 594.130 4.280 ;
        RECT 594.970 1.515 597.350 4.280 ;
        RECT 598.190 1.515 599.740 4.280 ;
      LAYER met3 ;
        RECT 4.400 732.680 595.600 733.545 ;
        RECT 3.990 731.360 596.555 732.680 ;
        RECT 3.990 730.680 595.600 731.360 ;
        RECT 4.400 729.960 595.600 730.680 ;
        RECT 4.400 729.280 596.555 729.960 ;
        RECT 3.990 728.640 596.555 729.280 ;
        RECT 3.990 727.280 595.600 728.640 ;
        RECT 4.400 727.240 595.600 727.280 ;
        RECT 4.400 725.920 596.555 727.240 ;
        RECT 4.400 725.880 595.600 725.920 ;
        RECT 3.990 724.560 595.600 725.880 ;
        RECT 4.400 724.520 595.600 724.560 ;
        RECT 4.400 723.200 596.555 724.520 ;
        RECT 4.400 723.160 595.600 723.200 ;
        RECT 3.990 721.800 595.600 723.160 ;
        RECT 3.990 721.160 596.555 721.800 ;
        RECT 4.400 720.480 596.555 721.160 ;
        RECT 4.400 719.760 595.600 720.480 ;
        RECT 3.990 719.080 595.600 719.760 ;
        RECT 3.990 717.760 596.555 719.080 ;
        RECT 4.400 716.360 595.600 717.760 ;
        RECT 3.990 715.040 596.555 716.360 ;
        RECT 3.990 714.360 595.600 715.040 ;
        RECT 4.400 713.640 595.600 714.360 ;
        RECT 4.400 712.960 596.555 713.640 ;
        RECT 3.990 712.320 596.555 712.960 ;
        RECT 3.990 711.640 595.600 712.320 ;
        RECT 4.400 710.920 595.600 711.640 ;
        RECT 4.400 710.240 596.555 710.920 ;
        RECT 3.990 709.600 596.555 710.240 ;
        RECT 3.990 708.240 595.600 709.600 ;
        RECT 4.400 708.200 595.600 708.240 ;
        RECT 4.400 706.880 596.555 708.200 ;
        RECT 4.400 706.840 595.600 706.880 ;
        RECT 3.990 705.480 595.600 706.840 ;
        RECT 3.990 704.840 596.555 705.480 ;
        RECT 4.400 704.160 596.555 704.840 ;
        RECT 4.400 703.440 595.600 704.160 ;
        RECT 3.990 702.760 595.600 703.440 ;
        RECT 3.990 702.120 596.555 702.760 ;
        RECT 4.400 701.440 596.555 702.120 ;
        RECT 4.400 700.720 595.600 701.440 ;
        RECT 3.990 700.040 595.600 700.720 ;
        RECT 3.990 698.720 596.555 700.040 ;
        RECT 4.400 697.320 595.600 698.720 ;
        RECT 3.990 696.000 596.555 697.320 ;
        RECT 3.990 695.320 595.600 696.000 ;
        RECT 4.400 694.600 595.600 695.320 ;
        RECT 4.400 693.920 596.555 694.600 ;
        RECT 3.990 693.280 596.555 693.920 ;
        RECT 3.990 691.920 595.600 693.280 ;
        RECT 4.400 691.880 595.600 691.920 ;
        RECT 4.400 690.560 596.555 691.880 ;
        RECT 4.400 690.520 595.600 690.560 ;
        RECT 3.990 689.200 595.600 690.520 ;
        RECT 4.400 689.160 595.600 689.200 ;
        RECT 4.400 687.840 596.555 689.160 ;
        RECT 4.400 687.800 595.600 687.840 ;
        RECT 3.990 686.440 595.600 687.800 ;
        RECT 3.990 685.800 596.555 686.440 ;
        RECT 4.400 685.120 596.555 685.800 ;
        RECT 4.400 684.400 595.600 685.120 ;
        RECT 3.990 683.720 595.600 684.400 ;
        RECT 3.990 682.400 596.555 683.720 ;
        RECT 4.400 681.000 595.600 682.400 ;
        RECT 3.990 679.680 596.555 681.000 ;
        RECT 4.400 678.280 595.600 679.680 ;
        RECT 3.990 676.960 596.555 678.280 ;
        RECT 3.990 676.280 595.600 676.960 ;
        RECT 4.400 675.560 595.600 676.280 ;
        RECT 4.400 674.880 596.555 675.560 ;
        RECT 3.990 674.240 596.555 674.880 ;
        RECT 3.990 672.880 595.600 674.240 ;
        RECT 4.400 672.840 595.600 672.880 ;
        RECT 4.400 671.520 596.555 672.840 ;
        RECT 4.400 671.480 595.600 671.520 ;
        RECT 3.990 670.120 595.600 671.480 ;
        RECT 3.990 669.480 596.555 670.120 ;
        RECT 4.400 668.800 596.555 669.480 ;
        RECT 4.400 668.080 595.600 668.800 ;
        RECT 3.990 667.400 595.600 668.080 ;
        RECT 3.990 666.760 596.555 667.400 ;
        RECT 4.400 666.080 596.555 666.760 ;
        RECT 4.400 665.360 595.600 666.080 ;
        RECT 3.990 664.680 595.600 665.360 ;
        RECT 3.990 663.360 596.555 664.680 ;
        RECT 4.400 661.960 595.600 663.360 ;
        RECT 3.990 660.640 596.555 661.960 ;
        RECT 3.990 659.960 595.600 660.640 ;
        RECT 4.400 659.240 595.600 659.960 ;
        RECT 4.400 658.560 596.555 659.240 ;
        RECT 3.990 657.920 596.555 658.560 ;
        RECT 3.990 656.560 595.600 657.920 ;
        RECT 4.400 656.520 595.600 656.560 ;
        RECT 4.400 655.160 596.555 656.520 ;
        RECT 3.990 654.520 596.555 655.160 ;
        RECT 3.990 653.840 595.600 654.520 ;
        RECT 4.400 653.120 595.600 653.840 ;
        RECT 4.400 652.440 596.555 653.120 ;
        RECT 3.990 651.800 596.555 652.440 ;
        RECT 3.990 650.440 595.600 651.800 ;
        RECT 4.400 650.400 595.600 650.440 ;
        RECT 4.400 649.080 596.555 650.400 ;
        RECT 4.400 649.040 595.600 649.080 ;
        RECT 3.990 647.680 595.600 649.040 ;
        RECT 3.990 647.040 596.555 647.680 ;
        RECT 4.400 646.360 596.555 647.040 ;
        RECT 4.400 645.640 595.600 646.360 ;
        RECT 3.990 644.960 595.600 645.640 ;
        RECT 3.990 644.320 596.555 644.960 ;
        RECT 4.400 643.640 596.555 644.320 ;
        RECT 4.400 642.920 595.600 643.640 ;
        RECT 3.990 642.240 595.600 642.920 ;
        RECT 3.990 640.920 596.555 642.240 ;
        RECT 4.400 639.520 595.600 640.920 ;
        RECT 3.990 638.200 596.555 639.520 ;
        RECT 3.990 637.520 595.600 638.200 ;
        RECT 4.400 636.800 595.600 637.520 ;
        RECT 4.400 636.120 596.555 636.800 ;
        RECT 3.990 635.480 596.555 636.120 ;
        RECT 3.990 634.120 595.600 635.480 ;
        RECT 4.400 634.080 595.600 634.120 ;
        RECT 4.400 632.760 596.555 634.080 ;
        RECT 4.400 632.720 595.600 632.760 ;
        RECT 3.990 631.400 595.600 632.720 ;
        RECT 4.400 631.360 595.600 631.400 ;
        RECT 4.400 630.040 596.555 631.360 ;
        RECT 4.400 630.000 595.600 630.040 ;
        RECT 3.990 628.640 595.600 630.000 ;
        RECT 3.990 628.000 596.555 628.640 ;
        RECT 4.400 627.320 596.555 628.000 ;
        RECT 4.400 626.600 595.600 627.320 ;
        RECT 3.990 625.920 595.600 626.600 ;
        RECT 3.990 624.600 596.555 625.920 ;
        RECT 4.400 623.200 595.600 624.600 ;
        RECT 3.990 621.880 596.555 623.200 ;
        RECT 4.400 620.480 595.600 621.880 ;
        RECT 3.990 619.160 596.555 620.480 ;
        RECT 3.990 618.480 595.600 619.160 ;
        RECT 4.400 617.760 595.600 618.480 ;
        RECT 4.400 617.080 596.555 617.760 ;
        RECT 3.990 616.440 596.555 617.080 ;
        RECT 3.990 615.080 595.600 616.440 ;
        RECT 4.400 615.040 595.600 615.080 ;
        RECT 4.400 613.720 596.555 615.040 ;
        RECT 4.400 613.680 595.600 613.720 ;
        RECT 3.990 612.320 595.600 613.680 ;
        RECT 3.990 611.680 596.555 612.320 ;
        RECT 4.400 611.000 596.555 611.680 ;
        RECT 4.400 610.280 595.600 611.000 ;
        RECT 3.990 609.600 595.600 610.280 ;
        RECT 3.990 608.960 596.555 609.600 ;
        RECT 4.400 608.280 596.555 608.960 ;
        RECT 4.400 607.560 595.600 608.280 ;
        RECT 3.990 606.880 595.600 607.560 ;
        RECT 3.990 605.560 596.555 606.880 ;
        RECT 4.400 604.160 595.600 605.560 ;
        RECT 3.990 602.840 596.555 604.160 ;
        RECT 3.990 602.160 595.600 602.840 ;
        RECT 4.400 601.440 595.600 602.160 ;
        RECT 4.400 600.760 596.555 601.440 ;
        RECT 3.990 600.120 596.555 600.760 ;
        RECT 3.990 599.440 595.600 600.120 ;
        RECT 4.400 598.720 595.600 599.440 ;
        RECT 4.400 598.040 596.555 598.720 ;
        RECT 3.990 597.400 596.555 598.040 ;
        RECT 3.990 596.040 595.600 597.400 ;
        RECT 4.400 596.000 595.600 596.040 ;
        RECT 4.400 594.680 596.555 596.000 ;
        RECT 4.400 594.640 595.600 594.680 ;
        RECT 3.990 593.280 595.600 594.640 ;
        RECT 3.990 592.640 596.555 593.280 ;
        RECT 4.400 591.960 596.555 592.640 ;
        RECT 4.400 591.240 595.600 591.960 ;
        RECT 3.990 590.560 595.600 591.240 ;
        RECT 3.990 589.240 596.555 590.560 ;
        RECT 4.400 587.840 595.600 589.240 ;
        RECT 3.990 586.520 596.555 587.840 ;
        RECT 4.400 585.120 595.600 586.520 ;
        RECT 3.990 583.800 596.555 585.120 ;
        RECT 3.990 583.120 595.600 583.800 ;
        RECT 4.400 582.400 595.600 583.120 ;
        RECT 4.400 581.720 596.555 582.400 ;
        RECT 3.990 581.080 596.555 581.720 ;
        RECT 3.990 579.720 595.600 581.080 ;
        RECT 4.400 579.680 595.600 579.720 ;
        RECT 4.400 578.360 596.555 579.680 ;
        RECT 4.400 578.320 595.600 578.360 ;
        RECT 3.990 576.960 595.600 578.320 ;
        RECT 3.990 576.320 596.555 576.960 ;
        RECT 4.400 575.640 596.555 576.320 ;
        RECT 4.400 574.920 595.600 575.640 ;
        RECT 3.990 574.240 595.600 574.920 ;
        RECT 3.990 573.600 596.555 574.240 ;
        RECT 4.400 572.240 596.555 573.600 ;
        RECT 4.400 572.200 595.600 572.240 ;
        RECT 3.990 570.840 595.600 572.200 ;
        RECT 3.990 570.200 596.555 570.840 ;
        RECT 4.400 569.520 596.555 570.200 ;
        RECT 4.400 568.800 595.600 569.520 ;
        RECT 3.990 568.120 595.600 568.800 ;
        RECT 3.990 566.800 596.555 568.120 ;
        RECT 4.400 565.400 595.600 566.800 ;
        RECT 3.990 564.080 596.555 565.400 ;
        RECT 4.400 562.680 595.600 564.080 ;
        RECT 3.990 561.360 596.555 562.680 ;
        RECT 3.990 560.680 595.600 561.360 ;
        RECT 4.400 559.960 595.600 560.680 ;
        RECT 4.400 559.280 596.555 559.960 ;
        RECT 3.990 558.640 596.555 559.280 ;
        RECT 3.990 557.280 595.600 558.640 ;
        RECT 4.400 557.240 595.600 557.280 ;
        RECT 4.400 555.920 596.555 557.240 ;
        RECT 4.400 555.880 595.600 555.920 ;
        RECT 3.990 554.520 595.600 555.880 ;
        RECT 3.990 553.880 596.555 554.520 ;
        RECT 4.400 553.200 596.555 553.880 ;
        RECT 4.400 552.480 595.600 553.200 ;
        RECT 3.990 551.800 595.600 552.480 ;
        RECT 3.990 551.160 596.555 551.800 ;
        RECT 4.400 550.480 596.555 551.160 ;
        RECT 4.400 549.760 595.600 550.480 ;
        RECT 3.990 549.080 595.600 549.760 ;
        RECT 3.990 547.760 596.555 549.080 ;
        RECT 4.400 546.360 595.600 547.760 ;
        RECT 3.990 545.040 596.555 546.360 ;
        RECT 3.990 544.360 595.600 545.040 ;
        RECT 4.400 543.640 595.600 544.360 ;
        RECT 4.400 542.960 596.555 543.640 ;
        RECT 3.990 542.320 596.555 542.960 ;
        RECT 3.990 541.640 595.600 542.320 ;
        RECT 4.400 540.920 595.600 541.640 ;
        RECT 4.400 540.240 596.555 540.920 ;
        RECT 3.990 539.600 596.555 540.240 ;
        RECT 3.990 538.240 595.600 539.600 ;
        RECT 4.400 538.200 595.600 538.240 ;
        RECT 4.400 536.880 596.555 538.200 ;
        RECT 4.400 536.840 595.600 536.880 ;
        RECT 3.990 535.480 595.600 536.840 ;
        RECT 3.990 534.840 596.555 535.480 ;
        RECT 4.400 534.160 596.555 534.840 ;
        RECT 4.400 533.440 595.600 534.160 ;
        RECT 3.990 532.760 595.600 533.440 ;
        RECT 3.990 531.440 596.555 532.760 ;
        RECT 4.400 530.040 595.600 531.440 ;
        RECT 3.990 528.720 596.555 530.040 ;
        RECT 4.400 527.320 595.600 528.720 ;
        RECT 3.990 526.000 596.555 527.320 ;
        RECT 3.990 525.320 595.600 526.000 ;
        RECT 4.400 524.600 595.600 525.320 ;
        RECT 4.400 523.920 596.555 524.600 ;
        RECT 3.990 523.280 596.555 523.920 ;
        RECT 3.990 521.920 595.600 523.280 ;
        RECT 4.400 521.880 595.600 521.920 ;
        RECT 4.400 520.560 596.555 521.880 ;
        RECT 4.400 520.520 595.600 520.560 ;
        RECT 3.990 519.200 595.600 520.520 ;
        RECT 4.400 519.160 595.600 519.200 ;
        RECT 4.400 517.840 596.555 519.160 ;
        RECT 4.400 517.800 595.600 517.840 ;
        RECT 3.990 516.440 595.600 517.800 ;
        RECT 3.990 515.800 596.555 516.440 ;
        RECT 4.400 515.120 596.555 515.800 ;
        RECT 4.400 514.400 595.600 515.120 ;
        RECT 3.990 513.720 595.600 514.400 ;
        RECT 3.990 512.400 596.555 513.720 ;
        RECT 4.400 511.000 595.600 512.400 ;
        RECT 3.990 509.680 596.555 511.000 ;
        RECT 3.990 509.000 595.600 509.680 ;
        RECT 4.400 508.280 595.600 509.000 ;
        RECT 4.400 507.600 596.555 508.280 ;
        RECT 3.990 506.960 596.555 507.600 ;
        RECT 3.990 506.280 595.600 506.960 ;
        RECT 4.400 505.560 595.600 506.280 ;
        RECT 4.400 504.880 596.555 505.560 ;
        RECT 3.990 504.240 596.555 504.880 ;
        RECT 3.990 502.880 595.600 504.240 ;
        RECT 4.400 502.840 595.600 502.880 ;
        RECT 4.400 501.520 596.555 502.840 ;
        RECT 4.400 501.480 595.600 501.520 ;
        RECT 3.990 500.120 595.600 501.480 ;
        RECT 3.990 499.480 596.555 500.120 ;
        RECT 4.400 498.800 596.555 499.480 ;
        RECT 4.400 498.080 595.600 498.800 ;
        RECT 3.990 497.400 595.600 498.080 ;
        RECT 3.990 496.080 596.555 497.400 ;
        RECT 4.400 494.680 595.600 496.080 ;
        RECT 3.990 493.360 596.555 494.680 ;
        RECT 4.400 491.960 595.600 493.360 ;
        RECT 3.990 489.960 596.555 491.960 ;
        RECT 4.400 488.560 595.600 489.960 ;
        RECT 3.990 487.240 596.555 488.560 ;
        RECT 3.990 486.560 595.600 487.240 ;
        RECT 4.400 485.840 595.600 486.560 ;
        RECT 4.400 485.160 596.555 485.840 ;
        RECT 3.990 484.520 596.555 485.160 ;
        RECT 3.990 483.840 595.600 484.520 ;
        RECT 4.400 483.120 595.600 483.840 ;
        RECT 4.400 482.440 596.555 483.120 ;
        RECT 3.990 481.800 596.555 482.440 ;
        RECT 3.990 480.440 595.600 481.800 ;
        RECT 4.400 480.400 595.600 480.440 ;
        RECT 4.400 479.080 596.555 480.400 ;
        RECT 4.400 479.040 595.600 479.080 ;
        RECT 3.990 477.680 595.600 479.040 ;
        RECT 3.990 477.040 596.555 477.680 ;
        RECT 4.400 476.360 596.555 477.040 ;
        RECT 4.400 475.640 595.600 476.360 ;
        RECT 3.990 474.960 595.600 475.640 ;
        RECT 3.990 473.640 596.555 474.960 ;
        RECT 4.400 472.240 595.600 473.640 ;
        RECT 3.990 470.920 596.555 472.240 ;
        RECT 4.400 469.520 595.600 470.920 ;
        RECT 3.990 468.200 596.555 469.520 ;
        RECT 3.990 467.520 595.600 468.200 ;
        RECT 4.400 466.800 595.600 467.520 ;
        RECT 4.400 466.120 596.555 466.800 ;
        RECT 3.990 465.480 596.555 466.120 ;
        RECT 3.990 464.120 595.600 465.480 ;
        RECT 4.400 464.080 595.600 464.120 ;
        RECT 4.400 462.760 596.555 464.080 ;
        RECT 4.400 462.720 595.600 462.760 ;
        RECT 3.990 461.400 595.600 462.720 ;
        RECT 4.400 461.360 595.600 461.400 ;
        RECT 4.400 460.040 596.555 461.360 ;
        RECT 4.400 460.000 595.600 460.040 ;
        RECT 3.990 458.640 595.600 460.000 ;
        RECT 3.990 458.000 596.555 458.640 ;
        RECT 4.400 457.320 596.555 458.000 ;
        RECT 4.400 456.600 595.600 457.320 ;
        RECT 3.990 455.920 595.600 456.600 ;
        RECT 3.990 454.600 596.555 455.920 ;
        RECT 4.400 453.200 595.600 454.600 ;
        RECT 3.990 451.880 596.555 453.200 ;
        RECT 3.990 451.200 595.600 451.880 ;
        RECT 4.400 450.480 595.600 451.200 ;
        RECT 4.400 449.800 596.555 450.480 ;
        RECT 3.990 449.160 596.555 449.800 ;
        RECT 3.990 448.480 595.600 449.160 ;
        RECT 4.400 447.760 595.600 448.480 ;
        RECT 4.400 447.080 596.555 447.760 ;
        RECT 3.990 446.440 596.555 447.080 ;
        RECT 3.990 445.080 595.600 446.440 ;
        RECT 4.400 445.040 595.600 445.080 ;
        RECT 4.400 443.720 596.555 445.040 ;
        RECT 4.400 443.680 595.600 443.720 ;
        RECT 3.990 442.320 595.600 443.680 ;
        RECT 3.990 441.680 596.555 442.320 ;
        RECT 4.400 441.000 596.555 441.680 ;
        RECT 4.400 440.280 595.600 441.000 ;
        RECT 3.990 439.600 595.600 440.280 ;
        RECT 3.990 438.280 596.555 439.600 ;
        RECT 4.400 436.880 595.600 438.280 ;
        RECT 3.990 435.560 596.555 436.880 ;
        RECT 4.400 434.160 595.600 435.560 ;
        RECT 3.990 432.840 596.555 434.160 ;
        RECT 3.990 432.160 595.600 432.840 ;
        RECT 4.400 431.440 595.600 432.160 ;
        RECT 4.400 430.760 596.555 431.440 ;
        RECT 3.990 430.120 596.555 430.760 ;
        RECT 3.990 428.760 595.600 430.120 ;
        RECT 4.400 428.720 595.600 428.760 ;
        RECT 4.400 427.400 596.555 428.720 ;
        RECT 4.400 427.360 595.600 427.400 ;
        RECT 3.990 426.040 595.600 427.360 ;
        RECT 4.400 426.000 595.600 426.040 ;
        RECT 4.400 424.680 596.555 426.000 ;
        RECT 4.400 424.640 595.600 424.680 ;
        RECT 3.990 423.280 595.600 424.640 ;
        RECT 3.990 422.640 596.555 423.280 ;
        RECT 4.400 421.960 596.555 422.640 ;
        RECT 4.400 421.240 595.600 421.960 ;
        RECT 3.990 420.560 595.600 421.240 ;
        RECT 3.990 419.240 596.555 420.560 ;
        RECT 4.400 417.840 595.600 419.240 ;
        RECT 3.990 416.520 596.555 417.840 ;
        RECT 3.990 415.840 595.600 416.520 ;
        RECT 4.400 415.120 595.600 415.840 ;
        RECT 4.400 414.440 596.555 415.120 ;
        RECT 3.990 413.800 596.555 414.440 ;
        RECT 3.990 413.120 595.600 413.800 ;
        RECT 4.400 412.400 595.600 413.120 ;
        RECT 4.400 411.720 596.555 412.400 ;
        RECT 3.990 411.080 596.555 411.720 ;
        RECT 3.990 409.720 595.600 411.080 ;
        RECT 4.400 409.680 595.600 409.720 ;
        RECT 4.400 408.320 596.555 409.680 ;
        RECT 3.990 407.680 596.555 408.320 ;
        RECT 3.990 406.320 595.600 407.680 ;
        RECT 4.400 406.280 595.600 406.320 ;
        RECT 4.400 404.960 596.555 406.280 ;
        RECT 4.400 404.920 595.600 404.960 ;
        RECT 3.990 403.600 595.600 404.920 ;
        RECT 4.400 403.560 595.600 403.600 ;
        RECT 4.400 402.240 596.555 403.560 ;
        RECT 4.400 402.200 595.600 402.240 ;
        RECT 3.990 400.840 595.600 402.200 ;
        RECT 3.990 400.200 596.555 400.840 ;
        RECT 4.400 399.520 596.555 400.200 ;
        RECT 4.400 398.800 595.600 399.520 ;
        RECT 3.990 398.120 595.600 398.800 ;
        RECT 3.990 396.800 596.555 398.120 ;
        RECT 4.400 395.400 595.600 396.800 ;
        RECT 3.990 394.080 596.555 395.400 ;
        RECT 3.990 393.400 595.600 394.080 ;
        RECT 4.400 392.680 595.600 393.400 ;
        RECT 4.400 392.000 596.555 392.680 ;
        RECT 3.990 391.360 596.555 392.000 ;
        RECT 3.990 390.680 595.600 391.360 ;
        RECT 4.400 389.960 595.600 390.680 ;
        RECT 4.400 389.280 596.555 389.960 ;
        RECT 3.990 388.640 596.555 389.280 ;
        RECT 3.990 387.280 595.600 388.640 ;
        RECT 4.400 387.240 595.600 387.280 ;
        RECT 4.400 385.920 596.555 387.240 ;
        RECT 4.400 385.880 595.600 385.920 ;
        RECT 3.990 384.520 595.600 385.880 ;
        RECT 3.990 383.880 596.555 384.520 ;
        RECT 4.400 383.200 596.555 383.880 ;
        RECT 4.400 382.480 595.600 383.200 ;
        RECT 3.990 381.800 595.600 382.480 ;
        RECT 3.990 381.160 596.555 381.800 ;
        RECT 4.400 380.480 596.555 381.160 ;
        RECT 4.400 379.760 595.600 380.480 ;
        RECT 3.990 379.080 595.600 379.760 ;
        RECT 3.990 377.760 596.555 379.080 ;
        RECT 4.400 376.360 595.600 377.760 ;
        RECT 3.990 375.040 596.555 376.360 ;
        RECT 3.990 374.360 595.600 375.040 ;
        RECT 4.400 373.640 595.600 374.360 ;
        RECT 4.400 372.960 596.555 373.640 ;
        RECT 3.990 372.320 596.555 372.960 ;
        RECT 3.990 370.960 595.600 372.320 ;
        RECT 4.400 370.920 595.600 370.960 ;
        RECT 4.400 369.600 596.555 370.920 ;
        RECT 4.400 369.560 595.600 369.600 ;
        RECT 3.990 368.240 595.600 369.560 ;
        RECT 4.400 368.200 595.600 368.240 ;
        RECT 4.400 366.880 596.555 368.200 ;
        RECT 4.400 366.840 595.600 366.880 ;
        RECT 3.990 365.480 595.600 366.840 ;
        RECT 3.990 364.840 596.555 365.480 ;
        RECT 4.400 364.160 596.555 364.840 ;
        RECT 4.400 363.440 595.600 364.160 ;
        RECT 3.990 362.760 595.600 363.440 ;
        RECT 3.990 361.440 596.555 362.760 ;
        RECT 4.400 360.040 595.600 361.440 ;
        RECT 3.990 358.720 596.555 360.040 ;
        RECT 3.990 358.040 595.600 358.720 ;
        RECT 4.400 357.320 595.600 358.040 ;
        RECT 4.400 356.640 596.555 357.320 ;
        RECT 3.990 356.000 596.555 356.640 ;
        RECT 3.990 355.320 595.600 356.000 ;
        RECT 4.400 354.600 595.600 355.320 ;
        RECT 4.400 353.920 596.555 354.600 ;
        RECT 3.990 353.280 596.555 353.920 ;
        RECT 3.990 351.920 595.600 353.280 ;
        RECT 4.400 351.880 595.600 351.920 ;
        RECT 4.400 350.560 596.555 351.880 ;
        RECT 4.400 350.520 595.600 350.560 ;
        RECT 3.990 349.160 595.600 350.520 ;
        RECT 3.990 348.520 596.555 349.160 ;
        RECT 4.400 347.840 596.555 348.520 ;
        RECT 4.400 347.120 595.600 347.840 ;
        RECT 3.990 346.440 595.600 347.120 ;
        RECT 3.990 345.800 596.555 346.440 ;
        RECT 4.400 345.120 596.555 345.800 ;
        RECT 4.400 344.400 595.600 345.120 ;
        RECT 3.990 343.720 595.600 344.400 ;
        RECT 3.990 342.400 596.555 343.720 ;
        RECT 4.400 341.000 595.600 342.400 ;
        RECT 3.990 339.680 596.555 341.000 ;
        RECT 3.990 339.000 595.600 339.680 ;
        RECT 4.400 338.280 595.600 339.000 ;
        RECT 4.400 337.600 596.555 338.280 ;
        RECT 3.990 336.960 596.555 337.600 ;
        RECT 3.990 335.600 595.600 336.960 ;
        RECT 4.400 335.560 595.600 335.600 ;
        RECT 4.400 334.240 596.555 335.560 ;
        RECT 4.400 334.200 595.600 334.240 ;
        RECT 3.990 332.880 595.600 334.200 ;
        RECT 4.400 332.840 595.600 332.880 ;
        RECT 4.400 331.520 596.555 332.840 ;
        RECT 4.400 331.480 595.600 331.520 ;
        RECT 3.990 330.120 595.600 331.480 ;
        RECT 3.990 329.480 596.555 330.120 ;
        RECT 4.400 328.120 596.555 329.480 ;
        RECT 4.400 328.080 595.600 328.120 ;
        RECT 3.990 326.720 595.600 328.080 ;
        RECT 3.990 326.080 596.555 326.720 ;
        RECT 4.400 325.400 596.555 326.080 ;
        RECT 4.400 324.680 595.600 325.400 ;
        RECT 3.990 324.000 595.600 324.680 ;
        RECT 3.990 323.360 596.555 324.000 ;
        RECT 4.400 322.680 596.555 323.360 ;
        RECT 4.400 321.960 595.600 322.680 ;
        RECT 3.990 321.280 595.600 321.960 ;
        RECT 3.990 319.960 596.555 321.280 ;
        RECT 4.400 318.560 595.600 319.960 ;
        RECT 3.990 317.240 596.555 318.560 ;
        RECT 3.990 316.560 595.600 317.240 ;
        RECT 4.400 315.840 595.600 316.560 ;
        RECT 4.400 315.160 596.555 315.840 ;
        RECT 3.990 314.520 596.555 315.160 ;
        RECT 3.990 313.160 595.600 314.520 ;
        RECT 4.400 313.120 595.600 313.160 ;
        RECT 4.400 311.800 596.555 313.120 ;
        RECT 4.400 311.760 595.600 311.800 ;
        RECT 3.990 310.440 595.600 311.760 ;
        RECT 4.400 310.400 595.600 310.440 ;
        RECT 4.400 309.080 596.555 310.400 ;
        RECT 4.400 309.040 595.600 309.080 ;
        RECT 3.990 307.680 595.600 309.040 ;
        RECT 3.990 307.040 596.555 307.680 ;
        RECT 4.400 306.360 596.555 307.040 ;
        RECT 4.400 305.640 595.600 306.360 ;
        RECT 3.990 304.960 595.600 305.640 ;
        RECT 3.990 303.640 596.555 304.960 ;
        RECT 4.400 302.240 595.600 303.640 ;
        RECT 3.990 300.920 596.555 302.240 ;
        RECT 4.400 299.520 595.600 300.920 ;
        RECT 3.990 298.200 596.555 299.520 ;
        RECT 3.990 297.520 595.600 298.200 ;
        RECT 4.400 296.800 595.600 297.520 ;
        RECT 4.400 296.120 596.555 296.800 ;
        RECT 3.990 295.480 596.555 296.120 ;
        RECT 3.990 294.120 595.600 295.480 ;
        RECT 4.400 294.080 595.600 294.120 ;
        RECT 4.400 292.760 596.555 294.080 ;
        RECT 4.400 292.720 595.600 292.760 ;
        RECT 3.990 291.360 595.600 292.720 ;
        RECT 3.990 290.720 596.555 291.360 ;
        RECT 4.400 290.040 596.555 290.720 ;
        RECT 4.400 289.320 595.600 290.040 ;
        RECT 3.990 288.640 595.600 289.320 ;
        RECT 3.990 288.000 596.555 288.640 ;
        RECT 4.400 287.320 596.555 288.000 ;
        RECT 4.400 286.600 595.600 287.320 ;
        RECT 3.990 285.920 595.600 286.600 ;
        RECT 3.990 284.600 596.555 285.920 ;
        RECT 4.400 283.200 595.600 284.600 ;
        RECT 3.990 281.880 596.555 283.200 ;
        RECT 3.990 281.200 595.600 281.880 ;
        RECT 4.400 280.480 595.600 281.200 ;
        RECT 4.400 279.800 596.555 280.480 ;
        RECT 3.990 279.160 596.555 279.800 ;
        RECT 3.990 277.800 595.600 279.160 ;
        RECT 4.400 277.760 595.600 277.800 ;
        RECT 4.400 276.440 596.555 277.760 ;
        RECT 4.400 276.400 595.600 276.440 ;
        RECT 3.990 275.080 595.600 276.400 ;
        RECT 4.400 275.040 595.600 275.080 ;
        RECT 4.400 273.720 596.555 275.040 ;
        RECT 4.400 273.680 595.600 273.720 ;
        RECT 3.990 272.320 595.600 273.680 ;
        RECT 3.990 271.680 596.555 272.320 ;
        RECT 4.400 271.000 596.555 271.680 ;
        RECT 4.400 270.280 595.600 271.000 ;
        RECT 3.990 269.600 595.600 270.280 ;
        RECT 3.990 268.280 596.555 269.600 ;
        RECT 4.400 266.880 595.600 268.280 ;
        RECT 3.990 265.560 596.555 266.880 ;
        RECT 4.400 264.160 595.600 265.560 ;
        RECT 3.990 262.840 596.555 264.160 ;
        RECT 3.990 262.160 595.600 262.840 ;
        RECT 4.400 261.440 595.600 262.160 ;
        RECT 4.400 260.760 596.555 261.440 ;
        RECT 3.990 260.120 596.555 260.760 ;
        RECT 3.990 258.760 595.600 260.120 ;
        RECT 4.400 258.720 595.600 258.760 ;
        RECT 4.400 257.400 596.555 258.720 ;
        RECT 4.400 257.360 595.600 257.400 ;
        RECT 3.990 256.000 595.600 257.360 ;
        RECT 3.990 255.360 596.555 256.000 ;
        RECT 4.400 254.680 596.555 255.360 ;
        RECT 4.400 253.960 595.600 254.680 ;
        RECT 3.990 253.280 595.600 253.960 ;
        RECT 3.990 252.640 596.555 253.280 ;
        RECT 4.400 251.960 596.555 252.640 ;
        RECT 4.400 251.240 595.600 251.960 ;
        RECT 3.990 250.560 595.600 251.240 ;
        RECT 3.990 249.240 596.555 250.560 ;
        RECT 4.400 247.840 595.600 249.240 ;
        RECT 3.990 245.840 596.555 247.840 ;
        RECT 4.400 244.440 595.600 245.840 ;
        RECT 3.990 243.120 596.555 244.440 ;
        RECT 4.400 241.720 595.600 243.120 ;
        RECT 3.990 240.400 596.555 241.720 ;
        RECT 3.990 239.720 595.600 240.400 ;
        RECT 4.400 239.000 595.600 239.720 ;
        RECT 4.400 238.320 596.555 239.000 ;
        RECT 3.990 237.680 596.555 238.320 ;
        RECT 3.990 236.320 595.600 237.680 ;
        RECT 4.400 236.280 595.600 236.320 ;
        RECT 4.400 234.960 596.555 236.280 ;
        RECT 4.400 234.920 595.600 234.960 ;
        RECT 3.990 233.560 595.600 234.920 ;
        RECT 3.990 232.920 596.555 233.560 ;
        RECT 4.400 232.240 596.555 232.920 ;
        RECT 4.400 231.520 595.600 232.240 ;
        RECT 3.990 230.840 595.600 231.520 ;
        RECT 3.990 230.200 596.555 230.840 ;
        RECT 4.400 229.520 596.555 230.200 ;
        RECT 4.400 228.800 595.600 229.520 ;
        RECT 3.990 228.120 595.600 228.800 ;
        RECT 3.990 226.800 596.555 228.120 ;
        RECT 4.400 225.400 595.600 226.800 ;
        RECT 3.990 224.080 596.555 225.400 ;
        RECT 3.990 223.400 595.600 224.080 ;
        RECT 4.400 222.680 595.600 223.400 ;
        RECT 4.400 222.000 596.555 222.680 ;
        RECT 3.990 221.360 596.555 222.000 ;
        RECT 3.990 220.000 595.600 221.360 ;
        RECT 4.400 219.960 595.600 220.000 ;
        RECT 4.400 218.640 596.555 219.960 ;
        RECT 4.400 218.600 595.600 218.640 ;
        RECT 3.990 217.280 595.600 218.600 ;
        RECT 4.400 217.240 595.600 217.280 ;
        RECT 4.400 215.920 596.555 217.240 ;
        RECT 4.400 215.880 595.600 215.920 ;
        RECT 3.990 214.520 595.600 215.880 ;
        RECT 3.990 213.880 596.555 214.520 ;
        RECT 4.400 213.200 596.555 213.880 ;
        RECT 4.400 212.480 595.600 213.200 ;
        RECT 3.990 211.800 595.600 212.480 ;
        RECT 3.990 210.480 596.555 211.800 ;
        RECT 4.400 209.080 595.600 210.480 ;
        RECT 3.990 207.760 596.555 209.080 ;
        RECT 4.400 206.360 595.600 207.760 ;
        RECT 3.990 205.040 596.555 206.360 ;
        RECT 3.990 204.360 595.600 205.040 ;
        RECT 4.400 203.640 595.600 204.360 ;
        RECT 4.400 202.960 596.555 203.640 ;
        RECT 3.990 202.320 596.555 202.960 ;
        RECT 3.990 200.960 595.600 202.320 ;
        RECT 4.400 200.920 595.600 200.960 ;
        RECT 4.400 199.600 596.555 200.920 ;
        RECT 4.400 199.560 595.600 199.600 ;
        RECT 3.990 198.200 595.600 199.560 ;
        RECT 3.990 197.560 596.555 198.200 ;
        RECT 4.400 196.880 596.555 197.560 ;
        RECT 4.400 196.160 595.600 196.880 ;
        RECT 3.990 195.480 595.600 196.160 ;
        RECT 3.990 194.840 596.555 195.480 ;
        RECT 4.400 194.160 596.555 194.840 ;
        RECT 4.400 193.440 595.600 194.160 ;
        RECT 3.990 192.760 595.600 193.440 ;
        RECT 3.990 191.440 596.555 192.760 ;
        RECT 4.400 190.040 595.600 191.440 ;
        RECT 3.990 188.720 596.555 190.040 ;
        RECT 3.990 188.040 595.600 188.720 ;
        RECT 4.400 187.320 595.600 188.040 ;
        RECT 4.400 186.640 596.555 187.320 ;
        RECT 3.990 186.000 596.555 186.640 ;
        RECT 3.990 185.320 595.600 186.000 ;
        RECT 4.400 184.600 595.600 185.320 ;
        RECT 4.400 183.920 596.555 184.600 ;
        RECT 3.990 183.280 596.555 183.920 ;
        RECT 3.990 181.920 595.600 183.280 ;
        RECT 4.400 181.880 595.600 181.920 ;
        RECT 4.400 180.560 596.555 181.880 ;
        RECT 4.400 180.520 595.600 180.560 ;
        RECT 3.990 179.160 595.600 180.520 ;
        RECT 3.990 178.520 596.555 179.160 ;
        RECT 4.400 177.840 596.555 178.520 ;
        RECT 4.400 177.120 595.600 177.840 ;
        RECT 3.990 176.440 595.600 177.120 ;
        RECT 3.990 175.120 596.555 176.440 ;
        RECT 4.400 173.720 595.600 175.120 ;
        RECT 3.990 172.400 596.555 173.720 ;
        RECT 4.400 171.000 595.600 172.400 ;
        RECT 3.990 169.680 596.555 171.000 ;
        RECT 3.990 169.000 595.600 169.680 ;
        RECT 4.400 168.280 595.600 169.000 ;
        RECT 4.400 167.600 596.555 168.280 ;
        RECT 3.990 166.960 596.555 167.600 ;
        RECT 3.990 165.600 595.600 166.960 ;
        RECT 4.400 165.560 595.600 165.600 ;
        RECT 4.400 164.200 596.555 165.560 ;
        RECT 3.990 163.560 596.555 164.200 ;
        RECT 3.990 162.880 595.600 163.560 ;
        RECT 4.400 162.160 595.600 162.880 ;
        RECT 4.400 161.480 596.555 162.160 ;
        RECT 3.990 160.840 596.555 161.480 ;
        RECT 3.990 159.480 595.600 160.840 ;
        RECT 4.400 159.440 595.600 159.480 ;
        RECT 4.400 158.120 596.555 159.440 ;
        RECT 4.400 158.080 595.600 158.120 ;
        RECT 3.990 156.720 595.600 158.080 ;
        RECT 3.990 156.080 596.555 156.720 ;
        RECT 4.400 155.400 596.555 156.080 ;
        RECT 4.400 154.680 595.600 155.400 ;
        RECT 3.990 154.000 595.600 154.680 ;
        RECT 3.990 152.680 596.555 154.000 ;
        RECT 4.400 151.280 595.600 152.680 ;
        RECT 3.990 149.960 596.555 151.280 ;
        RECT 4.400 148.560 595.600 149.960 ;
        RECT 3.990 147.240 596.555 148.560 ;
        RECT 3.990 146.560 595.600 147.240 ;
        RECT 4.400 145.840 595.600 146.560 ;
        RECT 4.400 145.160 596.555 145.840 ;
        RECT 3.990 144.520 596.555 145.160 ;
        RECT 3.990 143.160 595.600 144.520 ;
        RECT 4.400 143.120 595.600 143.160 ;
        RECT 4.400 141.800 596.555 143.120 ;
        RECT 4.400 141.760 595.600 141.800 ;
        RECT 3.990 140.400 595.600 141.760 ;
        RECT 3.990 139.760 596.555 140.400 ;
        RECT 4.400 139.080 596.555 139.760 ;
        RECT 4.400 138.360 595.600 139.080 ;
        RECT 3.990 137.680 595.600 138.360 ;
        RECT 3.990 137.040 596.555 137.680 ;
        RECT 4.400 136.360 596.555 137.040 ;
        RECT 4.400 135.640 595.600 136.360 ;
        RECT 3.990 134.960 595.600 135.640 ;
        RECT 3.990 133.640 596.555 134.960 ;
        RECT 4.400 132.240 595.600 133.640 ;
        RECT 3.990 130.920 596.555 132.240 ;
        RECT 3.990 130.240 595.600 130.920 ;
        RECT 4.400 129.520 595.600 130.240 ;
        RECT 4.400 128.840 596.555 129.520 ;
        RECT 3.990 128.200 596.555 128.840 ;
        RECT 3.990 127.520 595.600 128.200 ;
        RECT 4.400 126.800 595.600 127.520 ;
        RECT 4.400 126.120 596.555 126.800 ;
        RECT 3.990 125.480 596.555 126.120 ;
        RECT 3.990 124.120 595.600 125.480 ;
        RECT 4.400 124.080 595.600 124.120 ;
        RECT 4.400 122.760 596.555 124.080 ;
        RECT 4.400 122.720 595.600 122.760 ;
        RECT 3.990 121.360 595.600 122.720 ;
        RECT 3.990 120.720 596.555 121.360 ;
        RECT 4.400 120.040 596.555 120.720 ;
        RECT 4.400 119.320 595.600 120.040 ;
        RECT 3.990 118.640 595.600 119.320 ;
        RECT 3.990 117.320 596.555 118.640 ;
        RECT 4.400 115.920 595.600 117.320 ;
        RECT 3.990 114.600 596.555 115.920 ;
        RECT 4.400 113.200 595.600 114.600 ;
        RECT 3.990 111.880 596.555 113.200 ;
        RECT 3.990 111.200 595.600 111.880 ;
        RECT 4.400 110.480 595.600 111.200 ;
        RECT 4.400 109.800 596.555 110.480 ;
        RECT 3.990 109.160 596.555 109.800 ;
        RECT 3.990 107.800 595.600 109.160 ;
        RECT 4.400 107.760 595.600 107.800 ;
        RECT 4.400 106.440 596.555 107.760 ;
        RECT 4.400 106.400 595.600 106.440 ;
        RECT 3.990 105.080 595.600 106.400 ;
        RECT 4.400 105.040 595.600 105.080 ;
        RECT 4.400 103.720 596.555 105.040 ;
        RECT 4.400 103.680 595.600 103.720 ;
        RECT 3.990 102.320 595.600 103.680 ;
        RECT 3.990 101.680 596.555 102.320 ;
        RECT 4.400 101.000 596.555 101.680 ;
        RECT 4.400 100.280 595.600 101.000 ;
        RECT 3.990 99.600 595.600 100.280 ;
        RECT 3.990 98.280 596.555 99.600 ;
        RECT 4.400 96.880 595.600 98.280 ;
        RECT 3.990 95.560 596.555 96.880 ;
        RECT 3.990 94.880 595.600 95.560 ;
        RECT 4.400 94.160 595.600 94.880 ;
        RECT 4.400 93.480 596.555 94.160 ;
        RECT 3.990 92.840 596.555 93.480 ;
        RECT 3.990 92.160 595.600 92.840 ;
        RECT 4.400 91.440 595.600 92.160 ;
        RECT 4.400 90.760 596.555 91.440 ;
        RECT 3.990 90.120 596.555 90.760 ;
        RECT 3.990 88.760 595.600 90.120 ;
        RECT 4.400 88.720 595.600 88.760 ;
        RECT 4.400 87.400 596.555 88.720 ;
        RECT 4.400 87.360 595.600 87.400 ;
        RECT 3.990 86.000 595.600 87.360 ;
        RECT 3.990 85.360 596.555 86.000 ;
        RECT 4.400 84.680 596.555 85.360 ;
        RECT 4.400 83.960 595.600 84.680 ;
        RECT 3.990 83.280 595.600 83.960 ;
        RECT 3.990 82.640 596.555 83.280 ;
        RECT 4.400 81.280 596.555 82.640 ;
        RECT 4.400 81.240 595.600 81.280 ;
        RECT 3.990 79.880 595.600 81.240 ;
        RECT 3.990 79.240 596.555 79.880 ;
        RECT 4.400 78.560 596.555 79.240 ;
        RECT 4.400 77.840 595.600 78.560 ;
        RECT 3.990 77.160 595.600 77.840 ;
        RECT 3.990 75.840 596.555 77.160 ;
        RECT 4.400 74.440 595.600 75.840 ;
        RECT 3.990 73.120 596.555 74.440 ;
        RECT 3.990 72.440 595.600 73.120 ;
        RECT 4.400 71.720 595.600 72.440 ;
        RECT 4.400 71.040 596.555 71.720 ;
        RECT 3.990 70.400 596.555 71.040 ;
        RECT 3.990 69.720 595.600 70.400 ;
        RECT 4.400 69.000 595.600 69.720 ;
        RECT 4.400 68.320 596.555 69.000 ;
        RECT 3.990 67.680 596.555 68.320 ;
        RECT 3.990 66.320 595.600 67.680 ;
        RECT 4.400 66.280 595.600 66.320 ;
        RECT 4.400 64.960 596.555 66.280 ;
        RECT 4.400 64.920 595.600 64.960 ;
        RECT 3.990 63.560 595.600 64.920 ;
        RECT 3.990 62.920 596.555 63.560 ;
        RECT 4.400 62.240 596.555 62.920 ;
        RECT 4.400 61.520 595.600 62.240 ;
        RECT 3.990 60.840 595.600 61.520 ;
        RECT 3.990 59.520 596.555 60.840 ;
        RECT 4.400 58.120 595.600 59.520 ;
        RECT 3.990 56.800 596.555 58.120 ;
        RECT 4.400 55.400 595.600 56.800 ;
        RECT 3.990 54.080 596.555 55.400 ;
        RECT 3.990 53.400 595.600 54.080 ;
        RECT 4.400 52.680 595.600 53.400 ;
        RECT 4.400 52.000 596.555 52.680 ;
        RECT 3.990 51.360 596.555 52.000 ;
        RECT 3.990 50.000 595.600 51.360 ;
        RECT 4.400 49.960 595.600 50.000 ;
        RECT 4.400 48.640 596.555 49.960 ;
        RECT 4.400 48.600 595.600 48.640 ;
        RECT 3.990 47.280 595.600 48.600 ;
        RECT 4.400 47.240 595.600 47.280 ;
        RECT 4.400 45.920 596.555 47.240 ;
        RECT 4.400 45.880 595.600 45.920 ;
        RECT 3.990 44.520 595.600 45.880 ;
        RECT 3.990 43.880 596.555 44.520 ;
        RECT 4.400 43.200 596.555 43.880 ;
        RECT 4.400 42.480 595.600 43.200 ;
        RECT 3.990 41.800 595.600 42.480 ;
        RECT 3.990 40.480 596.555 41.800 ;
        RECT 4.400 39.080 595.600 40.480 ;
        RECT 3.990 37.760 596.555 39.080 ;
        RECT 3.990 37.080 595.600 37.760 ;
        RECT 4.400 36.360 595.600 37.080 ;
        RECT 4.400 35.680 596.555 36.360 ;
        RECT 3.990 35.040 596.555 35.680 ;
        RECT 3.990 34.360 595.600 35.040 ;
        RECT 4.400 33.640 595.600 34.360 ;
        RECT 4.400 32.960 596.555 33.640 ;
        RECT 3.990 32.320 596.555 32.960 ;
        RECT 3.990 30.960 595.600 32.320 ;
        RECT 4.400 30.920 595.600 30.960 ;
        RECT 4.400 29.600 596.555 30.920 ;
        RECT 4.400 29.560 595.600 29.600 ;
        RECT 3.990 28.200 595.600 29.560 ;
        RECT 3.990 27.560 596.555 28.200 ;
        RECT 4.400 26.880 596.555 27.560 ;
        RECT 4.400 26.160 595.600 26.880 ;
        RECT 3.990 25.480 595.600 26.160 ;
        RECT 3.990 24.840 596.555 25.480 ;
        RECT 4.400 24.160 596.555 24.840 ;
        RECT 4.400 23.440 595.600 24.160 ;
        RECT 3.990 22.760 595.600 23.440 ;
        RECT 3.990 21.440 596.555 22.760 ;
        RECT 4.400 20.040 595.600 21.440 ;
        RECT 3.990 18.720 596.555 20.040 ;
        RECT 3.990 18.040 595.600 18.720 ;
        RECT 4.400 17.320 595.600 18.040 ;
        RECT 4.400 16.640 596.555 17.320 ;
        RECT 3.990 16.000 596.555 16.640 ;
        RECT 3.990 14.640 595.600 16.000 ;
        RECT 4.400 14.600 595.600 14.640 ;
        RECT 4.400 13.280 596.555 14.600 ;
        RECT 4.400 13.240 595.600 13.280 ;
        RECT 3.990 11.920 595.600 13.240 ;
        RECT 4.400 11.880 595.600 11.920 ;
        RECT 4.400 10.560 596.555 11.880 ;
        RECT 4.400 10.520 595.600 10.560 ;
        RECT 3.990 9.160 595.600 10.520 ;
        RECT 3.990 8.520 596.555 9.160 ;
        RECT 4.400 7.840 596.555 8.520 ;
        RECT 4.400 7.120 595.600 7.840 ;
        RECT 3.990 6.440 595.600 7.120 ;
        RECT 3.990 5.120 596.555 6.440 ;
        RECT 4.400 3.720 595.600 5.120 ;
        RECT 3.990 2.400 596.555 3.720 ;
        RECT 4.400 1.535 595.600 2.400 ;
      LAYER met4 ;
        RECT 4.895 17.175 20.640 721.305 ;
        RECT 23.040 17.175 97.440 721.305 ;
        RECT 99.840 17.175 174.240 721.305 ;
        RECT 176.640 17.175 251.040 721.305 ;
        RECT 253.440 17.175 327.840 721.305 ;
        RECT 330.240 17.175 404.640 721.305 ;
        RECT 407.040 17.175 481.440 721.305 ;
        RECT 483.840 17.175 558.240 721.305 ;
        RECT 560.640 17.175 591.265 721.305 ;
  END
END main_controller
END LIBRARY

