VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO main_controller
  CLASS BLOCK ;
  FOREIGN main_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 300.000 ;
  PIN agent_1_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 296.000 1.750 300.000 ;
    END
  END agent_1_mem_ctrl_addr[0]
  PIN agent_1_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 296.000 37.170 300.000 ;
    END
  END agent_1_mem_ctrl_addr[10]
  PIN agent_1_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 296.000 40.850 300.000 ;
    END
  END agent_1_mem_ctrl_addr[11]
  PIN agent_1_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 296.000 44.530 300.000 ;
    END
  END agent_1_mem_ctrl_addr[12]
  PIN agent_1_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 296.000 48.210 300.000 ;
    END
  END agent_1_mem_ctrl_addr[13]
  PIN agent_1_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 296.000 4.970 300.000 ;
    END
  END agent_1_mem_ctrl_addr[1]
  PIN agent_1_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 296.000 8.650 300.000 ;
    END
  END agent_1_mem_ctrl_addr[2]
  PIN agent_1_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 296.000 12.330 300.000 ;
    END
  END agent_1_mem_ctrl_addr[3]
  PIN agent_1_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 296.000 16.010 300.000 ;
    END
  END agent_1_mem_ctrl_addr[4]
  PIN agent_1_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 296.000 19.230 300.000 ;
    END
  END agent_1_mem_ctrl_addr[5]
  PIN agent_1_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 296.000 22.910 300.000 ;
    END
  END agent_1_mem_ctrl_addr[6]
  PIN agent_1_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 296.000 26.590 300.000 ;
    END
  END agent_1_mem_ctrl_addr[7]
  PIN agent_1_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 296.000 30.270 300.000 ;
    END
  END agent_1_mem_ctrl_addr[8]
  PIN agent_1_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 296.000 33.950 300.000 ;
    END
  END agent_1_mem_ctrl_addr[9]
  PIN agent_1_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 296.000 51.890 300.000 ;
    END
  END agent_1_mem_ctrl_in[0]
  PIN agent_1_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 296.000 87.310 300.000 ;
    END
  END agent_1_mem_ctrl_in[10]
  PIN agent_1_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 296.000 90.990 300.000 ;
    END
  END agent_1_mem_ctrl_in[11]
  PIN agent_1_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 296.000 94.670 300.000 ;
    END
  END agent_1_mem_ctrl_in[12]
  PIN agent_1_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 296.000 98.350 300.000 ;
    END
  END agent_1_mem_ctrl_in[13]
  PIN agent_1_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 296.000 102.030 300.000 ;
    END
  END agent_1_mem_ctrl_in[14]
  PIN agent_1_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 296.000 105.250 300.000 ;
    END
  END agent_1_mem_ctrl_in[15]
  PIN agent_1_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 296.000 108.930 300.000 ;
    END
  END agent_1_mem_ctrl_in[16]
  PIN agent_1_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 296.000 112.610 300.000 ;
    END
  END agent_1_mem_ctrl_in[17]
  PIN agent_1_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 296.000 116.290 300.000 ;
    END
  END agent_1_mem_ctrl_in[18]
  PIN agent_1_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 296.000 119.970 300.000 ;
    END
  END agent_1_mem_ctrl_in[19]
  PIN agent_1_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 296.000 55.110 300.000 ;
    END
  END agent_1_mem_ctrl_in[1]
  PIN agent_1_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 296.000 123.190 300.000 ;
    END
  END agent_1_mem_ctrl_in[20]
  PIN agent_1_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 296.000 126.870 300.000 ;
    END
  END agent_1_mem_ctrl_in[21]
  PIN agent_1_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 296.000 130.550 300.000 ;
    END
  END agent_1_mem_ctrl_in[22]
  PIN agent_1_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 296.000 134.230 300.000 ;
    END
  END agent_1_mem_ctrl_in[23]
  PIN agent_1_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 296.000 137.450 300.000 ;
    END
  END agent_1_mem_ctrl_in[24]
  PIN agent_1_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 296.000 141.130 300.000 ;
    END
  END agent_1_mem_ctrl_in[25]
  PIN agent_1_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 296.000 144.810 300.000 ;
    END
  END agent_1_mem_ctrl_in[26]
  PIN agent_1_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 296.000 148.490 300.000 ;
    END
  END agent_1_mem_ctrl_in[27]
  PIN agent_1_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 296.000 152.170 300.000 ;
    END
  END agent_1_mem_ctrl_in[28]
  PIN agent_1_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 296.000 155.390 300.000 ;
    END
  END agent_1_mem_ctrl_in[29]
  PIN agent_1_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 296.000 58.790 300.000 ;
    END
  END agent_1_mem_ctrl_in[2]
  PIN agent_1_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 296.000 159.070 300.000 ;
    END
  END agent_1_mem_ctrl_in[30]
  PIN agent_1_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 296.000 162.750 300.000 ;
    END
  END agent_1_mem_ctrl_in[31]
  PIN agent_1_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 296.000 62.470 300.000 ;
    END
  END agent_1_mem_ctrl_in[3]
  PIN agent_1_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 296.000 66.150 300.000 ;
    END
  END agent_1_mem_ctrl_in[4]
  PIN agent_1_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 296.000 69.370 300.000 ;
    END
  END agent_1_mem_ctrl_in[5]
  PIN agent_1_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 296.000 73.050 300.000 ;
    END
  END agent_1_mem_ctrl_in[6]
  PIN agent_1_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 296.000 76.730 300.000 ;
    END
  END agent_1_mem_ctrl_in[7]
  PIN agent_1_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 296.000 80.410 300.000 ;
    END
  END agent_1_mem_ctrl_in[8]
  PIN agent_1_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 296.000 84.090 300.000 ;
    END
  END agent_1_mem_ctrl_in[9]
  PIN agent_1_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 296.000 166.430 300.000 ;
    END
  END agent_1_mem_ctrl_out[0]
  PIN agent_1_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 296.000 202.310 300.000 ;
    END
  END agent_1_mem_ctrl_out[10]
  PIN agent_1_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 296.000 205.530 300.000 ;
    END
  END agent_1_mem_ctrl_out[11]
  PIN agent_1_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 296.000 209.210 300.000 ;
    END
  END agent_1_mem_ctrl_out[12]
  PIN agent_1_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 296.000 212.890 300.000 ;
    END
  END agent_1_mem_ctrl_out[13]
  PIN agent_1_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 296.000 216.570 300.000 ;
    END
  END agent_1_mem_ctrl_out[14]
  PIN agent_1_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 296.000 220.250 300.000 ;
    END
  END agent_1_mem_ctrl_out[15]
  PIN agent_1_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 296.000 223.470 300.000 ;
    END
  END agent_1_mem_ctrl_out[16]
  PIN agent_1_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 296.000 227.150 300.000 ;
    END
  END agent_1_mem_ctrl_out[17]
  PIN agent_1_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 296.000 230.830 300.000 ;
    END
  END agent_1_mem_ctrl_out[18]
  PIN agent_1_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 296.000 234.510 300.000 ;
    END
  END agent_1_mem_ctrl_out[19]
  PIN agent_1_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 296.000 170.110 300.000 ;
    END
  END agent_1_mem_ctrl_out[1]
  PIN agent_1_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 296.000 238.190 300.000 ;
    END
  END agent_1_mem_ctrl_out[20]
  PIN agent_1_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 296.000 241.410 300.000 ;
    END
  END agent_1_mem_ctrl_out[21]
  PIN agent_1_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 296.000 245.090 300.000 ;
    END
  END agent_1_mem_ctrl_out[22]
  PIN agent_1_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 296.000 248.770 300.000 ;
    END
  END agent_1_mem_ctrl_out[23]
  PIN agent_1_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 296.000 252.450 300.000 ;
    END
  END agent_1_mem_ctrl_out[24]
  PIN agent_1_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 296.000 255.670 300.000 ;
    END
  END agent_1_mem_ctrl_out[25]
  PIN agent_1_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 296.000 259.350 300.000 ;
    END
  END agent_1_mem_ctrl_out[26]
  PIN agent_1_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 296.000 263.030 300.000 ;
    END
  END agent_1_mem_ctrl_out[27]
  PIN agent_1_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 296.000 266.710 300.000 ;
    END
  END agent_1_mem_ctrl_out[28]
  PIN agent_1_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 296.000 270.390 300.000 ;
    END
  END agent_1_mem_ctrl_out[29]
  PIN agent_1_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 296.000 173.330 300.000 ;
    END
  END agent_1_mem_ctrl_out[2]
  PIN agent_1_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 296.000 273.610 300.000 ;
    END
  END agent_1_mem_ctrl_out[30]
  PIN agent_1_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 296.000 277.290 300.000 ;
    END
  END agent_1_mem_ctrl_out[31]
  PIN agent_1_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 296.000 177.010 300.000 ;
    END
  END agent_1_mem_ctrl_out[3]
  PIN agent_1_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 296.000 180.690 300.000 ;
    END
  END agent_1_mem_ctrl_out[4]
  PIN agent_1_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 296.000 184.370 300.000 ;
    END
  END agent_1_mem_ctrl_out[5]
  PIN agent_1_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 296.000 187.590 300.000 ;
    END
  END agent_1_mem_ctrl_out[6]
  PIN agent_1_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 296.000 191.270 300.000 ;
    END
  END agent_1_mem_ctrl_out[7]
  PIN agent_1_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 296.000 194.950 300.000 ;
    END
  END agent_1_mem_ctrl_out[8]
  PIN agent_1_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 296.000 198.630 300.000 ;
    END
  END agent_1_mem_ctrl_out[9]
  PIN agent_1_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 296.000 280.970 300.000 ;
    END
  END agent_1_mem_ctrl_req
  PIN agent_1_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 296.000 284.650 300.000 ;
    END
  END agent_1_mem_ctrl_vld
  PIN agent_1_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 296.000 288.330 300.000 ;
    END
  END agent_1_mem_ctrl_we
  PIN agent_1_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END agent_1_sram0_csb0
  PIN agent_1_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END agent_1_sram0_dout0[0]
  PIN agent_1_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END agent_1_sram0_dout0[10]
  PIN agent_1_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END agent_1_sram0_dout0[11]
  PIN agent_1_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END agent_1_sram0_dout0[12]
  PIN agent_1_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END agent_1_sram0_dout0[13]
  PIN agent_1_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END agent_1_sram0_dout0[14]
  PIN agent_1_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END agent_1_sram0_dout0[15]
  PIN agent_1_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END agent_1_sram0_dout0[16]
  PIN agent_1_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END agent_1_sram0_dout0[17]
  PIN agent_1_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END agent_1_sram0_dout0[18]
  PIN agent_1_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END agent_1_sram0_dout0[19]
  PIN agent_1_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END agent_1_sram0_dout0[1]
  PIN agent_1_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END agent_1_sram0_dout0[20]
  PIN agent_1_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END agent_1_sram0_dout0[21]
  PIN agent_1_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END agent_1_sram0_dout0[22]
  PIN agent_1_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END agent_1_sram0_dout0[23]
  PIN agent_1_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END agent_1_sram0_dout0[24]
  PIN agent_1_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END agent_1_sram0_dout0[25]
  PIN agent_1_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END agent_1_sram0_dout0[26]
  PIN agent_1_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END agent_1_sram0_dout0[27]
  PIN agent_1_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END agent_1_sram0_dout0[28]
  PIN agent_1_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END agent_1_sram0_dout0[29]
  PIN agent_1_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END agent_1_sram0_dout0[2]
  PIN agent_1_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END agent_1_sram0_dout0[30]
  PIN agent_1_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END agent_1_sram0_dout0[31]
  PIN agent_1_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END agent_1_sram0_dout0[3]
  PIN agent_1_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END agent_1_sram0_dout0[4]
  PIN agent_1_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END agent_1_sram0_dout0[5]
  PIN agent_1_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END agent_1_sram0_dout0[6]
  PIN agent_1_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END agent_1_sram0_dout0[7]
  PIN agent_1_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END agent_1_sram0_dout0[8]
  PIN agent_1_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END agent_1_sram0_dout0[9]
  PIN agent_1_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END agent_1_sram0_web0
  PIN agent_1_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END agent_1_sram1_csb0
  PIN agent_1_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END agent_1_sram1_dout0[0]
  PIN agent_1_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END agent_1_sram1_dout0[10]
  PIN agent_1_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END agent_1_sram1_dout0[11]
  PIN agent_1_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END agent_1_sram1_dout0[12]
  PIN agent_1_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END agent_1_sram1_dout0[13]
  PIN agent_1_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END agent_1_sram1_dout0[14]
  PIN agent_1_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END agent_1_sram1_dout0[15]
  PIN agent_1_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END agent_1_sram1_dout0[16]
  PIN agent_1_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END agent_1_sram1_dout0[17]
  PIN agent_1_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END agent_1_sram1_dout0[18]
  PIN agent_1_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END agent_1_sram1_dout0[19]
  PIN agent_1_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END agent_1_sram1_dout0[1]
  PIN agent_1_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END agent_1_sram1_dout0[20]
  PIN agent_1_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END agent_1_sram1_dout0[21]
  PIN agent_1_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END agent_1_sram1_dout0[22]
  PIN agent_1_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END agent_1_sram1_dout0[23]
  PIN agent_1_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END agent_1_sram1_dout0[24]
  PIN agent_1_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END agent_1_sram1_dout0[25]
  PIN agent_1_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END agent_1_sram1_dout0[26]
  PIN agent_1_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END agent_1_sram1_dout0[27]
  PIN agent_1_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END agent_1_sram1_dout0[28]
  PIN agent_1_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END agent_1_sram1_dout0[29]
  PIN agent_1_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END agent_1_sram1_dout0[2]
  PIN agent_1_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END agent_1_sram1_dout0[30]
  PIN agent_1_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END agent_1_sram1_dout0[31]
  PIN agent_1_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END agent_1_sram1_dout0[3]
  PIN agent_1_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END agent_1_sram1_dout0[4]
  PIN agent_1_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END agent_1_sram1_dout0[5]
  PIN agent_1_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END agent_1_sram1_dout0[6]
  PIN agent_1_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END agent_1_sram1_dout0[7]
  PIN agent_1_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END agent_1_sram1_dout0[8]
  PIN agent_1_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END agent_1_sram1_dout0[9]
  PIN agent_1_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END agent_1_sram1_web0
  PIN agent_1_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END agent_1_sram2_csb0
  PIN agent_1_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END agent_1_sram2_dout0[0]
  PIN agent_1_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END agent_1_sram2_dout0[10]
  PIN agent_1_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END agent_1_sram2_dout0[11]
  PIN agent_1_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END agent_1_sram2_dout0[12]
  PIN agent_1_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END agent_1_sram2_dout0[13]
  PIN agent_1_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END agent_1_sram2_dout0[14]
  PIN agent_1_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END agent_1_sram2_dout0[15]
  PIN agent_1_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END agent_1_sram2_dout0[16]
  PIN agent_1_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END agent_1_sram2_dout0[17]
  PIN agent_1_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END agent_1_sram2_dout0[18]
  PIN agent_1_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END agent_1_sram2_dout0[19]
  PIN agent_1_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END agent_1_sram2_dout0[1]
  PIN agent_1_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END agent_1_sram2_dout0[20]
  PIN agent_1_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END agent_1_sram2_dout0[21]
  PIN agent_1_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END agent_1_sram2_dout0[22]
  PIN agent_1_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END agent_1_sram2_dout0[23]
  PIN agent_1_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END agent_1_sram2_dout0[24]
  PIN agent_1_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END agent_1_sram2_dout0[25]
  PIN agent_1_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END agent_1_sram2_dout0[26]
  PIN agent_1_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END agent_1_sram2_dout0[27]
  PIN agent_1_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END agent_1_sram2_dout0[28]
  PIN agent_1_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END agent_1_sram2_dout0[29]
  PIN agent_1_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END agent_1_sram2_dout0[2]
  PIN agent_1_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END agent_1_sram2_dout0[30]
  PIN agent_1_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END agent_1_sram2_dout0[31]
  PIN agent_1_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END agent_1_sram2_dout0[3]
  PIN agent_1_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END agent_1_sram2_dout0[4]
  PIN agent_1_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END agent_1_sram2_dout0[5]
  PIN agent_1_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END agent_1_sram2_dout0[6]
  PIN agent_1_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END agent_1_sram2_dout0[7]
  PIN agent_1_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END agent_1_sram2_dout0[8]
  PIN agent_1_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END agent_1_sram2_dout0[9]
  PIN agent_1_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END agent_1_sram2_web0
  PIN agent_1_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END agent_1_sram_comm_addr0[0]
  PIN agent_1_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END agent_1_sram_comm_addr0[1]
  PIN agent_1_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END agent_1_sram_comm_addr0[2]
  PIN agent_1_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END agent_1_sram_comm_addr0[3]
  PIN agent_1_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END agent_1_sram_comm_addr0[4]
  PIN agent_1_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END agent_1_sram_comm_addr0[5]
  PIN agent_1_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END agent_1_sram_comm_addr0[6]
  PIN agent_1_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END agent_1_sram_comm_addr0[7]
  PIN agent_1_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END agent_1_sram_comm_addr0[8]
  PIN agent_1_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END agent_1_sram_comm_din0[0]
  PIN agent_1_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END agent_1_sram_comm_din0[10]
  PIN agent_1_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END agent_1_sram_comm_din0[11]
  PIN agent_1_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END agent_1_sram_comm_din0[12]
  PIN agent_1_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END agent_1_sram_comm_din0[13]
  PIN agent_1_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END agent_1_sram_comm_din0[14]
  PIN agent_1_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END agent_1_sram_comm_din0[15]
  PIN agent_1_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END agent_1_sram_comm_din0[16]
  PIN agent_1_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END agent_1_sram_comm_din0[17]
  PIN agent_1_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END agent_1_sram_comm_din0[18]
  PIN agent_1_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END agent_1_sram_comm_din0[19]
  PIN agent_1_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END agent_1_sram_comm_din0[1]
  PIN agent_1_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END agent_1_sram_comm_din0[20]
  PIN agent_1_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END agent_1_sram_comm_din0[21]
  PIN agent_1_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END agent_1_sram_comm_din0[22]
  PIN agent_1_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END agent_1_sram_comm_din0[23]
  PIN agent_1_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END agent_1_sram_comm_din0[24]
  PIN agent_1_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END agent_1_sram_comm_din0[25]
  PIN agent_1_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END agent_1_sram_comm_din0[26]
  PIN agent_1_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END agent_1_sram_comm_din0[27]
  PIN agent_1_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END agent_1_sram_comm_din0[28]
  PIN agent_1_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END agent_1_sram_comm_din0[29]
  PIN agent_1_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END agent_1_sram_comm_din0[2]
  PIN agent_1_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END agent_1_sram_comm_din0[30]
  PIN agent_1_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END agent_1_sram_comm_din0[31]
  PIN agent_1_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END agent_1_sram_comm_din0[3]
  PIN agent_1_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END agent_1_sram_comm_din0[4]
  PIN agent_1_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END agent_1_sram_comm_din0[5]
  PIN agent_1_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END agent_1_sram_comm_din0[6]
  PIN agent_1_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END agent_1_sram_comm_din0[7]
  PIN agent_1_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END agent_1_sram_comm_din0[8]
  PIN agent_1_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END agent_1_sram_comm_din0[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END clk
  PIN cm_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 296.000 581.810 300.000 ;
    END
  END cm_mem_ctrl_addr[0]
  PIN cm_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 296.000 617.690 300.000 ;
    END
  END cm_mem_ctrl_addr[10]
  PIN cm_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 296.000 621.370 300.000 ;
    END
  END cm_mem_ctrl_addr[11]
  PIN cm_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 296.000 625.050 300.000 ;
    END
  END cm_mem_ctrl_addr[12]
  PIN cm_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 296.000 628.270 300.000 ;
    END
  END cm_mem_ctrl_addr[13]
  PIN cm_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 296.000 585.490 300.000 ;
    END
  END cm_mem_ctrl_addr[1]
  PIN cm_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 296.000 589.170 300.000 ;
    END
  END cm_mem_ctrl_addr[2]
  PIN cm_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 296.000 592.850 300.000 ;
    END
  END cm_mem_ctrl_addr[3]
  PIN cm_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 296.000 596.070 300.000 ;
    END
  END cm_mem_ctrl_addr[4]
  PIN cm_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 296.000 599.750 300.000 ;
    END
  END cm_mem_ctrl_addr[5]
  PIN cm_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 296.000 603.430 300.000 ;
    END
  END cm_mem_ctrl_addr[6]
  PIN cm_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 296.000 607.110 300.000 ;
    END
  END cm_mem_ctrl_addr[7]
  PIN cm_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 296.000 610.330 300.000 ;
    END
  END cm_mem_ctrl_addr[8]
  PIN cm_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 296.000 614.010 300.000 ;
    END
  END cm_mem_ctrl_addr[9]
  PIN cm_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 296.000 631.950 300.000 ;
    END
  END cm_mem_ctrl_in[0]
  PIN cm_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 296.000 667.830 300.000 ;
    END
  END cm_mem_ctrl_in[10]
  PIN cm_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 296.000 671.510 300.000 ;
    END
  END cm_mem_ctrl_in[11]
  PIN cm_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 296.000 675.190 300.000 ;
    END
  END cm_mem_ctrl_in[12]
  PIN cm_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 296.000 678.410 300.000 ;
    END
  END cm_mem_ctrl_in[13]
  PIN cm_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 296.000 682.090 300.000 ;
    END
  END cm_mem_ctrl_in[14]
  PIN cm_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 296.000 685.770 300.000 ;
    END
  END cm_mem_ctrl_in[15]
  PIN cm_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 296.000 689.450 300.000 ;
    END
  END cm_mem_ctrl_in[16]
  PIN cm_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 296.000 693.130 300.000 ;
    END
  END cm_mem_ctrl_in[17]
  PIN cm_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 296.000 696.350 300.000 ;
    END
  END cm_mem_ctrl_in[18]
  PIN cm_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 296.000 700.030 300.000 ;
    END
  END cm_mem_ctrl_in[19]
  PIN cm_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 296.000 635.630 300.000 ;
    END
  END cm_mem_ctrl_in[1]
  PIN cm_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 296.000 703.710 300.000 ;
    END
  END cm_mem_ctrl_in[20]
  PIN cm_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 296.000 707.390 300.000 ;
    END
  END cm_mem_ctrl_in[21]
  PIN cm_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 296.000 711.070 300.000 ;
    END
  END cm_mem_ctrl_in[22]
  PIN cm_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 296.000 714.290 300.000 ;
    END
  END cm_mem_ctrl_in[23]
  PIN cm_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 296.000 717.970 300.000 ;
    END
  END cm_mem_ctrl_in[24]
  PIN cm_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 296.000 721.650 300.000 ;
    END
  END cm_mem_ctrl_in[25]
  PIN cm_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 296.000 725.330 300.000 ;
    END
  END cm_mem_ctrl_in[26]
  PIN cm_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 296.000 728.550 300.000 ;
    END
  END cm_mem_ctrl_in[27]
  PIN cm_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 296.000 732.230 300.000 ;
    END
  END cm_mem_ctrl_in[28]
  PIN cm_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 296.000 735.910 300.000 ;
    END
  END cm_mem_ctrl_in[29]
  PIN cm_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 296.000 639.310 300.000 ;
    END
  END cm_mem_ctrl_in[2]
  PIN cm_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 296.000 739.590 300.000 ;
    END
  END cm_mem_ctrl_in[30]
  PIN cm_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 296.000 743.270 300.000 ;
    END
  END cm_mem_ctrl_in[31]
  PIN cm_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 296.000 642.990 300.000 ;
    END
  END cm_mem_ctrl_in[3]
  PIN cm_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 296.000 646.210 300.000 ;
    END
  END cm_mem_ctrl_in[4]
  PIN cm_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 296.000 649.890 300.000 ;
    END
  END cm_mem_ctrl_in[5]
  PIN cm_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 296.000 653.570 300.000 ;
    END
  END cm_mem_ctrl_in[6]
  PIN cm_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 296.000 657.250 300.000 ;
    END
  END cm_mem_ctrl_in[7]
  PIN cm_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 296.000 660.930 300.000 ;
    END
  END cm_mem_ctrl_in[8]
  PIN cm_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 296.000 664.150 300.000 ;
    END
  END cm_mem_ctrl_in[9]
  PIN cm_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 296.000 746.490 300.000 ;
    END
  END cm_mem_ctrl_out[0]
  PIN cm_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 296.000 782.370 300.000 ;
    END
  END cm_mem_ctrl_out[10]
  PIN cm_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 296.000 786.050 300.000 ;
    END
  END cm_mem_ctrl_out[11]
  PIN cm_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 296.000 789.730 300.000 ;
    END
  END cm_mem_ctrl_out[12]
  PIN cm_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 296.000 793.410 300.000 ;
    END
  END cm_mem_ctrl_out[13]
  PIN cm_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 296.000 796.630 300.000 ;
    END
  END cm_mem_ctrl_out[14]
  PIN cm_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 296.000 800.310 300.000 ;
    END
  END cm_mem_ctrl_out[15]
  PIN cm_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 296.000 803.990 300.000 ;
    END
  END cm_mem_ctrl_out[16]
  PIN cm_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 296.000 807.670 300.000 ;
    END
  END cm_mem_ctrl_out[17]
  PIN cm_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 296.000 811.350 300.000 ;
    END
  END cm_mem_ctrl_out[18]
  PIN cm_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 296.000 814.570 300.000 ;
    END
  END cm_mem_ctrl_out[19]
  PIN cm_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 296.000 750.170 300.000 ;
    END
  END cm_mem_ctrl_out[1]
  PIN cm_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 296.000 818.250 300.000 ;
    END
  END cm_mem_ctrl_out[20]
  PIN cm_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 296.000 821.930 300.000 ;
    END
  END cm_mem_ctrl_out[21]
  PIN cm_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 296.000 825.610 300.000 ;
    END
  END cm_mem_ctrl_out[22]
  PIN cm_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 296.000 829.290 300.000 ;
    END
  END cm_mem_ctrl_out[23]
  PIN cm_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 296.000 832.510 300.000 ;
    END
  END cm_mem_ctrl_out[24]
  PIN cm_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 296.000 836.190 300.000 ;
    END
  END cm_mem_ctrl_out[25]
  PIN cm_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 296.000 839.870 300.000 ;
    END
  END cm_mem_ctrl_out[26]
  PIN cm_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 296.000 843.550 300.000 ;
    END
  END cm_mem_ctrl_out[27]
  PIN cm_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 296.000 846.770 300.000 ;
    END
  END cm_mem_ctrl_out[28]
  PIN cm_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 296.000 850.450 300.000 ;
    END
  END cm_mem_ctrl_out[29]
  PIN cm_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 296.000 753.850 300.000 ;
    END
  END cm_mem_ctrl_out[2]
  PIN cm_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 296.000 854.130 300.000 ;
    END
  END cm_mem_ctrl_out[30]
  PIN cm_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.530 296.000 857.810 300.000 ;
    END
  END cm_mem_ctrl_out[31]
  PIN cm_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 296.000 757.530 300.000 ;
    END
  END cm_mem_ctrl_out[3]
  PIN cm_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 296.000 761.210 300.000 ;
    END
  END cm_mem_ctrl_out[4]
  PIN cm_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 296.000 764.430 300.000 ;
    END
  END cm_mem_ctrl_out[5]
  PIN cm_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 296.000 768.110 300.000 ;
    END
  END cm_mem_ctrl_out[6]
  PIN cm_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 296.000 771.790 300.000 ;
    END
  END cm_mem_ctrl_out[7]
  PIN cm_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 296.000 775.470 300.000 ;
    END
  END cm_mem_ctrl_out[8]
  PIN cm_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 296.000 779.150 300.000 ;
    END
  END cm_mem_ctrl_out[9]
  PIN cm_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 296.000 861.490 300.000 ;
    END
  END cm_mem_ctrl_req
  PIN cm_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 296.000 864.710 300.000 ;
    END
  END cm_mem_ctrl_vld
  PIN cm_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 296.000 868.390 300.000 ;
    END
  END cm_mem_ctrl_we
  PIN cm_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END cm_sram0_csb0
  PIN cm_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 0.000 813.650 4.000 ;
    END
  END cm_sram0_dout0[0]
  PIN cm_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 0.000 835.730 4.000 ;
    END
  END cm_sram0_dout0[10]
  PIN cm_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 0.000 838.030 4.000 ;
    END
  END cm_sram0_dout0[11]
  PIN cm_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END cm_sram0_dout0[12]
  PIN cm_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END cm_sram0_dout0[13]
  PIN cm_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 0.000 844.470 4.000 ;
    END
  END cm_sram0_dout0[14]
  PIN cm_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 0.000 846.770 4.000 ;
    END
  END cm_sram0_dout0[15]
  PIN cm_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END cm_sram0_dout0[16]
  PIN cm_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 0.000 850.910 4.000 ;
    END
  END cm_sram0_dout0[17]
  PIN cm_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END cm_sram0_dout0[18]
  PIN cm_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.230 0.000 855.510 4.000 ;
    END
  END cm_sram0_dout0[19]
  PIN cm_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 4.000 ;
    END
  END cm_sram0_dout0[1]
  PIN cm_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.530 0.000 857.810 4.000 ;
    END
  END cm_sram0_dout0[20]
  PIN cm_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 0.000 859.650 4.000 ;
    END
  END cm_sram0_dout0[21]
  PIN cm_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END cm_sram0_dout0[22]
  PIN cm_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 4.000 ;
    END
  END cm_sram0_dout0[23]
  PIN cm_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END cm_sram0_dout0[24]
  PIN cm_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 0.000 868.850 4.000 ;
    END
  END cm_sram0_dout0[25]
  PIN cm_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END cm_sram0_dout0[26]
  PIN cm_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END cm_sram0_dout0[27]
  PIN cm_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END cm_sram0_dout0[28]
  PIN cm_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 0.000 877.590 4.000 ;
    END
  END cm_sram0_dout0[29]
  PIN cm_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END cm_sram0_dout0[2]
  PIN cm_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END cm_sram0_dout0[30]
  PIN cm_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END cm_sram0_dout0[31]
  PIN cm_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END cm_sram0_dout0[3]
  PIN cm_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END cm_sram0_dout0[4]
  PIN cm_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END cm_sram0_dout0[5]
  PIN cm_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 0.000 826.990 4.000 ;
    END
  END cm_sram0_dout0[6]
  PIN cm_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 4.000 ;
    END
  END cm_sram0_dout0[7]
  PIN cm_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END cm_sram0_dout0[8]
  PIN cm_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END cm_sram0_dout0[9]
  PIN cm_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.750 0.000 884.030 4.000 ;
    END
  END cm_sram0_web0
  PIN cm_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 0.000 886.330 4.000 ;
    END
  END cm_sram1_csb0
  PIN cm_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END cm_sram1_dout0[0]
  PIN cm_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END cm_sram1_dout0[10]
  PIN cm_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 0.000 912.550 4.000 ;
    END
  END cm_sram1_dout0[11]
  PIN cm_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END cm_sram1_dout0[12]
  PIN cm_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END cm_sram1_dout0[13]
  PIN cm_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.170 0.000 919.450 4.000 ;
    END
  END cm_sram1_dout0[14]
  PIN cm_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 0.000 921.750 4.000 ;
    END
  END cm_sram1_dout0[15]
  PIN cm_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.310 0.000 923.590 4.000 ;
    END
  END cm_sram1_dout0[16]
  PIN cm_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 4.000 ;
    END
  END cm_sram1_dout0[17]
  PIN cm_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END cm_sram1_dout0[18]
  PIN cm_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 0.000 930.490 4.000 ;
    END
  END cm_sram1_dout0[19]
  PIN cm_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.650 0.000 890.930 4.000 ;
    END
  END cm_sram1_dout0[1]
  PIN cm_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END cm_sram1_dout0[20]
  PIN cm_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 0.000 934.630 4.000 ;
    END
  END cm_sram1_dout0[21]
  PIN cm_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END cm_sram1_dout0[22]
  PIN cm_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 0.000 939.230 4.000 ;
    END
  END cm_sram1_dout0[23]
  PIN cm_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 4.000 ;
    END
  END cm_sram1_dout0[24]
  PIN cm_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 0.000 943.370 4.000 ;
    END
  END cm_sram1_dout0[25]
  PIN cm_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END cm_sram1_dout0[26]
  PIN cm_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 0.000 947.970 4.000 ;
    END
  END cm_sram1_dout0[27]
  PIN cm_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END cm_sram1_dout0[28]
  PIN cm_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 0.000 952.570 4.000 ;
    END
  END cm_sram1_dout0[29]
  PIN cm_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 4.000 ;
    END
  END cm_sram1_dout0[2]
  PIN cm_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END cm_sram1_dout0[30]
  PIN cm_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END cm_sram1_dout0[31]
  PIN cm_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 0.000 895.070 4.000 ;
    END
  END cm_sram1_dout0[3]
  PIN cm_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END cm_sram1_dout0[4]
  PIN cm_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END cm_sram1_dout0[5]
  PIN cm_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END cm_sram1_dout0[6]
  PIN cm_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END cm_sram1_dout0[7]
  PIN cm_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.830 0.000 906.110 4.000 ;
    END
  END cm_sram1_dout0[8]
  PIN cm_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END cm_sram1_dout0[9]
  PIN cm_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END cm_sram1_web0
  PIN cm_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 0.000 961.310 4.000 ;
    END
  END cm_sram2_csb0
  PIN cm_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END cm_sram2_dout0[0]
  PIN cm_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END cm_sram2_dout0[10]
  PIN cm_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END cm_sram2_dout0[11]
  PIN cm_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 0.000 989.830 4.000 ;
    END
  END cm_sram2_dout0[12]
  PIN cm_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END cm_sram2_dout0[13]
  PIN cm_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 0.000 994.430 4.000 ;
    END
  END cm_sram2_dout0[14]
  PIN cm_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 4.000 ;
    END
  END cm_sram2_dout0[15]
  PIN cm_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END cm_sram2_dout0[16]
  PIN cm_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 4.000 ;
    END
  END cm_sram2_dout0[17]
  PIN cm_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 0.000 1003.170 4.000 ;
    END
  END cm_sram2_dout0[18]
  PIN cm_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END cm_sram2_dout0[19]
  PIN cm_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END cm_sram2_dout0[1]
  PIN cm_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.030 0.000 1007.310 4.000 ;
    END
  END cm_sram2_dout0[20]
  PIN cm_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 4.000 ;
    END
  END cm_sram2_dout0[21]
  PIN cm_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 0.000 1011.910 4.000 ;
    END
  END cm_sram2_dout0[22]
  PIN cm_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 0.000 1014.210 4.000 ;
    END
  END cm_sram2_dout0[23]
  PIN cm_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 0.000 1016.050 4.000 ;
    END
  END cm_sram2_dout0[24]
  PIN cm_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 0.000 1018.350 4.000 ;
    END
  END cm_sram2_dout0[25]
  PIN cm_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 4.000 ;
    END
  END cm_sram2_dout0[26]
  PIN cm_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.670 0.000 1022.950 4.000 ;
    END
  END cm_sram2_dout0[27]
  PIN cm_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 0.000 1025.250 4.000 ;
    END
  END cm_sram2_dout0[28]
  PIN cm_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.810 0.000 1027.090 4.000 ;
    END
  END cm_sram2_dout0[29]
  PIN cm_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 4.000 ;
    END
  END cm_sram2_dout0[2]
  PIN cm_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END cm_sram2_dout0[30]
  PIN cm_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.410 0.000 1031.690 4.000 ;
    END
  END cm_sram2_dout0[31]
  PIN cm_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 0.000 970.050 4.000 ;
    END
  END cm_sram2_dout0[3]
  PIN cm_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END cm_sram2_dout0[4]
  PIN cm_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.910 0.000 974.190 4.000 ;
    END
  END cm_sram2_dout0[5]
  PIN cm_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END cm_sram2_dout0[6]
  PIN cm_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.510 0.000 978.790 4.000 ;
    END
  END cm_sram2_dout0[7]
  PIN cm_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 4.000 ;
    END
  END cm_sram2_dout0[8]
  PIN cm_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 0.000 983.390 4.000 ;
    END
  END cm_sram2_dout0[9]
  PIN cm_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END cm_sram2_web0
  PIN cm_sram3_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 0.000 1035.830 4.000 ;
    END
  END cm_sram3_csb0
  PIN cm_sram3_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 0.000 1038.130 4.000 ;
    END
  END cm_sram3_dout0[0]
  PIN cm_sram3_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 0.000 1060.210 4.000 ;
    END
  END cm_sram3_dout0[10]
  PIN cm_sram3_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 0.000 1062.510 4.000 ;
    END
  END cm_sram3_dout0[11]
  PIN cm_sram3_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END cm_sram3_dout0[12]
  PIN cm_sram3_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 0.000 1066.650 4.000 ;
    END
  END cm_sram3_dout0[13]
  PIN cm_sram3_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.670 0.000 1068.950 4.000 ;
    END
  END cm_sram3_dout0[14]
  PIN cm_sram3_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.970 0.000 1071.250 4.000 ;
    END
  END cm_sram3_dout0[15]
  PIN cm_sram3_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END cm_sram3_dout0[16]
  PIN cm_sram3_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END cm_sram3_dout0[17]
  PIN cm_sram3_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END cm_sram3_dout0[18]
  PIN cm_sram3_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 4.000 ;
    END
  END cm_sram3_dout0[19]
  PIN cm_sram3_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END cm_sram3_dout0[1]
  PIN cm_sram3_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END cm_sram3_dout0[20]
  PIN cm_sram3_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 0.000 1084.590 4.000 ;
    END
  END cm_sram3_dout0[21]
  PIN cm_sram3_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 0.000 1086.890 4.000 ;
    END
  END cm_sram3_dout0[22]
  PIN cm_sram3_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END cm_sram3_dout0[23]
  PIN cm_sram3_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 0.000 1091.030 4.000 ;
    END
  END cm_sram3_dout0[24]
  PIN cm_sram3_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 0.000 1093.330 4.000 ;
    END
  END cm_sram3_dout0[25]
  PIN cm_sram3_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 0.000 1095.630 4.000 ;
    END
  END cm_sram3_dout0[26]
  PIN cm_sram3_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.650 0.000 1097.930 4.000 ;
    END
  END cm_sram3_dout0[27]
  PIN cm_sram3_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.490 0.000 1099.770 4.000 ;
    END
  END cm_sram3_dout0[28]
  PIN cm_sram3_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 0.000 1102.070 4.000 ;
    END
  END cm_sram3_dout0[29]
  PIN cm_sram3_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 4.000 ;
    END
  END cm_sram3_dout0[2]
  PIN cm_sram3_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END cm_sram3_dout0[30]
  PIN cm_sram3_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.390 0.000 1106.670 4.000 ;
    END
  END cm_sram3_dout0[31]
  PIN cm_sram3_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 0.000 1045.030 4.000 ;
    END
  END cm_sram3_dout0[3]
  PIN cm_sram3_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END cm_sram3_dout0[4]
  PIN cm_sram3_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 0.000 1049.170 4.000 ;
    END
  END cm_sram3_dout0[5]
  PIN cm_sram3_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 0.000 1051.470 4.000 ;
    END
  END cm_sram3_dout0[6]
  PIN cm_sram3_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.490 0.000 1053.770 4.000 ;
    END
  END cm_sram3_dout0[7]
  PIN cm_sram3_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END cm_sram3_dout0[8]
  PIN cm_sram3_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.630 0.000 1057.910 4.000 ;
    END
  END cm_sram3_dout0[9]
  PIN cm_sram3_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 4.000 ;
    END
  END cm_sram3_web0
  PIN cm_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.530 0.000 1110.810 4.000 ;
    END
  END cm_sram_comm_addr0[0]
  PIN cm_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.830 0.000 1113.110 4.000 ;
    END
  END cm_sram_comm_addr0[1]
  PIN cm_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 0.000 1115.410 4.000 ;
    END
  END cm_sram_comm_addr0[2]
  PIN cm_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END cm_sram_comm_addr0[3]
  PIN cm_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.270 0.000 1119.550 4.000 ;
    END
  END cm_sram_comm_addr0[4]
  PIN cm_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.570 0.000 1121.850 4.000 ;
    END
  END cm_sram_comm_addr0[5]
  PIN cm_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END cm_sram_comm_addr0[6]
  PIN cm_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.170 0.000 1126.450 4.000 ;
    END
  END cm_sram_comm_addr0[7]
  PIN cm_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 0.000 1128.750 4.000 ;
    END
  END cm_sram_comm_addr0[8]
  PIN cm_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END cm_sram_comm_din0[0]
  PIN cm_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.390 0.000 1152.670 4.000 ;
    END
  END cm_sram_comm_din0[10]
  PIN cm_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 0.000 1154.970 4.000 ;
    END
  END cm_sram_comm_din0[11]
  PIN cm_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 0.000 1157.270 4.000 ;
    END
  END cm_sram_comm_din0[12]
  PIN cm_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END cm_sram_comm_din0[13]
  PIN cm_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.130 0.000 1161.410 4.000 ;
    END
  END cm_sram_comm_din0[14]
  PIN cm_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.430 0.000 1163.710 4.000 ;
    END
  END cm_sram_comm_din0[15]
  PIN cm_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END cm_sram_comm_din0[16]
  PIN cm_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 0.000 1168.310 4.000 ;
    END
  END cm_sram_comm_din0[17]
  PIN cm_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 0.000 1170.150 4.000 ;
    END
  END cm_sram_comm_din0[18]
  PIN cm_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END cm_sram_comm_din0[19]
  PIN cm_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.610 0.000 1132.890 4.000 ;
    END
  END cm_sram_comm_din0[1]
  PIN cm_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.470 0.000 1174.750 4.000 ;
    END
  END cm_sram_comm_din0[20]
  PIN cm_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END cm_sram_comm_din0[21]
  PIN cm_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.070 0.000 1179.350 4.000 ;
    END
  END cm_sram_comm_din0[22]
  PIN cm_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END cm_sram_comm_din0[23]
  PIN cm_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 0.000 1183.490 4.000 ;
    END
  END cm_sram_comm_din0[24]
  PIN cm_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 0.000 1185.790 4.000 ;
    END
  END cm_sram_comm_din0[25]
  PIN cm_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END cm_sram_comm_din0[26]
  PIN cm_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 0.000 1190.390 4.000 ;
    END
  END cm_sram_comm_din0[27]
  PIN cm_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 4.000 ;
    END
  END cm_sram_comm_din0[28]
  PIN cm_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END cm_sram_comm_din0[29]
  PIN cm_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END cm_sram_comm_din0[2]
  PIN cm_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.550 0.000 1196.830 4.000 ;
    END
  END cm_sram_comm_din0[30]
  PIN cm_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.850 0.000 1199.130 4.000 ;
    END
  END cm_sram_comm_din0[31]
  PIN cm_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END cm_sram_comm_din0[3]
  PIN cm_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.050 0.000 1139.330 4.000 ;
    END
  END cm_sram_comm_din0[4]
  PIN cm_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END cm_sram_comm_din0[5]
  PIN cm_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END cm_sram_comm_din0[6]
  PIN cm_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 0.000 1146.230 4.000 ;
    END
  END cm_sram_comm_din0[7]
  PIN cm_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 0.000 1148.530 4.000 ;
    END
  END cm_sram_comm_din0[8]
  PIN cm_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 4.000 ;
    END
  END cm_sram_comm_din0[9]
  PIN ct_mem_ctrl_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 296.000 291.550 300.000 ;
    END
  END ct_mem_ctrl_addr[0]
  PIN ct_mem_ctrl_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 296.000 327.430 300.000 ;
    END
  END ct_mem_ctrl_addr[10]
  PIN ct_mem_ctrl_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 296.000 331.110 300.000 ;
    END
  END ct_mem_ctrl_addr[11]
  PIN ct_mem_ctrl_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 296.000 334.790 300.000 ;
    END
  END ct_mem_ctrl_addr[12]
  PIN ct_mem_ctrl_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 296.000 338.470 300.000 ;
    END
  END ct_mem_ctrl_addr[13]
  PIN ct_mem_ctrl_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 296.000 295.230 300.000 ;
    END
  END ct_mem_ctrl_addr[1]
  PIN ct_mem_ctrl_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 296.000 298.910 300.000 ;
    END
  END ct_mem_ctrl_addr[2]
  PIN ct_mem_ctrl_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 296.000 302.590 300.000 ;
    END
  END ct_mem_ctrl_addr[3]
  PIN ct_mem_ctrl_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 296.000 305.810 300.000 ;
    END
  END ct_mem_ctrl_addr[4]
  PIN ct_mem_ctrl_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 296.000 309.490 300.000 ;
    END
  END ct_mem_ctrl_addr[5]
  PIN ct_mem_ctrl_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 296.000 313.170 300.000 ;
    END
  END ct_mem_ctrl_addr[6]
  PIN ct_mem_ctrl_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 296.000 316.850 300.000 ;
    END
  END ct_mem_ctrl_addr[7]
  PIN ct_mem_ctrl_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 296.000 320.530 300.000 ;
    END
  END ct_mem_ctrl_addr[8]
  PIN ct_mem_ctrl_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 296.000 323.750 300.000 ;
    END
  END ct_mem_ctrl_addr[9]
  PIN ct_mem_ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 296.000 341.690 300.000 ;
    END
  END ct_mem_ctrl_in[0]
  PIN ct_mem_ctrl_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 296.000 377.570 300.000 ;
    END
  END ct_mem_ctrl_in[10]
  PIN ct_mem_ctrl_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 296.000 381.250 300.000 ;
    END
  END ct_mem_ctrl_in[11]
  PIN ct_mem_ctrl_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 296.000 384.930 300.000 ;
    END
  END ct_mem_ctrl_in[12]
  PIN ct_mem_ctrl_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 296.000 388.610 300.000 ;
    END
  END ct_mem_ctrl_in[13]
  PIN ct_mem_ctrl_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 296.000 391.830 300.000 ;
    END
  END ct_mem_ctrl_in[14]
  PIN ct_mem_ctrl_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 296.000 395.510 300.000 ;
    END
  END ct_mem_ctrl_in[15]
  PIN ct_mem_ctrl_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 296.000 399.190 300.000 ;
    END
  END ct_mem_ctrl_in[16]
  PIN ct_mem_ctrl_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 296.000 402.870 300.000 ;
    END
  END ct_mem_ctrl_in[17]
  PIN ct_mem_ctrl_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 296.000 406.550 300.000 ;
    END
  END ct_mem_ctrl_in[18]
  PIN ct_mem_ctrl_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 296.000 409.770 300.000 ;
    END
  END ct_mem_ctrl_in[19]
  PIN ct_mem_ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 296.000 345.370 300.000 ;
    END
  END ct_mem_ctrl_in[1]
  PIN ct_mem_ctrl_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 296.000 413.450 300.000 ;
    END
  END ct_mem_ctrl_in[20]
  PIN ct_mem_ctrl_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 296.000 417.130 300.000 ;
    END
  END ct_mem_ctrl_in[21]
  PIN ct_mem_ctrl_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 296.000 420.810 300.000 ;
    END
  END ct_mem_ctrl_in[22]
  PIN ct_mem_ctrl_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 296.000 424.030 300.000 ;
    END
  END ct_mem_ctrl_in[23]
  PIN ct_mem_ctrl_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 296.000 427.710 300.000 ;
    END
  END ct_mem_ctrl_in[24]
  PIN ct_mem_ctrl_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 296.000 431.390 300.000 ;
    END
  END ct_mem_ctrl_in[25]
  PIN ct_mem_ctrl_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 296.000 435.070 300.000 ;
    END
  END ct_mem_ctrl_in[26]
  PIN ct_mem_ctrl_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 296.000 438.750 300.000 ;
    END
  END ct_mem_ctrl_in[27]
  PIN ct_mem_ctrl_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 296.000 441.970 300.000 ;
    END
  END ct_mem_ctrl_in[28]
  PIN ct_mem_ctrl_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 296.000 445.650 300.000 ;
    END
  END ct_mem_ctrl_in[29]
  PIN ct_mem_ctrl_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 296.000 349.050 300.000 ;
    END
  END ct_mem_ctrl_in[2]
  PIN ct_mem_ctrl_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 296.000 449.330 300.000 ;
    END
  END ct_mem_ctrl_in[30]
  PIN ct_mem_ctrl_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 296.000 453.010 300.000 ;
    END
  END ct_mem_ctrl_in[31]
  PIN ct_mem_ctrl_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 296.000 352.730 300.000 ;
    END
  END ct_mem_ctrl_in[3]
  PIN ct_mem_ctrl_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 296.000 356.410 300.000 ;
    END
  END ct_mem_ctrl_in[4]
  PIN ct_mem_ctrl_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 296.000 359.630 300.000 ;
    END
  END ct_mem_ctrl_in[5]
  PIN ct_mem_ctrl_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 296.000 363.310 300.000 ;
    END
  END ct_mem_ctrl_in[6]
  PIN ct_mem_ctrl_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 296.000 366.990 300.000 ;
    END
  END ct_mem_ctrl_in[7]
  PIN ct_mem_ctrl_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 296.000 370.670 300.000 ;
    END
  END ct_mem_ctrl_in[8]
  PIN ct_mem_ctrl_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 296.000 373.890 300.000 ;
    END
  END ct_mem_ctrl_in[9]
  PIN ct_mem_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 296.000 456.690 300.000 ;
    END
  END ct_mem_ctrl_out[0]
  PIN ct_mem_ctrl_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 296.000 492.110 300.000 ;
    END
  END ct_mem_ctrl_out[10]
  PIN ct_mem_ctrl_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 296.000 495.790 300.000 ;
    END
  END ct_mem_ctrl_out[11]
  PIN ct_mem_ctrl_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 296.000 499.470 300.000 ;
    END
  END ct_mem_ctrl_out[12]
  PIN ct_mem_ctrl_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 296.000 503.150 300.000 ;
    END
  END ct_mem_ctrl_out[13]
  PIN ct_mem_ctrl_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 296.000 506.830 300.000 ;
    END
  END ct_mem_ctrl_out[14]
  PIN ct_mem_ctrl_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 296.000 510.050 300.000 ;
    END
  END ct_mem_ctrl_out[15]
  PIN ct_mem_ctrl_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 296.000 513.730 300.000 ;
    END
  END ct_mem_ctrl_out[16]
  PIN ct_mem_ctrl_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 296.000 517.410 300.000 ;
    END
  END ct_mem_ctrl_out[17]
  PIN ct_mem_ctrl_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 296.000 521.090 300.000 ;
    END
  END ct_mem_ctrl_out[18]
  PIN ct_mem_ctrl_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 296.000 524.770 300.000 ;
    END
  END ct_mem_ctrl_out[19]
  PIN ct_mem_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 296.000 459.910 300.000 ;
    END
  END ct_mem_ctrl_out[1]
  PIN ct_mem_ctrl_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 296.000 527.990 300.000 ;
    END
  END ct_mem_ctrl_out[20]
  PIN ct_mem_ctrl_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 296.000 531.670 300.000 ;
    END
  END ct_mem_ctrl_out[21]
  PIN ct_mem_ctrl_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 296.000 535.350 300.000 ;
    END
  END ct_mem_ctrl_out[22]
  PIN ct_mem_ctrl_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 296.000 539.030 300.000 ;
    END
  END ct_mem_ctrl_out[23]
  PIN ct_mem_ctrl_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 296.000 542.250 300.000 ;
    END
  END ct_mem_ctrl_out[24]
  PIN ct_mem_ctrl_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 296.000 545.930 300.000 ;
    END
  END ct_mem_ctrl_out[25]
  PIN ct_mem_ctrl_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 296.000 549.610 300.000 ;
    END
  END ct_mem_ctrl_out[26]
  PIN ct_mem_ctrl_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 296.000 553.290 300.000 ;
    END
  END ct_mem_ctrl_out[27]
  PIN ct_mem_ctrl_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 296.000 556.970 300.000 ;
    END
  END ct_mem_ctrl_out[28]
  PIN ct_mem_ctrl_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 296.000 560.190 300.000 ;
    END
  END ct_mem_ctrl_out[29]
  PIN ct_mem_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 296.000 463.590 300.000 ;
    END
  END ct_mem_ctrl_out[2]
  PIN ct_mem_ctrl_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 296.000 563.870 300.000 ;
    END
  END ct_mem_ctrl_out[30]
  PIN ct_mem_ctrl_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 296.000 567.550 300.000 ;
    END
  END ct_mem_ctrl_out[31]
  PIN ct_mem_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 296.000 467.270 300.000 ;
    END
  END ct_mem_ctrl_out[3]
  PIN ct_mem_ctrl_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 296.000 470.950 300.000 ;
    END
  END ct_mem_ctrl_out[4]
  PIN ct_mem_ctrl_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 296.000 474.630 300.000 ;
    END
  END ct_mem_ctrl_out[5]
  PIN ct_mem_ctrl_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 296.000 477.850 300.000 ;
    END
  END ct_mem_ctrl_out[6]
  PIN ct_mem_ctrl_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 296.000 481.530 300.000 ;
    END
  END ct_mem_ctrl_out[7]
  PIN ct_mem_ctrl_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 296.000 485.210 300.000 ;
    END
  END ct_mem_ctrl_out[8]
  PIN ct_mem_ctrl_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 296.000 488.890 300.000 ;
    END
  END ct_mem_ctrl_out[9]
  PIN ct_mem_ctrl_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 296.000 571.230 300.000 ;
    END
  END ct_mem_ctrl_req
  PIN ct_mem_ctrl_vld
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 296.000 574.910 300.000 ;
    END
  END ct_mem_ctrl_vld
  PIN ct_mem_ctrl_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 296.000 578.130 300.000 ;
    END
  END ct_mem_ctrl_we
  PIN ct_sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END ct_sram0_csb0
  PIN ct_sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END ct_sram0_dout0[0]
  PIN ct_sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END ct_sram0_dout0[10]
  PIN ct_sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END ct_sram0_dout0[11]
  PIN ct_sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END ct_sram0_dout0[12]
  PIN ct_sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END ct_sram0_dout0[13]
  PIN ct_sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END ct_sram0_dout0[14]
  PIN ct_sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END ct_sram0_dout0[15]
  PIN ct_sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END ct_sram0_dout0[16]
  PIN ct_sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END ct_sram0_dout0[17]
  PIN ct_sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END ct_sram0_dout0[18]
  PIN ct_sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END ct_sram0_dout0[19]
  PIN ct_sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END ct_sram0_dout0[1]
  PIN ct_sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END ct_sram0_dout0[20]
  PIN ct_sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END ct_sram0_dout0[21]
  PIN ct_sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END ct_sram0_dout0[22]
  PIN ct_sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END ct_sram0_dout0[23]
  PIN ct_sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END ct_sram0_dout0[24]
  PIN ct_sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END ct_sram0_dout0[25]
  PIN ct_sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END ct_sram0_dout0[26]
  PIN ct_sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END ct_sram0_dout0[27]
  PIN ct_sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END ct_sram0_dout0[28]
  PIN ct_sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END ct_sram0_dout0[29]
  PIN ct_sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END ct_sram0_dout0[2]
  PIN ct_sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END ct_sram0_dout0[30]
  PIN ct_sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END ct_sram0_dout0[31]
  PIN ct_sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END ct_sram0_dout0[3]
  PIN ct_sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END ct_sram0_dout0[4]
  PIN ct_sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END ct_sram0_dout0[5]
  PIN ct_sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END ct_sram0_dout0[6]
  PIN ct_sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END ct_sram0_dout0[7]
  PIN ct_sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END ct_sram0_dout0[8]
  PIN ct_sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END ct_sram0_dout0[9]
  PIN ct_sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END ct_sram0_web0
  PIN ct_sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END ct_sram1_csb0
  PIN ct_sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END ct_sram1_dout0[0]
  PIN ct_sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END ct_sram1_dout0[10]
  PIN ct_sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END ct_sram1_dout0[11]
  PIN ct_sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END ct_sram1_dout0[12]
  PIN ct_sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END ct_sram1_dout0[13]
  PIN ct_sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END ct_sram1_dout0[14]
  PIN ct_sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END ct_sram1_dout0[15]
  PIN ct_sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END ct_sram1_dout0[16]
  PIN ct_sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END ct_sram1_dout0[17]
  PIN ct_sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END ct_sram1_dout0[18]
  PIN ct_sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END ct_sram1_dout0[19]
  PIN ct_sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END ct_sram1_dout0[1]
  PIN ct_sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END ct_sram1_dout0[20]
  PIN ct_sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END ct_sram1_dout0[21]
  PIN ct_sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END ct_sram1_dout0[22]
  PIN ct_sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END ct_sram1_dout0[23]
  PIN ct_sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END ct_sram1_dout0[24]
  PIN ct_sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END ct_sram1_dout0[25]
  PIN ct_sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END ct_sram1_dout0[26]
  PIN ct_sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END ct_sram1_dout0[27]
  PIN ct_sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END ct_sram1_dout0[28]
  PIN ct_sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END ct_sram1_dout0[29]
  PIN ct_sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END ct_sram1_dout0[2]
  PIN ct_sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END ct_sram1_dout0[30]
  PIN ct_sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END ct_sram1_dout0[31]
  PIN ct_sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END ct_sram1_dout0[3]
  PIN ct_sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END ct_sram1_dout0[4]
  PIN ct_sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END ct_sram1_dout0[5]
  PIN ct_sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END ct_sram1_dout0[6]
  PIN ct_sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END ct_sram1_dout0[7]
  PIN ct_sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END ct_sram1_dout0[8]
  PIN ct_sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END ct_sram1_dout0[9]
  PIN ct_sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END ct_sram1_web0
  PIN ct_sram2_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END ct_sram2_csb0
  PIN ct_sram2_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END ct_sram2_dout0[0]
  PIN ct_sram2_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END ct_sram2_dout0[10]
  PIN ct_sram2_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END ct_sram2_dout0[11]
  PIN ct_sram2_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END ct_sram2_dout0[12]
  PIN ct_sram2_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END ct_sram2_dout0[13]
  PIN ct_sram2_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END ct_sram2_dout0[14]
  PIN ct_sram2_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END ct_sram2_dout0[15]
  PIN ct_sram2_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END ct_sram2_dout0[16]
  PIN ct_sram2_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END ct_sram2_dout0[17]
  PIN ct_sram2_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END ct_sram2_dout0[18]
  PIN ct_sram2_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END ct_sram2_dout0[19]
  PIN ct_sram2_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END ct_sram2_dout0[1]
  PIN ct_sram2_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END ct_sram2_dout0[20]
  PIN ct_sram2_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END ct_sram2_dout0[21]
  PIN ct_sram2_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END ct_sram2_dout0[22]
  PIN ct_sram2_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END ct_sram2_dout0[23]
  PIN ct_sram2_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END ct_sram2_dout0[24]
  PIN ct_sram2_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END ct_sram2_dout0[25]
  PIN ct_sram2_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END ct_sram2_dout0[26]
  PIN ct_sram2_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END ct_sram2_dout0[27]
  PIN ct_sram2_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END ct_sram2_dout0[28]
  PIN ct_sram2_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END ct_sram2_dout0[29]
  PIN ct_sram2_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END ct_sram2_dout0[2]
  PIN ct_sram2_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END ct_sram2_dout0[30]
  PIN ct_sram2_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END ct_sram2_dout0[31]
  PIN ct_sram2_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END ct_sram2_dout0[3]
  PIN ct_sram2_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END ct_sram2_dout0[4]
  PIN ct_sram2_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END ct_sram2_dout0[5]
  PIN ct_sram2_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END ct_sram2_dout0[6]
  PIN ct_sram2_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END ct_sram2_dout0[7]
  PIN ct_sram2_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END ct_sram2_dout0[8]
  PIN ct_sram2_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END ct_sram2_dout0[9]
  PIN ct_sram2_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END ct_sram2_web0
  PIN ct_sram3_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END ct_sram3_csb0
  PIN ct_sram3_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END ct_sram3_dout0[0]
  PIN ct_sram3_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END ct_sram3_dout0[10]
  PIN ct_sram3_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END ct_sram3_dout0[11]
  PIN ct_sram3_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END ct_sram3_dout0[12]
  PIN ct_sram3_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 0.000 602.050 4.000 ;
    END
  END ct_sram3_dout0[13]
  PIN ct_sram3_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END ct_sram3_dout0[14]
  PIN ct_sram3_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END ct_sram3_dout0[15]
  PIN ct_sram3_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END ct_sram3_dout0[16]
  PIN ct_sram3_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END ct_sram3_dout0[17]
  PIN ct_sram3_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END ct_sram3_dout0[18]
  PIN ct_sram3_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END ct_sram3_dout0[19]
  PIN ct_sram3_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END ct_sram3_dout0[1]
  PIN ct_sram3_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END ct_sram3_dout0[20]
  PIN ct_sram3_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END ct_sram3_dout0[21]
  PIN ct_sram3_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END ct_sram3_dout0[22]
  PIN ct_sram3_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END ct_sram3_dout0[23]
  PIN ct_sram3_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END ct_sram3_dout0[24]
  PIN ct_sram3_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END ct_sram3_dout0[25]
  PIN ct_sram3_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END ct_sram3_dout0[26]
  PIN ct_sram3_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END ct_sram3_dout0[27]
  PIN ct_sram3_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END ct_sram3_dout0[28]
  PIN ct_sram3_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END ct_sram3_dout0[29]
  PIN ct_sram3_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END ct_sram3_dout0[2]
  PIN ct_sram3_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END ct_sram3_dout0[30]
  PIN ct_sram3_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 4.000 ;
    END
  END ct_sram3_dout0[31]
  PIN ct_sram3_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END ct_sram3_dout0[3]
  PIN ct_sram3_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END ct_sram3_dout0[4]
  PIN ct_sram3_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END ct_sram3_dout0[5]
  PIN ct_sram3_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END ct_sram3_dout0[6]
  PIN ct_sram3_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END ct_sram3_dout0[7]
  PIN ct_sram3_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END ct_sram3_dout0[8]
  PIN ct_sram3_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END ct_sram3_dout0[9]
  PIN ct_sram3_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END ct_sram3_web0
  PIN ct_sram4_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END ct_sram4_csb0
  PIN ct_sram4_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 0.000 648.510 4.000 ;
    END
  END ct_sram4_dout0[0]
  PIN ct_sram4_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END ct_sram4_dout0[10]
  PIN ct_sram4_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END ct_sram4_dout0[11]
  PIN ct_sram4_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END ct_sram4_dout0[12]
  PIN ct_sram4_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END ct_sram4_dout0[13]
  PIN ct_sram4_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END ct_sram4_dout0[14]
  PIN ct_sram4_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END ct_sram4_dout0[15]
  PIN ct_sram4_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END ct_sram4_dout0[16]
  PIN ct_sram4_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END ct_sram4_dout0[17]
  PIN ct_sram4_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END ct_sram4_dout0[18]
  PIN ct_sram4_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END ct_sram4_dout0[19]
  PIN ct_sram4_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END ct_sram4_dout0[1]
  PIN ct_sram4_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END ct_sram4_dout0[20]
  PIN ct_sram4_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END ct_sram4_dout0[21]
  PIN ct_sram4_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END ct_sram4_dout0[22]
  PIN ct_sram4_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END ct_sram4_dout0[23]
  PIN ct_sram4_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 0.000 701.410 4.000 ;
    END
  END ct_sram4_dout0[24]
  PIN ct_sram4_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 0.000 703.710 4.000 ;
    END
  END ct_sram4_dout0[25]
  PIN ct_sram4_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END ct_sram4_dout0[26]
  PIN ct_sram4_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END ct_sram4_dout0[27]
  PIN ct_sram4_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 0.000 710.150 4.000 ;
    END
  END ct_sram4_dout0[28]
  PIN ct_sram4_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END ct_sram4_dout0[29]
  PIN ct_sram4_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END ct_sram4_dout0[2]
  PIN ct_sram4_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END ct_sram4_dout0[30]
  PIN ct_sram4_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END ct_sram4_dout0[31]
  PIN ct_sram4_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 0.000 654.950 4.000 ;
    END
  END ct_sram4_dout0[3]
  PIN ct_sram4_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END ct_sram4_dout0[4]
  PIN ct_sram4_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 4.000 ;
    END
  END ct_sram4_dout0[5]
  PIN ct_sram4_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END ct_sram4_dout0[6]
  PIN ct_sram4_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END ct_sram4_dout0[7]
  PIN ct_sram4_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END ct_sram4_dout0[8]
  PIN ct_sram4_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END ct_sram4_dout0[9]
  PIN ct_sram4_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END ct_sram4_web0
  PIN ct_sram_comm_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END ct_sram_comm_addr0[0]
  PIN ct_sram_comm_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END ct_sram_comm_addr0[1]
  PIN ct_sram_comm_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END ct_sram_comm_addr0[2]
  PIN ct_sram_comm_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END ct_sram_comm_addr0[3]
  PIN ct_sram_comm_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END ct_sram_comm_addr0[4]
  PIN ct_sram_comm_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END ct_sram_comm_addr0[5]
  PIN ct_sram_comm_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END ct_sram_comm_addr0[6]
  PIN ct_sram_comm_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END ct_sram_comm_addr0[7]
  PIN ct_sram_comm_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END ct_sram_comm_addr0[8]
  PIN ct_sram_comm_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END ct_sram_comm_din0[0]
  PIN ct_sram_comm_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END ct_sram_comm_din0[10]
  PIN ct_sram_comm_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END ct_sram_comm_din0[11]
  PIN ct_sram_comm_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 0.000 767.190 4.000 ;
    END
  END ct_sram_comm_din0[12]
  PIN ct_sram_comm_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END ct_sram_comm_din0[13]
  PIN ct_sram_comm_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END ct_sram_comm_din0[14]
  PIN ct_sram_comm_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END ct_sram_comm_din0[15]
  PIN ct_sram_comm_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END ct_sram_comm_din0[16]
  PIN ct_sram_comm_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END ct_sram_comm_din0[17]
  PIN ct_sram_comm_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END ct_sram_comm_din0[18]
  PIN ct_sram_comm_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END ct_sram_comm_din0[19]
  PIN ct_sram_comm_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 0.000 743.270 4.000 ;
    END
  END ct_sram_comm_din0[1]
  PIN ct_sram_comm_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END ct_sram_comm_din0[20]
  PIN ct_sram_comm_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END ct_sram_comm_din0[21]
  PIN ct_sram_comm_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END ct_sram_comm_din0[22]
  PIN ct_sram_comm_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 4.000 ;
    END
  END ct_sram_comm_din0[23]
  PIN ct_sram_comm_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END ct_sram_comm_din0[24]
  PIN ct_sram_comm_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END ct_sram_comm_din0[25]
  PIN ct_sram_comm_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END ct_sram_comm_din0[26]
  PIN ct_sram_comm_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END ct_sram_comm_din0[27]
  PIN ct_sram_comm_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END ct_sram_comm_din0[28]
  PIN ct_sram_comm_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END ct_sram_comm_din0[29]
  PIN ct_sram_comm_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END ct_sram_comm_din0[2]
  PIN ct_sram_comm_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 0.000 807.210 4.000 ;
    END
  END ct_sram_comm_din0[30]
  PIN ct_sram_comm_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 0.000 809.050 4.000 ;
    END
  END ct_sram_comm_din0[31]
  PIN ct_sram_comm_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END ct_sram_comm_din0[3]
  PIN ct_sram_comm_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END ct_sram_comm_din0[4]
  PIN ct_sram_comm_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 0.000 752.010 4.000 ;
    END
  END ct_sram_comm_din0[5]
  PIN ct_sram_comm_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END ct_sram_comm_din0[6]
  PIN ct_sram_comm_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 4.000 ;
    END
  END ct_sram_comm_din0[7]
  PIN ct_sram_comm_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END ct_sram_comm_din0[8]
  PIN ct_sram_comm_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 4.000 ;
    END
  END ct_sram_comm_din0[9]
  PIN main_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 296.000 872.070 300.000 ;
    END
  END main_mem_addr[0]
  PIN main_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.470 296.000 875.750 300.000 ;
    END
  END main_mem_addr[1]
  PIN main_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 296.000 879.430 300.000 ;
    END
  END main_mem_addr[2]
  PIN main_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 296.000 882.650 300.000 ;
    END
  END main_mem_addr[3]
  PIN main_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 296.000 886.330 300.000 ;
    END
  END main_mem_addr[4]
  PIN main_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 296.000 890.010 300.000 ;
    END
  END main_mem_addr[5]
  PIN main_mem_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 296.000 893.690 300.000 ;
    END
  END main_mem_in[0]
  PIN main_mem_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 296.000 929.570 300.000 ;
    END
  END main_mem_in[10]
  PIN main_mem_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 296.000 932.790 300.000 ;
    END
  END main_mem_in[11]
  PIN main_mem_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 296.000 936.470 300.000 ;
    END
  END main_mem_in[12]
  PIN main_mem_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 296.000 940.150 300.000 ;
    END
  END main_mem_in[13]
  PIN main_mem_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 296.000 943.830 300.000 ;
    END
  END main_mem_in[14]
  PIN main_mem_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 296.000 947.510 300.000 ;
    END
  END main_mem_in[15]
  PIN main_mem_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 296.000 950.730 300.000 ;
    END
  END main_mem_in[16]
  PIN main_mem_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 296.000 954.410 300.000 ;
    END
  END main_mem_in[17]
  PIN main_mem_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 296.000 958.090 300.000 ;
    END
  END main_mem_in[18]
  PIN main_mem_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 296.000 961.770 300.000 ;
    END
  END main_mem_in[19]
  PIN main_mem_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 296.000 897.370 300.000 ;
    END
  END main_mem_in[1]
  PIN main_mem_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 296.000 964.990 300.000 ;
    END
  END main_mem_in[20]
  PIN main_mem_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 296.000 968.670 300.000 ;
    END
  END main_mem_in[21]
  PIN main_mem_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 296.000 972.350 300.000 ;
    END
  END main_mem_in[22]
  PIN main_mem_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 296.000 976.030 300.000 ;
    END
  END main_mem_in[23]
  PIN main_mem_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 296.000 979.710 300.000 ;
    END
  END main_mem_in[24]
  PIN main_mem_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 296.000 982.930 300.000 ;
    END
  END main_mem_in[25]
  PIN main_mem_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 296.000 986.610 300.000 ;
    END
  END main_mem_in[26]
  PIN main_mem_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 296.000 990.290 300.000 ;
    END
  END main_mem_in[27]
  PIN main_mem_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 296.000 993.970 300.000 ;
    END
  END main_mem_in[28]
  PIN main_mem_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.370 296.000 997.650 300.000 ;
    END
  END main_mem_in[29]
  PIN main_mem_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 296.000 900.590 300.000 ;
    END
  END main_mem_in[2]
  PIN main_mem_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 296.000 1000.870 300.000 ;
    END
  END main_mem_in[30]
  PIN main_mem_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.270 296.000 1004.550 300.000 ;
    END
  END main_mem_in[31]
  PIN main_mem_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 296.000 904.270 300.000 ;
    END
  END main_mem_in[3]
  PIN main_mem_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 296.000 907.950 300.000 ;
    END
  END main_mem_in[4]
  PIN main_mem_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 296.000 911.630 300.000 ;
    END
  END main_mem_in[5]
  PIN main_mem_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 296.000 914.850 300.000 ;
    END
  END main_mem_in[6]
  PIN main_mem_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 296.000 918.530 300.000 ;
    END
  END main_mem_in[7]
  PIN main_mem_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 296.000 922.210 300.000 ;
    END
  END main_mem_in[8]
  PIN main_mem_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 296.000 925.890 300.000 ;
    END
  END main_mem_in[9]
  PIN main_mem_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 296.000 1008.230 300.000 ;
    END
  END main_mem_out[0]
  PIN main_mem_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.830 296.000 1044.110 300.000 ;
    END
  END main_mem_out[10]
  PIN main_mem_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 296.000 1047.790 300.000 ;
    END
  END main_mem_out[11]
  PIN main_mem_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 296.000 1051.010 300.000 ;
    END
  END main_mem_out[12]
  PIN main_mem_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 296.000 1054.690 300.000 ;
    END
  END main_mem_out[13]
  PIN main_mem_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 296.000 1058.370 300.000 ;
    END
  END main_mem_out[14]
  PIN main_mem_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 296.000 1062.050 300.000 ;
    END
  END main_mem_out[15]
  PIN main_mem_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 296.000 1065.730 300.000 ;
    END
  END main_mem_out[16]
  PIN main_mem_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.670 296.000 1068.950 300.000 ;
    END
  END main_mem_out[17]
  PIN main_mem_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 296.000 1072.630 300.000 ;
    END
  END main_mem_out[18]
  PIN main_mem_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 296.000 1076.310 300.000 ;
    END
  END main_mem_out[19]
  PIN main_mem_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 296.000 1011.910 300.000 ;
    END
  END main_mem_out[1]
  PIN main_mem_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 296.000 1079.990 300.000 ;
    END
  END main_mem_out[20]
  PIN main_mem_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 296.000 1083.210 300.000 ;
    END
  END main_mem_out[21]
  PIN main_mem_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 296.000 1086.890 300.000 ;
    END
  END main_mem_out[22]
  PIN main_mem_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 296.000 1090.570 300.000 ;
    END
  END main_mem_out[23]
  PIN main_mem_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 296.000 1094.250 300.000 ;
    END
  END main_mem_out[24]
  PIN main_mem_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.650 296.000 1097.930 300.000 ;
    END
  END main_mem_out[25]
  PIN main_mem_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.870 296.000 1101.150 300.000 ;
    END
  END main_mem_out[26]
  PIN main_mem_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 296.000 1104.830 300.000 ;
    END
  END main_mem_out[27]
  PIN main_mem_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 296.000 1108.510 300.000 ;
    END
  END main_mem_out[28]
  PIN main_mem_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 296.000 1112.190 300.000 ;
    END
  END main_mem_out[29]
  PIN main_mem_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.310 296.000 1015.590 300.000 ;
    END
  END main_mem_out[2]
  PIN main_mem_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.590 296.000 1115.870 300.000 ;
    END
  END main_mem_out[30]
  PIN main_mem_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.810 296.000 1119.090 300.000 ;
    END
  END main_mem_out[31]
  PIN main_mem_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 296.000 1018.810 300.000 ;
    END
  END main_mem_out[3]
  PIN main_mem_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 296.000 1022.490 300.000 ;
    END
  END main_mem_out[4]
  PIN main_mem_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.890 296.000 1026.170 300.000 ;
    END
  END main_mem_out[5]
  PIN main_mem_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 296.000 1029.850 300.000 ;
    END
  END main_mem_out[6]
  PIN main_mem_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.790 296.000 1033.070 300.000 ;
    END
  END main_mem_out[7]
  PIN main_mem_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.470 296.000 1036.750 300.000 ;
    END
  END main_mem_out[8]
  PIN main_mem_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 296.000 1040.430 300.000 ;
    END
  END main_mem_out[9]
  PIN main_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.490 296.000 1122.770 300.000 ;
    END
  END main_mem_we
  PIN program_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 187.040 1200.000 187.640 ;
    END
  END program_sel[0]
  PIN program_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 261.840 1200.000 262.440 ;
    END
  END program_sel[1]
  PIN r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 296.000 1172.910 300.000 ;
    END
  END r_data[0]
  PIN r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.310 296.000 1176.590 300.000 ;
    END
  END r_data[1]
  PIN r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.990 296.000 1180.270 300.000 ;
    END
  END r_data[2]
  PIN r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 296.000 1183.950 300.000 ;
    END
  END r_data[3]
  PIN r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 296.000 1187.170 300.000 ;
    END
  END r_data[4]
  PIN r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.570 296.000 1190.850 300.000 ;
    END
  END r_data[5]
  PIN r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 296.000 1194.530 300.000 ;
    END
  END r_data[6]
  PIN r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 296.000 1198.210 300.000 ;
    END
  END r_data[7]
  PIN rd_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.850 296.000 1130.130 300.000 ;
    END
  END rd_uart
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 37.440 1200.000 38.040 ;
    END
  END rst
  PIN rst_asserted
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 112.240 1200.000 112.840 ;
    END
  END rst_asserted
  PIN rx_empty
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 296.000 1169.230 300.000 ;
    END
  END rx_empty
  PIN rx_fifo_flush_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.170 296.000 1126.450 300.000 ;
    END
  END rx_fifo_flush_enable
  PIN sram_const_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END sram_const_addr1[0]
  PIN sram_const_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END sram_const_addr1[1]
  PIN sram_const_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END sram_const_addr1[2]
  PIN sram_const_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END sram_const_addr1[3]
  PIN sram_const_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END sram_const_addr1[4]
  PIN sram_const_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END sram_const_addr1[5]
  PIN sram_const_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END sram_const_addr1[6]
  PIN sram_const_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END sram_const_addr1[7]
  PIN sram_const_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END sram_const_addr1[8]
  PIN sram_const_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END sram_const_csb1
  PIN sram_const_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END sram_const_wmask0[0]
  PIN sram_const_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END sram_const_wmask0[1]
  PIN sram_const_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END sram_const_wmask0[2]
  PIN sram_const_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END sram_const_wmask0[3]
  PIN tx_full
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 296.000 1166.010 300.000 ;
    END
  END tx_full
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 288.560 ;
    END
  END vssd1
  PIN w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 296.000 1137.030 300.000 ;
    END
  END w_data[0]
  PIN w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.430 296.000 1140.710 300.000 ;
    END
  END w_data[1]
  PIN w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.110 296.000 1144.390 300.000 ;
    END
  END w_data[2]
  PIN w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 296.000 1148.070 300.000 ;
    END
  END w_data[3]
  PIN w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.010 296.000 1151.290 300.000 ;
    END
  END w_data[4]
  PIN w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 296.000 1154.970 300.000 ;
    END
  END w_data[5]
  PIN w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.370 296.000 1158.650 300.000 ;
    END
  END w_data[6]
  PIN w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 296.000 1162.330 300.000 ;
    END
  END w_data[7]
  PIN wr_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 296.000 1133.810 300.000 ;
    END
  END wr_uart
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 288.405 ;
      LAYER met1 ;
        RECT 0.990 0.720 1199.150 299.840 ;
      LAYER met2 ;
        RECT 1.020 295.720 1.190 299.870 ;
        RECT 2.030 295.720 4.410 299.870 ;
        RECT 5.250 295.720 8.090 299.870 ;
        RECT 8.930 295.720 11.770 299.870 ;
        RECT 12.610 295.720 15.450 299.870 ;
        RECT 16.290 295.720 18.670 299.870 ;
        RECT 19.510 295.720 22.350 299.870 ;
        RECT 23.190 295.720 26.030 299.870 ;
        RECT 26.870 295.720 29.710 299.870 ;
        RECT 30.550 295.720 33.390 299.870 ;
        RECT 34.230 295.720 36.610 299.870 ;
        RECT 37.450 295.720 40.290 299.870 ;
        RECT 41.130 295.720 43.970 299.870 ;
        RECT 44.810 295.720 47.650 299.870 ;
        RECT 48.490 295.720 51.330 299.870 ;
        RECT 52.170 295.720 54.550 299.870 ;
        RECT 55.390 295.720 58.230 299.870 ;
        RECT 59.070 295.720 61.910 299.870 ;
        RECT 62.750 295.720 65.590 299.870 ;
        RECT 66.430 295.720 68.810 299.870 ;
        RECT 69.650 295.720 72.490 299.870 ;
        RECT 73.330 295.720 76.170 299.870 ;
        RECT 77.010 295.720 79.850 299.870 ;
        RECT 80.690 295.720 83.530 299.870 ;
        RECT 84.370 295.720 86.750 299.870 ;
        RECT 87.590 295.720 90.430 299.870 ;
        RECT 91.270 295.720 94.110 299.870 ;
        RECT 94.950 295.720 97.790 299.870 ;
        RECT 98.630 295.720 101.470 299.870 ;
        RECT 102.310 295.720 104.690 299.870 ;
        RECT 105.530 295.720 108.370 299.870 ;
        RECT 109.210 295.720 112.050 299.870 ;
        RECT 112.890 295.720 115.730 299.870 ;
        RECT 116.570 295.720 119.410 299.870 ;
        RECT 120.250 295.720 122.630 299.870 ;
        RECT 123.470 295.720 126.310 299.870 ;
        RECT 127.150 295.720 129.990 299.870 ;
        RECT 130.830 295.720 133.670 299.870 ;
        RECT 134.510 295.720 136.890 299.870 ;
        RECT 137.730 295.720 140.570 299.870 ;
        RECT 141.410 295.720 144.250 299.870 ;
        RECT 145.090 295.720 147.930 299.870 ;
        RECT 148.770 295.720 151.610 299.870 ;
        RECT 152.450 295.720 154.830 299.870 ;
        RECT 155.670 295.720 158.510 299.870 ;
        RECT 159.350 295.720 162.190 299.870 ;
        RECT 163.030 295.720 165.870 299.870 ;
        RECT 166.710 295.720 169.550 299.870 ;
        RECT 170.390 295.720 172.770 299.870 ;
        RECT 173.610 295.720 176.450 299.870 ;
        RECT 177.290 295.720 180.130 299.870 ;
        RECT 180.970 295.720 183.810 299.870 ;
        RECT 184.650 295.720 187.030 299.870 ;
        RECT 187.870 295.720 190.710 299.870 ;
        RECT 191.550 295.720 194.390 299.870 ;
        RECT 195.230 295.720 198.070 299.870 ;
        RECT 198.910 295.720 201.750 299.870 ;
        RECT 202.590 295.720 204.970 299.870 ;
        RECT 205.810 295.720 208.650 299.870 ;
        RECT 209.490 295.720 212.330 299.870 ;
        RECT 213.170 295.720 216.010 299.870 ;
        RECT 216.850 295.720 219.690 299.870 ;
        RECT 220.530 295.720 222.910 299.870 ;
        RECT 223.750 295.720 226.590 299.870 ;
        RECT 227.430 295.720 230.270 299.870 ;
        RECT 231.110 295.720 233.950 299.870 ;
        RECT 234.790 295.720 237.630 299.870 ;
        RECT 238.470 295.720 240.850 299.870 ;
        RECT 241.690 295.720 244.530 299.870 ;
        RECT 245.370 295.720 248.210 299.870 ;
        RECT 249.050 295.720 251.890 299.870 ;
        RECT 252.730 295.720 255.110 299.870 ;
        RECT 255.950 295.720 258.790 299.870 ;
        RECT 259.630 295.720 262.470 299.870 ;
        RECT 263.310 295.720 266.150 299.870 ;
        RECT 266.990 295.720 269.830 299.870 ;
        RECT 270.670 295.720 273.050 299.870 ;
        RECT 273.890 295.720 276.730 299.870 ;
        RECT 277.570 295.720 280.410 299.870 ;
        RECT 281.250 295.720 284.090 299.870 ;
        RECT 284.930 295.720 287.770 299.870 ;
        RECT 288.610 295.720 290.990 299.870 ;
        RECT 291.830 295.720 294.670 299.870 ;
        RECT 295.510 295.720 298.350 299.870 ;
        RECT 299.190 295.720 302.030 299.870 ;
        RECT 302.870 295.720 305.250 299.870 ;
        RECT 306.090 295.720 308.930 299.870 ;
        RECT 309.770 295.720 312.610 299.870 ;
        RECT 313.450 295.720 316.290 299.870 ;
        RECT 317.130 295.720 319.970 299.870 ;
        RECT 320.810 295.720 323.190 299.870 ;
        RECT 324.030 295.720 326.870 299.870 ;
        RECT 327.710 295.720 330.550 299.870 ;
        RECT 331.390 295.720 334.230 299.870 ;
        RECT 335.070 295.720 337.910 299.870 ;
        RECT 338.750 295.720 341.130 299.870 ;
        RECT 341.970 295.720 344.810 299.870 ;
        RECT 345.650 295.720 348.490 299.870 ;
        RECT 349.330 295.720 352.170 299.870 ;
        RECT 353.010 295.720 355.850 299.870 ;
        RECT 356.690 295.720 359.070 299.870 ;
        RECT 359.910 295.720 362.750 299.870 ;
        RECT 363.590 295.720 366.430 299.870 ;
        RECT 367.270 295.720 370.110 299.870 ;
        RECT 370.950 295.720 373.330 299.870 ;
        RECT 374.170 295.720 377.010 299.870 ;
        RECT 377.850 295.720 380.690 299.870 ;
        RECT 381.530 295.720 384.370 299.870 ;
        RECT 385.210 295.720 388.050 299.870 ;
        RECT 388.890 295.720 391.270 299.870 ;
        RECT 392.110 295.720 394.950 299.870 ;
        RECT 395.790 295.720 398.630 299.870 ;
        RECT 399.470 295.720 402.310 299.870 ;
        RECT 403.150 295.720 405.990 299.870 ;
        RECT 406.830 295.720 409.210 299.870 ;
        RECT 410.050 295.720 412.890 299.870 ;
        RECT 413.730 295.720 416.570 299.870 ;
        RECT 417.410 295.720 420.250 299.870 ;
        RECT 421.090 295.720 423.470 299.870 ;
        RECT 424.310 295.720 427.150 299.870 ;
        RECT 427.990 295.720 430.830 299.870 ;
        RECT 431.670 295.720 434.510 299.870 ;
        RECT 435.350 295.720 438.190 299.870 ;
        RECT 439.030 295.720 441.410 299.870 ;
        RECT 442.250 295.720 445.090 299.870 ;
        RECT 445.930 295.720 448.770 299.870 ;
        RECT 449.610 295.720 452.450 299.870 ;
        RECT 453.290 295.720 456.130 299.870 ;
        RECT 456.970 295.720 459.350 299.870 ;
        RECT 460.190 295.720 463.030 299.870 ;
        RECT 463.870 295.720 466.710 299.870 ;
        RECT 467.550 295.720 470.390 299.870 ;
        RECT 471.230 295.720 474.070 299.870 ;
        RECT 474.910 295.720 477.290 299.870 ;
        RECT 478.130 295.720 480.970 299.870 ;
        RECT 481.810 295.720 484.650 299.870 ;
        RECT 485.490 295.720 488.330 299.870 ;
        RECT 489.170 295.720 491.550 299.870 ;
        RECT 492.390 295.720 495.230 299.870 ;
        RECT 496.070 295.720 498.910 299.870 ;
        RECT 499.750 295.720 502.590 299.870 ;
        RECT 503.430 295.720 506.270 299.870 ;
        RECT 507.110 295.720 509.490 299.870 ;
        RECT 510.330 295.720 513.170 299.870 ;
        RECT 514.010 295.720 516.850 299.870 ;
        RECT 517.690 295.720 520.530 299.870 ;
        RECT 521.370 295.720 524.210 299.870 ;
        RECT 525.050 295.720 527.430 299.870 ;
        RECT 528.270 295.720 531.110 299.870 ;
        RECT 531.950 295.720 534.790 299.870 ;
        RECT 535.630 295.720 538.470 299.870 ;
        RECT 539.310 295.720 541.690 299.870 ;
        RECT 542.530 295.720 545.370 299.870 ;
        RECT 546.210 295.720 549.050 299.870 ;
        RECT 549.890 295.720 552.730 299.870 ;
        RECT 553.570 295.720 556.410 299.870 ;
        RECT 557.250 295.720 559.630 299.870 ;
        RECT 560.470 295.720 563.310 299.870 ;
        RECT 564.150 295.720 566.990 299.870 ;
        RECT 567.830 295.720 570.670 299.870 ;
        RECT 571.510 295.720 574.350 299.870 ;
        RECT 575.190 295.720 577.570 299.870 ;
        RECT 578.410 295.720 581.250 299.870 ;
        RECT 582.090 295.720 584.930 299.870 ;
        RECT 585.770 295.720 588.610 299.870 ;
        RECT 589.450 295.720 592.290 299.870 ;
        RECT 593.130 295.720 595.510 299.870 ;
        RECT 596.350 295.720 599.190 299.870 ;
        RECT 600.030 295.720 602.870 299.870 ;
        RECT 603.710 295.720 606.550 299.870 ;
        RECT 607.390 295.720 609.770 299.870 ;
        RECT 610.610 295.720 613.450 299.870 ;
        RECT 614.290 295.720 617.130 299.870 ;
        RECT 617.970 295.720 620.810 299.870 ;
        RECT 621.650 295.720 624.490 299.870 ;
        RECT 625.330 295.720 627.710 299.870 ;
        RECT 628.550 295.720 631.390 299.870 ;
        RECT 632.230 295.720 635.070 299.870 ;
        RECT 635.910 295.720 638.750 299.870 ;
        RECT 639.590 295.720 642.430 299.870 ;
        RECT 643.270 295.720 645.650 299.870 ;
        RECT 646.490 295.720 649.330 299.870 ;
        RECT 650.170 295.720 653.010 299.870 ;
        RECT 653.850 295.720 656.690 299.870 ;
        RECT 657.530 295.720 660.370 299.870 ;
        RECT 661.210 295.720 663.590 299.870 ;
        RECT 664.430 295.720 667.270 299.870 ;
        RECT 668.110 295.720 670.950 299.870 ;
        RECT 671.790 295.720 674.630 299.870 ;
        RECT 675.470 295.720 677.850 299.870 ;
        RECT 678.690 295.720 681.530 299.870 ;
        RECT 682.370 295.720 685.210 299.870 ;
        RECT 686.050 295.720 688.890 299.870 ;
        RECT 689.730 295.720 692.570 299.870 ;
        RECT 693.410 295.720 695.790 299.870 ;
        RECT 696.630 295.720 699.470 299.870 ;
        RECT 700.310 295.720 703.150 299.870 ;
        RECT 703.990 295.720 706.830 299.870 ;
        RECT 707.670 295.720 710.510 299.870 ;
        RECT 711.350 295.720 713.730 299.870 ;
        RECT 714.570 295.720 717.410 299.870 ;
        RECT 718.250 295.720 721.090 299.870 ;
        RECT 721.930 295.720 724.770 299.870 ;
        RECT 725.610 295.720 727.990 299.870 ;
        RECT 728.830 295.720 731.670 299.870 ;
        RECT 732.510 295.720 735.350 299.870 ;
        RECT 736.190 295.720 739.030 299.870 ;
        RECT 739.870 295.720 742.710 299.870 ;
        RECT 743.550 295.720 745.930 299.870 ;
        RECT 746.770 295.720 749.610 299.870 ;
        RECT 750.450 295.720 753.290 299.870 ;
        RECT 754.130 295.720 756.970 299.870 ;
        RECT 757.810 295.720 760.650 299.870 ;
        RECT 761.490 295.720 763.870 299.870 ;
        RECT 764.710 295.720 767.550 299.870 ;
        RECT 768.390 295.720 771.230 299.870 ;
        RECT 772.070 295.720 774.910 299.870 ;
        RECT 775.750 295.720 778.590 299.870 ;
        RECT 779.430 295.720 781.810 299.870 ;
        RECT 782.650 295.720 785.490 299.870 ;
        RECT 786.330 295.720 789.170 299.870 ;
        RECT 790.010 295.720 792.850 299.870 ;
        RECT 793.690 295.720 796.070 299.870 ;
        RECT 796.910 295.720 799.750 299.870 ;
        RECT 800.590 295.720 803.430 299.870 ;
        RECT 804.270 295.720 807.110 299.870 ;
        RECT 807.950 295.720 810.790 299.870 ;
        RECT 811.630 295.720 814.010 299.870 ;
        RECT 814.850 295.720 817.690 299.870 ;
        RECT 818.530 295.720 821.370 299.870 ;
        RECT 822.210 295.720 825.050 299.870 ;
        RECT 825.890 295.720 828.730 299.870 ;
        RECT 829.570 295.720 831.950 299.870 ;
        RECT 832.790 295.720 835.630 299.870 ;
        RECT 836.470 295.720 839.310 299.870 ;
        RECT 840.150 295.720 842.990 299.870 ;
        RECT 843.830 295.720 846.210 299.870 ;
        RECT 847.050 295.720 849.890 299.870 ;
        RECT 850.730 295.720 853.570 299.870 ;
        RECT 854.410 295.720 857.250 299.870 ;
        RECT 858.090 295.720 860.930 299.870 ;
        RECT 861.770 295.720 864.150 299.870 ;
        RECT 864.990 295.720 867.830 299.870 ;
        RECT 868.670 295.720 871.510 299.870 ;
        RECT 872.350 295.720 875.190 299.870 ;
        RECT 876.030 295.720 878.870 299.870 ;
        RECT 879.710 295.720 882.090 299.870 ;
        RECT 882.930 295.720 885.770 299.870 ;
        RECT 886.610 295.720 889.450 299.870 ;
        RECT 890.290 295.720 893.130 299.870 ;
        RECT 893.970 295.720 896.810 299.870 ;
        RECT 897.650 295.720 900.030 299.870 ;
        RECT 900.870 295.720 903.710 299.870 ;
        RECT 904.550 295.720 907.390 299.870 ;
        RECT 908.230 295.720 911.070 299.870 ;
        RECT 911.910 295.720 914.290 299.870 ;
        RECT 915.130 295.720 917.970 299.870 ;
        RECT 918.810 295.720 921.650 299.870 ;
        RECT 922.490 295.720 925.330 299.870 ;
        RECT 926.170 295.720 929.010 299.870 ;
        RECT 929.850 295.720 932.230 299.870 ;
        RECT 933.070 295.720 935.910 299.870 ;
        RECT 936.750 295.720 939.590 299.870 ;
        RECT 940.430 295.720 943.270 299.870 ;
        RECT 944.110 295.720 946.950 299.870 ;
        RECT 947.790 295.720 950.170 299.870 ;
        RECT 951.010 295.720 953.850 299.870 ;
        RECT 954.690 295.720 957.530 299.870 ;
        RECT 958.370 295.720 961.210 299.870 ;
        RECT 962.050 295.720 964.430 299.870 ;
        RECT 965.270 295.720 968.110 299.870 ;
        RECT 968.950 295.720 971.790 299.870 ;
        RECT 972.630 295.720 975.470 299.870 ;
        RECT 976.310 295.720 979.150 299.870 ;
        RECT 979.990 295.720 982.370 299.870 ;
        RECT 983.210 295.720 986.050 299.870 ;
        RECT 986.890 295.720 989.730 299.870 ;
        RECT 990.570 295.720 993.410 299.870 ;
        RECT 994.250 295.720 997.090 299.870 ;
        RECT 997.930 295.720 1000.310 299.870 ;
        RECT 1001.150 295.720 1003.990 299.870 ;
        RECT 1004.830 295.720 1007.670 299.870 ;
        RECT 1008.510 295.720 1011.350 299.870 ;
        RECT 1012.190 295.720 1015.030 299.870 ;
        RECT 1015.870 295.720 1018.250 299.870 ;
        RECT 1019.090 295.720 1021.930 299.870 ;
        RECT 1022.770 295.720 1025.610 299.870 ;
        RECT 1026.450 295.720 1029.290 299.870 ;
        RECT 1030.130 295.720 1032.510 299.870 ;
        RECT 1033.350 295.720 1036.190 299.870 ;
        RECT 1037.030 295.720 1039.870 299.870 ;
        RECT 1040.710 295.720 1043.550 299.870 ;
        RECT 1044.390 295.720 1047.230 299.870 ;
        RECT 1048.070 295.720 1050.450 299.870 ;
        RECT 1051.290 295.720 1054.130 299.870 ;
        RECT 1054.970 295.720 1057.810 299.870 ;
        RECT 1058.650 295.720 1061.490 299.870 ;
        RECT 1062.330 295.720 1065.170 299.870 ;
        RECT 1066.010 295.720 1068.390 299.870 ;
        RECT 1069.230 295.720 1072.070 299.870 ;
        RECT 1072.910 295.720 1075.750 299.870 ;
        RECT 1076.590 295.720 1079.430 299.870 ;
        RECT 1080.270 295.720 1082.650 299.870 ;
        RECT 1083.490 295.720 1086.330 299.870 ;
        RECT 1087.170 295.720 1090.010 299.870 ;
        RECT 1090.850 295.720 1093.690 299.870 ;
        RECT 1094.530 295.720 1097.370 299.870 ;
        RECT 1098.210 295.720 1100.590 299.870 ;
        RECT 1101.430 295.720 1104.270 299.870 ;
        RECT 1105.110 295.720 1107.950 299.870 ;
        RECT 1108.790 295.720 1111.630 299.870 ;
        RECT 1112.470 295.720 1115.310 299.870 ;
        RECT 1116.150 295.720 1118.530 299.870 ;
        RECT 1119.370 295.720 1122.210 299.870 ;
        RECT 1123.050 295.720 1125.890 299.870 ;
        RECT 1126.730 295.720 1129.570 299.870 ;
        RECT 1130.410 295.720 1133.250 299.870 ;
        RECT 1134.090 295.720 1136.470 299.870 ;
        RECT 1137.310 295.720 1140.150 299.870 ;
        RECT 1140.990 295.720 1143.830 299.870 ;
        RECT 1144.670 295.720 1147.510 299.870 ;
        RECT 1148.350 295.720 1150.730 299.870 ;
        RECT 1151.570 295.720 1154.410 299.870 ;
        RECT 1155.250 295.720 1158.090 299.870 ;
        RECT 1158.930 295.720 1161.770 299.870 ;
        RECT 1162.610 295.720 1165.450 299.870 ;
        RECT 1166.290 295.720 1168.670 299.870 ;
        RECT 1169.510 295.720 1172.350 299.870 ;
        RECT 1173.190 295.720 1176.030 299.870 ;
        RECT 1176.870 295.720 1179.710 299.870 ;
        RECT 1180.550 295.720 1183.390 299.870 ;
        RECT 1184.230 295.720 1186.610 299.870 ;
        RECT 1187.450 295.720 1190.290 299.870 ;
        RECT 1191.130 295.720 1193.970 299.870 ;
        RECT 1194.810 295.720 1197.650 299.870 ;
        RECT 1198.490 295.720 1199.120 299.870 ;
        RECT 1.020 4.280 1199.120 295.720 ;
        RECT 1.570 0.690 2.570 4.280 ;
        RECT 3.410 0.690 4.870 4.280 ;
        RECT 5.710 0.690 7.170 4.280 ;
        RECT 8.010 0.690 9.470 4.280 ;
        RECT 10.310 0.690 11.310 4.280 ;
        RECT 12.150 0.690 13.610 4.280 ;
        RECT 14.450 0.690 15.910 4.280 ;
        RECT 16.750 0.690 18.210 4.280 ;
        RECT 19.050 0.690 20.510 4.280 ;
        RECT 21.350 0.690 22.350 4.280 ;
        RECT 23.190 0.690 24.650 4.280 ;
        RECT 25.490 0.690 26.950 4.280 ;
        RECT 27.790 0.690 29.250 4.280 ;
        RECT 30.090 0.690 31.550 4.280 ;
        RECT 32.390 0.690 33.390 4.280 ;
        RECT 34.230 0.690 35.690 4.280 ;
        RECT 36.530 0.690 37.990 4.280 ;
        RECT 38.830 0.690 40.290 4.280 ;
        RECT 41.130 0.690 42.130 4.280 ;
        RECT 42.970 0.690 44.430 4.280 ;
        RECT 45.270 0.690 46.730 4.280 ;
        RECT 47.570 0.690 49.030 4.280 ;
        RECT 49.870 0.690 51.330 4.280 ;
        RECT 52.170 0.690 53.170 4.280 ;
        RECT 54.010 0.690 55.470 4.280 ;
        RECT 56.310 0.690 57.770 4.280 ;
        RECT 58.610 0.690 60.070 4.280 ;
        RECT 60.910 0.690 62.370 4.280 ;
        RECT 63.210 0.690 64.210 4.280 ;
        RECT 65.050 0.690 66.510 4.280 ;
        RECT 67.350 0.690 68.810 4.280 ;
        RECT 69.650 0.690 71.110 4.280 ;
        RECT 71.950 0.690 72.950 4.280 ;
        RECT 73.790 0.690 75.250 4.280 ;
        RECT 76.090 0.690 77.550 4.280 ;
        RECT 78.390 0.690 79.850 4.280 ;
        RECT 80.690 0.690 82.150 4.280 ;
        RECT 82.990 0.690 83.990 4.280 ;
        RECT 84.830 0.690 86.290 4.280 ;
        RECT 87.130 0.690 88.590 4.280 ;
        RECT 89.430 0.690 90.890 4.280 ;
        RECT 91.730 0.690 93.190 4.280 ;
        RECT 94.030 0.690 95.030 4.280 ;
        RECT 95.870 0.690 97.330 4.280 ;
        RECT 98.170 0.690 99.630 4.280 ;
        RECT 100.470 0.690 101.930 4.280 ;
        RECT 102.770 0.690 103.770 4.280 ;
        RECT 104.610 0.690 106.070 4.280 ;
        RECT 106.910 0.690 108.370 4.280 ;
        RECT 109.210 0.690 110.670 4.280 ;
        RECT 111.510 0.690 112.970 4.280 ;
        RECT 113.810 0.690 114.810 4.280 ;
        RECT 115.650 0.690 117.110 4.280 ;
        RECT 117.950 0.690 119.410 4.280 ;
        RECT 120.250 0.690 121.710 4.280 ;
        RECT 122.550 0.690 124.010 4.280 ;
        RECT 124.850 0.690 125.850 4.280 ;
        RECT 126.690 0.690 128.150 4.280 ;
        RECT 128.990 0.690 130.450 4.280 ;
        RECT 131.290 0.690 132.750 4.280 ;
        RECT 133.590 0.690 135.050 4.280 ;
        RECT 135.890 0.690 136.890 4.280 ;
        RECT 137.730 0.690 139.190 4.280 ;
        RECT 140.030 0.690 141.490 4.280 ;
        RECT 142.330 0.690 143.790 4.280 ;
        RECT 144.630 0.690 145.630 4.280 ;
        RECT 146.470 0.690 147.930 4.280 ;
        RECT 148.770 0.690 150.230 4.280 ;
        RECT 151.070 0.690 152.530 4.280 ;
        RECT 153.370 0.690 154.830 4.280 ;
        RECT 155.670 0.690 156.670 4.280 ;
        RECT 157.510 0.690 158.970 4.280 ;
        RECT 159.810 0.690 161.270 4.280 ;
        RECT 162.110 0.690 163.570 4.280 ;
        RECT 164.410 0.690 165.870 4.280 ;
        RECT 166.710 0.690 167.710 4.280 ;
        RECT 168.550 0.690 170.010 4.280 ;
        RECT 170.850 0.690 172.310 4.280 ;
        RECT 173.150 0.690 174.610 4.280 ;
        RECT 175.450 0.690 176.450 4.280 ;
        RECT 177.290 0.690 178.750 4.280 ;
        RECT 179.590 0.690 181.050 4.280 ;
        RECT 181.890 0.690 183.350 4.280 ;
        RECT 184.190 0.690 185.650 4.280 ;
        RECT 186.490 0.690 187.490 4.280 ;
        RECT 188.330 0.690 189.790 4.280 ;
        RECT 190.630 0.690 192.090 4.280 ;
        RECT 192.930 0.690 194.390 4.280 ;
        RECT 195.230 0.690 196.690 4.280 ;
        RECT 197.530 0.690 198.530 4.280 ;
        RECT 199.370 0.690 200.830 4.280 ;
        RECT 201.670 0.690 203.130 4.280 ;
        RECT 203.970 0.690 205.430 4.280 ;
        RECT 206.270 0.690 207.270 4.280 ;
        RECT 208.110 0.690 209.570 4.280 ;
        RECT 210.410 0.690 211.870 4.280 ;
        RECT 212.710 0.690 214.170 4.280 ;
        RECT 215.010 0.690 216.470 4.280 ;
        RECT 217.310 0.690 218.310 4.280 ;
        RECT 219.150 0.690 220.610 4.280 ;
        RECT 221.450 0.690 222.910 4.280 ;
        RECT 223.750 0.690 225.210 4.280 ;
        RECT 226.050 0.690 227.510 4.280 ;
        RECT 228.350 0.690 229.350 4.280 ;
        RECT 230.190 0.690 231.650 4.280 ;
        RECT 232.490 0.690 233.950 4.280 ;
        RECT 234.790 0.690 236.250 4.280 ;
        RECT 237.090 0.690 238.550 4.280 ;
        RECT 239.390 0.690 240.390 4.280 ;
        RECT 241.230 0.690 242.690 4.280 ;
        RECT 243.530 0.690 244.990 4.280 ;
        RECT 245.830 0.690 247.290 4.280 ;
        RECT 248.130 0.690 249.130 4.280 ;
        RECT 249.970 0.690 251.430 4.280 ;
        RECT 252.270 0.690 253.730 4.280 ;
        RECT 254.570 0.690 256.030 4.280 ;
        RECT 256.870 0.690 258.330 4.280 ;
        RECT 259.170 0.690 260.170 4.280 ;
        RECT 261.010 0.690 262.470 4.280 ;
        RECT 263.310 0.690 264.770 4.280 ;
        RECT 265.610 0.690 267.070 4.280 ;
        RECT 267.910 0.690 269.370 4.280 ;
        RECT 270.210 0.690 271.210 4.280 ;
        RECT 272.050 0.690 273.510 4.280 ;
        RECT 274.350 0.690 275.810 4.280 ;
        RECT 276.650 0.690 278.110 4.280 ;
        RECT 278.950 0.690 279.950 4.280 ;
        RECT 280.790 0.690 282.250 4.280 ;
        RECT 283.090 0.690 284.550 4.280 ;
        RECT 285.390 0.690 286.850 4.280 ;
        RECT 287.690 0.690 289.150 4.280 ;
        RECT 289.990 0.690 290.990 4.280 ;
        RECT 291.830 0.690 293.290 4.280 ;
        RECT 294.130 0.690 295.590 4.280 ;
        RECT 296.430 0.690 297.890 4.280 ;
        RECT 298.730 0.690 300.190 4.280 ;
        RECT 301.030 0.690 302.030 4.280 ;
        RECT 302.870 0.690 304.330 4.280 ;
        RECT 305.170 0.690 306.630 4.280 ;
        RECT 307.470 0.690 308.930 4.280 ;
        RECT 309.770 0.690 310.770 4.280 ;
        RECT 311.610 0.690 313.070 4.280 ;
        RECT 313.910 0.690 315.370 4.280 ;
        RECT 316.210 0.690 317.670 4.280 ;
        RECT 318.510 0.690 319.970 4.280 ;
        RECT 320.810 0.690 321.810 4.280 ;
        RECT 322.650 0.690 324.110 4.280 ;
        RECT 324.950 0.690 326.410 4.280 ;
        RECT 327.250 0.690 328.710 4.280 ;
        RECT 329.550 0.690 331.010 4.280 ;
        RECT 331.850 0.690 332.850 4.280 ;
        RECT 333.690 0.690 335.150 4.280 ;
        RECT 335.990 0.690 337.450 4.280 ;
        RECT 338.290 0.690 339.750 4.280 ;
        RECT 340.590 0.690 342.050 4.280 ;
        RECT 342.890 0.690 343.890 4.280 ;
        RECT 344.730 0.690 346.190 4.280 ;
        RECT 347.030 0.690 348.490 4.280 ;
        RECT 349.330 0.690 350.790 4.280 ;
        RECT 351.630 0.690 352.630 4.280 ;
        RECT 353.470 0.690 354.930 4.280 ;
        RECT 355.770 0.690 357.230 4.280 ;
        RECT 358.070 0.690 359.530 4.280 ;
        RECT 360.370 0.690 361.830 4.280 ;
        RECT 362.670 0.690 363.670 4.280 ;
        RECT 364.510 0.690 365.970 4.280 ;
        RECT 366.810 0.690 368.270 4.280 ;
        RECT 369.110 0.690 370.570 4.280 ;
        RECT 371.410 0.690 372.870 4.280 ;
        RECT 373.710 0.690 374.710 4.280 ;
        RECT 375.550 0.690 377.010 4.280 ;
        RECT 377.850 0.690 379.310 4.280 ;
        RECT 380.150 0.690 381.610 4.280 ;
        RECT 382.450 0.690 383.450 4.280 ;
        RECT 384.290 0.690 385.750 4.280 ;
        RECT 386.590 0.690 388.050 4.280 ;
        RECT 388.890 0.690 390.350 4.280 ;
        RECT 391.190 0.690 392.650 4.280 ;
        RECT 393.490 0.690 394.490 4.280 ;
        RECT 395.330 0.690 396.790 4.280 ;
        RECT 397.630 0.690 399.090 4.280 ;
        RECT 399.930 0.690 401.390 4.280 ;
        RECT 402.230 0.690 403.690 4.280 ;
        RECT 404.530 0.690 405.530 4.280 ;
        RECT 406.370 0.690 407.830 4.280 ;
        RECT 408.670 0.690 410.130 4.280 ;
        RECT 410.970 0.690 412.430 4.280 ;
        RECT 413.270 0.690 414.270 4.280 ;
        RECT 415.110 0.690 416.570 4.280 ;
        RECT 417.410 0.690 418.870 4.280 ;
        RECT 419.710 0.690 421.170 4.280 ;
        RECT 422.010 0.690 423.470 4.280 ;
        RECT 424.310 0.690 425.310 4.280 ;
        RECT 426.150 0.690 427.610 4.280 ;
        RECT 428.450 0.690 429.910 4.280 ;
        RECT 430.750 0.690 432.210 4.280 ;
        RECT 433.050 0.690 434.510 4.280 ;
        RECT 435.350 0.690 436.350 4.280 ;
        RECT 437.190 0.690 438.650 4.280 ;
        RECT 439.490 0.690 440.950 4.280 ;
        RECT 441.790 0.690 443.250 4.280 ;
        RECT 444.090 0.690 445.550 4.280 ;
        RECT 446.390 0.690 447.390 4.280 ;
        RECT 448.230 0.690 449.690 4.280 ;
        RECT 450.530 0.690 451.990 4.280 ;
        RECT 452.830 0.690 454.290 4.280 ;
        RECT 455.130 0.690 456.130 4.280 ;
        RECT 456.970 0.690 458.430 4.280 ;
        RECT 459.270 0.690 460.730 4.280 ;
        RECT 461.570 0.690 463.030 4.280 ;
        RECT 463.870 0.690 465.330 4.280 ;
        RECT 466.170 0.690 467.170 4.280 ;
        RECT 468.010 0.690 469.470 4.280 ;
        RECT 470.310 0.690 471.770 4.280 ;
        RECT 472.610 0.690 474.070 4.280 ;
        RECT 474.910 0.690 476.370 4.280 ;
        RECT 477.210 0.690 478.210 4.280 ;
        RECT 479.050 0.690 480.510 4.280 ;
        RECT 481.350 0.690 482.810 4.280 ;
        RECT 483.650 0.690 485.110 4.280 ;
        RECT 485.950 0.690 486.950 4.280 ;
        RECT 487.790 0.690 489.250 4.280 ;
        RECT 490.090 0.690 491.550 4.280 ;
        RECT 492.390 0.690 493.850 4.280 ;
        RECT 494.690 0.690 496.150 4.280 ;
        RECT 496.990 0.690 497.990 4.280 ;
        RECT 498.830 0.690 500.290 4.280 ;
        RECT 501.130 0.690 502.590 4.280 ;
        RECT 503.430 0.690 504.890 4.280 ;
        RECT 505.730 0.690 507.190 4.280 ;
        RECT 508.030 0.690 509.030 4.280 ;
        RECT 509.870 0.690 511.330 4.280 ;
        RECT 512.170 0.690 513.630 4.280 ;
        RECT 514.470 0.690 515.930 4.280 ;
        RECT 516.770 0.690 517.770 4.280 ;
        RECT 518.610 0.690 520.070 4.280 ;
        RECT 520.910 0.690 522.370 4.280 ;
        RECT 523.210 0.690 524.670 4.280 ;
        RECT 525.510 0.690 526.970 4.280 ;
        RECT 527.810 0.690 528.810 4.280 ;
        RECT 529.650 0.690 531.110 4.280 ;
        RECT 531.950 0.690 533.410 4.280 ;
        RECT 534.250 0.690 535.710 4.280 ;
        RECT 536.550 0.690 538.010 4.280 ;
        RECT 538.850 0.690 539.850 4.280 ;
        RECT 540.690 0.690 542.150 4.280 ;
        RECT 542.990 0.690 544.450 4.280 ;
        RECT 545.290 0.690 546.750 4.280 ;
        RECT 547.590 0.690 549.050 4.280 ;
        RECT 549.890 0.690 550.890 4.280 ;
        RECT 551.730 0.690 553.190 4.280 ;
        RECT 554.030 0.690 555.490 4.280 ;
        RECT 556.330 0.690 557.790 4.280 ;
        RECT 558.630 0.690 559.630 4.280 ;
        RECT 560.470 0.690 561.930 4.280 ;
        RECT 562.770 0.690 564.230 4.280 ;
        RECT 565.070 0.690 566.530 4.280 ;
        RECT 567.370 0.690 568.830 4.280 ;
        RECT 569.670 0.690 570.670 4.280 ;
        RECT 571.510 0.690 572.970 4.280 ;
        RECT 573.810 0.690 575.270 4.280 ;
        RECT 576.110 0.690 577.570 4.280 ;
        RECT 578.410 0.690 579.870 4.280 ;
        RECT 580.710 0.690 581.710 4.280 ;
        RECT 582.550 0.690 584.010 4.280 ;
        RECT 584.850 0.690 586.310 4.280 ;
        RECT 587.150 0.690 588.610 4.280 ;
        RECT 589.450 0.690 590.450 4.280 ;
        RECT 591.290 0.690 592.750 4.280 ;
        RECT 593.590 0.690 595.050 4.280 ;
        RECT 595.890 0.690 597.350 4.280 ;
        RECT 598.190 0.690 599.650 4.280 ;
        RECT 600.490 0.690 601.490 4.280 ;
        RECT 602.330 0.690 603.790 4.280 ;
        RECT 604.630 0.690 606.090 4.280 ;
        RECT 606.930 0.690 608.390 4.280 ;
        RECT 609.230 0.690 610.690 4.280 ;
        RECT 611.530 0.690 612.530 4.280 ;
        RECT 613.370 0.690 614.830 4.280 ;
        RECT 615.670 0.690 617.130 4.280 ;
        RECT 617.970 0.690 619.430 4.280 ;
        RECT 620.270 0.690 621.270 4.280 ;
        RECT 622.110 0.690 623.570 4.280 ;
        RECT 624.410 0.690 625.870 4.280 ;
        RECT 626.710 0.690 628.170 4.280 ;
        RECT 629.010 0.690 630.470 4.280 ;
        RECT 631.310 0.690 632.310 4.280 ;
        RECT 633.150 0.690 634.610 4.280 ;
        RECT 635.450 0.690 636.910 4.280 ;
        RECT 637.750 0.690 639.210 4.280 ;
        RECT 640.050 0.690 641.510 4.280 ;
        RECT 642.350 0.690 643.350 4.280 ;
        RECT 644.190 0.690 645.650 4.280 ;
        RECT 646.490 0.690 647.950 4.280 ;
        RECT 648.790 0.690 650.250 4.280 ;
        RECT 651.090 0.690 652.090 4.280 ;
        RECT 652.930 0.690 654.390 4.280 ;
        RECT 655.230 0.690 656.690 4.280 ;
        RECT 657.530 0.690 658.990 4.280 ;
        RECT 659.830 0.690 661.290 4.280 ;
        RECT 662.130 0.690 663.130 4.280 ;
        RECT 663.970 0.690 665.430 4.280 ;
        RECT 666.270 0.690 667.730 4.280 ;
        RECT 668.570 0.690 670.030 4.280 ;
        RECT 670.870 0.690 672.330 4.280 ;
        RECT 673.170 0.690 674.170 4.280 ;
        RECT 675.010 0.690 676.470 4.280 ;
        RECT 677.310 0.690 678.770 4.280 ;
        RECT 679.610 0.690 681.070 4.280 ;
        RECT 681.910 0.690 683.370 4.280 ;
        RECT 684.210 0.690 685.210 4.280 ;
        RECT 686.050 0.690 687.510 4.280 ;
        RECT 688.350 0.690 689.810 4.280 ;
        RECT 690.650 0.690 692.110 4.280 ;
        RECT 692.950 0.690 693.950 4.280 ;
        RECT 694.790 0.690 696.250 4.280 ;
        RECT 697.090 0.690 698.550 4.280 ;
        RECT 699.390 0.690 700.850 4.280 ;
        RECT 701.690 0.690 703.150 4.280 ;
        RECT 703.990 0.690 704.990 4.280 ;
        RECT 705.830 0.690 707.290 4.280 ;
        RECT 708.130 0.690 709.590 4.280 ;
        RECT 710.430 0.690 711.890 4.280 ;
        RECT 712.730 0.690 714.190 4.280 ;
        RECT 715.030 0.690 716.030 4.280 ;
        RECT 716.870 0.690 718.330 4.280 ;
        RECT 719.170 0.690 720.630 4.280 ;
        RECT 721.470 0.690 722.930 4.280 ;
        RECT 723.770 0.690 724.770 4.280 ;
        RECT 725.610 0.690 727.070 4.280 ;
        RECT 727.910 0.690 729.370 4.280 ;
        RECT 730.210 0.690 731.670 4.280 ;
        RECT 732.510 0.690 733.970 4.280 ;
        RECT 734.810 0.690 735.810 4.280 ;
        RECT 736.650 0.690 738.110 4.280 ;
        RECT 738.950 0.690 740.410 4.280 ;
        RECT 741.250 0.690 742.710 4.280 ;
        RECT 743.550 0.690 745.010 4.280 ;
        RECT 745.850 0.690 746.850 4.280 ;
        RECT 747.690 0.690 749.150 4.280 ;
        RECT 749.990 0.690 751.450 4.280 ;
        RECT 752.290 0.690 753.750 4.280 ;
        RECT 754.590 0.690 755.590 4.280 ;
        RECT 756.430 0.690 757.890 4.280 ;
        RECT 758.730 0.690 760.190 4.280 ;
        RECT 761.030 0.690 762.490 4.280 ;
        RECT 763.330 0.690 764.790 4.280 ;
        RECT 765.630 0.690 766.630 4.280 ;
        RECT 767.470 0.690 768.930 4.280 ;
        RECT 769.770 0.690 771.230 4.280 ;
        RECT 772.070 0.690 773.530 4.280 ;
        RECT 774.370 0.690 775.830 4.280 ;
        RECT 776.670 0.690 777.670 4.280 ;
        RECT 778.510 0.690 779.970 4.280 ;
        RECT 780.810 0.690 782.270 4.280 ;
        RECT 783.110 0.690 784.570 4.280 ;
        RECT 785.410 0.690 786.870 4.280 ;
        RECT 787.710 0.690 788.710 4.280 ;
        RECT 789.550 0.690 791.010 4.280 ;
        RECT 791.850 0.690 793.310 4.280 ;
        RECT 794.150 0.690 795.610 4.280 ;
        RECT 796.450 0.690 797.450 4.280 ;
        RECT 798.290 0.690 799.750 4.280 ;
        RECT 800.590 0.690 802.050 4.280 ;
        RECT 802.890 0.690 804.350 4.280 ;
        RECT 805.190 0.690 806.650 4.280 ;
        RECT 807.490 0.690 808.490 4.280 ;
        RECT 809.330 0.690 810.790 4.280 ;
        RECT 811.630 0.690 813.090 4.280 ;
        RECT 813.930 0.690 815.390 4.280 ;
        RECT 816.230 0.690 817.690 4.280 ;
        RECT 818.530 0.690 819.530 4.280 ;
        RECT 820.370 0.690 821.830 4.280 ;
        RECT 822.670 0.690 824.130 4.280 ;
        RECT 824.970 0.690 826.430 4.280 ;
        RECT 827.270 0.690 828.270 4.280 ;
        RECT 829.110 0.690 830.570 4.280 ;
        RECT 831.410 0.690 832.870 4.280 ;
        RECT 833.710 0.690 835.170 4.280 ;
        RECT 836.010 0.690 837.470 4.280 ;
        RECT 838.310 0.690 839.310 4.280 ;
        RECT 840.150 0.690 841.610 4.280 ;
        RECT 842.450 0.690 843.910 4.280 ;
        RECT 844.750 0.690 846.210 4.280 ;
        RECT 847.050 0.690 848.510 4.280 ;
        RECT 849.350 0.690 850.350 4.280 ;
        RECT 851.190 0.690 852.650 4.280 ;
        RECT 853.490 0.690 854.950 4.280 ;
        RECT 855.790 0.690 857.250 4.280 ;
        RECT 858.090 0.690 859.090 4.280 ;
        RECT 859.930 0.690 861.390 4.280 ;
        RECT 862.230 0.690 863.690 4.280 ;
        RECT 864.530 0.690 865.990 4.280 ;
        RECT 866.830 0.690 868.290 4.280 ;
        RECT 869.130 0.690 870.130 4.280 ;
        RECT 870.970 0.690 872.430 4.280 ;
        RECT 873.270 0.690 874.730 4.280 ;
        RECT 875.570 0.690 877.030 4.280 ;
        RECT 877.870 0.690 879.330 4.280 ;
        RECT 880.170 0.690 881.170 4.280 ;
        RECT 882.010 0.690 883.470 4.280 ;
        RECT 884.310 0.690 885.770 4.280 ;
        RECT 886.610 0.690 888.070 4.280 ;
        RECT 888.910 0.690 890.370 4.280 ;
        RECT 891.210 0.690 892.210 4.280 ;
        RECT 893.050 0.690 894.510 4.280 ;
        RECT 895.350 0.690 896.810 4.280 ;
        RECT 897.650 0.690 899.110 4.280 ;
        RECT 899.950 0.690 900.950 4.280 ;
        RECT 901.790 0.690 903.250 4.280 ;
        RECT 904.090 0.690 905.550 4.280 ;
        RECT 906.390 0.690 907.850 4.280 ;
        RECT 908.690 0.690 910.150 4.280 ;
        RECT 910.990 0.690 911.990 4.280 ;
        RECT 912.830 0.690 914.290 4.280 ;
        RECT 915.130 0.690 916.590 4.280 ;
        RECT 917.430 0.690 918.890 4.280 ;
        RECT 919.730 0.690 921.190 4.280 ;
        RECT 922.030 0.690 923.030 4.280 ;
        RECT 923.870 0.690 925.330 4.280 ;
        RECT 926.170 0.690 927.630 4.280 ;
        RECT 928.470 0.690 929.930 4.280 ;
        RECT 930.770 0.690 931.770 4.280 ;
        RECT 932.610 0.690 934.070 4.280 ;
        RECT 934.910 0.690 936.370 4.280 ;
        RECT 937.210 0.690 938.670 4.280 ;
        RECT 939.510 0.690 940.970 4.280 ;
        RECT 941.810 0.690 942.810 4.280 ;
        RECT 943.650 0.690 945.110 4.280 ;
        RECT 945.950 0.690 947.410 4.280 ;
        RECT 948.250 0.690 949.710 4.280 ;
        RECT 950.550 0.690 952.010 4.280 ;
        RECT 952.850 0.690 953.850 4.280 ;
        RECT 954.690 0.690 956.150 4.280 ;
        RECT 956.990 0.690 958.450 4.280 ;
        RECT 959.290 0.690 960.750 4.280 ;
        RECT 961.590 0.690 962.590 4.280 ;
        RECT 963.430 0.690 964.890 4.280 ;
        RECT 965.730 0.690 967.190 4.280 ;
        RECT 968.030 0.690 969.490 4.280 ;
        RECT 970.330 0.690 971.790 4.280 ;
        RECT 972.630 0.690 973.630 4.280 ;
        RECT 974.470 0.690 975.930 4.280 ;
        RECT 976.770 0.690 978.230 4.280 ;
        RECT 979.070 0.690 980.530 4.280 ;
        RECT 981.370 0.690 982.830 4.280 ;
        RECT 983.670 0.690 984.670 4.280 ;
        RECT 985.510 0.690 986.970 4.280 ;
        RECT 987.810 0.690 989.270 4.280 ;
        RECT 990.110 0.690 991.570 4.280 ;
        RECT 992.410 0.690 993.870 4.280 ;
        RECT 994.710 0.690 995.710 4.280 ;
        RECT 996.550 0.690 998.010 4.280 ;
        RECT 998.850 0.690 1000.310 4.280 ;
        RECT 1001.150 0.690 1002.610 4.280 ;
        RECT 1003.450 0.690 1004.450 4.280 ;
        RECT 1005.290 0.690 1006.750 4.280 ;
        RECT 1007.590 0.690 1009.050 4.280 ;
        RECT 1009.890 0.690 1011.350 4.280 ;
        RECT 1012.190 0.690 1013.650 4.280 ;
        RECT 1014.490 0.690 1015.490 4.280 ;
        RECT 1016.330 0.690 1017.790 4.280 ;
        RECT 1018.630 0.690 1020.090 4.280 ;
        RECT 1020.930 0.690 1022.390 4.280 ;
        RECT 1023.230 0.690 1024.690 4.280 ;
        RECT 1025.530 0.690 1026.530 4.280 ;
        RECT 1027.370 0.690 1028.830 4.280 ;
        RECT 1029.670 0.690 1031.130 4.280 ;
        RECT 1031.970 0.690 1033.430 4.280 ;
        RECT 1034.270 0.690 1035.270 4.280 ;
        RECT 1036.110 0.690 1037.570 4.280 ;
        RECT 1038.410 0.690 1039.870 4.280 ;
        RECT 1040.710 0.690 1042.170 4.280 ;
        RECT 1043.010 0.690 1044.470 4.280 ;
        RECT 1045.310 0.690 1046.310 4.280 ;
        RECT 1047.150 0.690 1048.610 4.280 ;
        RECT 1049.450 0.690 1050.910 4.280 ;
        RECT 1051.750 0.690 1053.210 4.280 ;
        RECT 1054.050 0.690 1055.510 4.280 ;
        RECT 1056.350 0.690 1057.350 4.280 ;
        RECT 1058.190 0.690 1059.650 4.280 ;
        RECT 1060.490 0.690 1061.950 4.280 ;
        RECT 1062.790 0.690 1064.250 4.280 ;
        RECT 1065.090 0.690 1066.090 4.280 ;
        RECT 1066.930 0.690 1068.390 4.280 ;
        RECT 1069.230 0.690 1070.690 4.280 ;
        RECT 1071.530 0.690 1072.990 4.280 ;
        RECT 1073.830 0.690 1075.290 4.280 ;
        RECT 1076.130 0.690 1077.130 4.280 ;
        RECT 1077.970 0.690 1079.430 4.280 ;
        RECT 1080.270 0.690 1081.730 4.280 ;
        RECT 1082.570 0.690 1084.030 4.280 ;
        RECT 1084.870 0.690 1086.330 4.280 ;
        RECT 1087.170 0.690 1088.170 4.280 ;
        RECT 1089.010 0.690 1090.470 4.280 ;
        RECT 1091.310 0.690 1092.770 4.280 ;
        RECT 1093.610 0.690 1095.070 4.280 ;
        RECT 1095.910 0.690 1097.370 4.280 ;
        RECT 1098.210 0.690 1099.210 4.280 ;
        RECT 1100.050 0.690 1101.510 4.280 ;
        RECT 1102.350 0.690 1103.810 4.280 ;
        RECT 1104.650 0.690 1106.110 4.280 ;
        RECT 1106.950 0.690 1107.950 4.280 ;
        RECT 1108.790 0.690 1110.250 4.280 ;
        RECT 1111.090 0.690 1112.550 4.280 ;
        RECT 1113.390 0.690 1114.850 4.280 ;
        RECT 1115.690 0.690 1117.150 4.280 ;
        RECT 1117.990 0.690 1118.990 4.280 ;
        RECT 1119.830 0.690 1121.290 4.280 ;
        RECT 1122.130 0.690 1123.590 4.280 ;
        RECT 1124.430 0.690 1125.890 4.280 ;
        RECT 1126.730 0.690 1128.190 4.280 ;
        RECT 1129.030 0.690 1130.030 4.280 ;
        RECT 1130.870 0.690 1132.330 4.280 ;
        RECT 1133.170 0.690 1134.630 4.280 ;
        RECT 1135.470 0.690 1136.930 4.280 ;
        RECT 1137.770 0.690 1138.770 4.280 ;
        RECT 1139.610 0.690 1141.070 4.280 ;
        RECT 1141.910 0.690 1143.370 4.280 ;
        RECT 1144.210 0.690 1145.670 4.280 ;
        RECT 1146.510 0.690 1147.970 4.280 ;
        RECT 1148.810 0.690 1149.810 4.280 ;
        RECT 1150.650 0.690 1152.110 4.280 ;
        RECT 1152.950 0.690 1154.410 4.280 ;
        RECT 1155.250 0.690 1156.710 4.280 ;
        RECT 1157.550 0.690 1159.010 4.280 ;
        RECT 1159.850 0.690 1160.850 4.280 ;
        RECT 1161.690 0.690 1163.150 4.280 ;
        RECT 1163.990 0.690 1165.450 4.280 ;
        RECT 1166.290 0.690 1167.750 4.280 ;
        RECT 1168.590 0.690 1169.590 4.280 ;
        RECT 1170.430 0.690 1171.890 4.280 ;
        RECT 1172.730 0.690 1174.190 4.280 ;
        RECT 1175.030 0.690 1176.490 4.280 ;
        RECT 1177.330 0.690 1178.790 4.280 ;
        RECT 1179.630 0.690 1180.630 4.280 ;
        RECT 1181.470 0.690 1182.930 4.280 ;
        RECT 1183.770 0.690 1185.230 4.280 ;
        RECT 1186.070 0.690 1187.530 4.280 ;
        RECT 1188.370 0.690 1189.830 4.280 ;
        RECT 1190.670 0.690 1191.670 4.280 ;
        RECT 1192.510 0.690 1193.970 4.280 ;
        RECT 1194.810 0.690 1196.270 4.280 ;
        RECT 1197.110 0.690 1198.570 4.280 ;
      LAYER met3 ;
        RECT 4.000 262.840 1196.000 296.300 ;
        RECT 4.000 261.440 1195.600 262.840 ;
        RECT 4.000 188.040 1196.000 261.440 ;
        RECT 4.000 186.640 1195.600 188.040 ;
        RECT 4.000 150.640 1196.000 186.640 ;
        RECT 4.400 149.240 1196.000 150.640 ;
        RECT 4.000 113.240 1196.000 149.240 ;
        RECT 4.000 111.840 1195.600 113.240 ;
        RECT 4.000 38.440 1196.000 111.840 ;
        RECT 4.000 37.040 1195.600 38.440 ;
        RECT 4.000 0.855 1196.000 37.040 ;
      LAYER met4 ;
        RECT 96.895 288.960 1112.905 296.305 ;
        RECT 96.895 10.240 97.440 288.960 ;
        RECT 99.840 10.240 174.240 288.960 ;
        RECT 176.640 10.240 251.040 288.960 ;
        RECT 253.440 10.240 327.840 288.960 ;
        RECT 330.240 10.240 404.640 288.960 ;
        RECT 407.040 10.240 481.440 288.960 ;
        RECT 483.840 10.240 558.240 288.960 ;
        RECT 560.640 10.240 635.040 288.960 ;
        RECT 637.440 10.240 711.840 288.960 ;
        RECT 714.240 10.240 788.640 288.960 ;
        RECT 791.040 10.240 865.440 288.960 ;
        RECT 867.840 10.240 942.240 288.960 ;
        RECT 944.640 10.240 1019.040 288.960 ;
        RECT 1021.440 10.240 1095.840 288.960 ;
        RECT 1098.240 10.240 1112.905 288.960 ;
        RECT 96.895 1.535 1112.905 10.240 ;
  END
END main_controller
END LIBRARY

