VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.330 2934.450 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 154.330 2934.450 157.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 294.330 2934.450 297.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 434.330 2934.450 437.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 574.330 2934.450 577.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 714.330 2934.450 717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 288.970 779.630 2532.070 782.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 854.330 2934.450 857.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 994.330 2934.450 997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1134.330 2934.450 1137.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1274.330 2934.450 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1414.330 2934.450 1417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1554.330 2934.450 1557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1694.330 2934.450 1697.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1828.970 1759.630 2112.070 1762.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1834.330 2934.450 1837.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1974.330 2934.450 1977.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2114.330 2934.450 2117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 288.970 2189.030 852.070 2192.130 ;
    END
    PORT
      LAYER met5 ;
        RECT 988.970 2189.030 1552.070 2192.130 ;
    END
    PORT
      LAYER met5 ;
        RECT 1968.970 2189.030 2532.070 2192.130 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2254.330 2934.450 2257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2394.330 2934.450 2397.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2534.330 2934.450 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2674.330 2934.450 2677.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 288.970 2739.630 2532.070 2742.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2814.330 2934.450 2817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2954.330 2934.450 2957.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3094.330 2934.450 3097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3234.330 2934.450 3237.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3374.330 2934.450 3377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 -9.470 292.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.970 -9.470 432.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 -9.470 572.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 -9.470 712.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.970 -9.470 852.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 988.970 -9.470 992.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.970 -9.470 1132.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -9.470 1272.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 -9.470 1412.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.970 -9.470 1552.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 -9.470 1692.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 -9.470 1972.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 -9.470 2112.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.970 -9.470 2252.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2388.970 -9.470 2392.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -9.470 2532.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 726.540 292.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.970 726.540 432.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 726.540 572.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 726.540 712.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.970 726.540 852.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 988.970 726.540 992.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.970 726.540 1132.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 726.540 1272.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 726.540 1412.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.970 726.540 1552.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 726.540 1692.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 726.540 1972.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 726.540 2112.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.970 726.540 2252.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2388.970 726.540 2392.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 726.540 2532.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 988.970 1261.540 992.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.970 1261.540 1132.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 1261.540 1272.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 1261.540 1412.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.970 1261.540 1552.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1828.970 -9.470 1832.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 1261.540 1972.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 1261.540 2112.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2388.970 1261.540 2392.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1261.540 2532.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 1261.540 292.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.970 1261.540 432.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 1261.540 572.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 1261.540 712.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.970 1261.540 852.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1828.970 1710.495 1832.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 1710.495 1972.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 1710.495 2112.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.970 1261.540 2252.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2388.970 1645.000 2392.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1645.000 2532.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 2135.165 292.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.970 2135.165 432.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 2135.165 572.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 2135.165 712.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.970 2135.165 852.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 988.970 2130.000 992.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.970 2130.000 1132.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 2130.000 1272.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 2130.000 1412.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.970 2130.000 1552.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 1261.540 1692.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 2145.495 1972.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 2145.495 2112.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.970 2145.495 2252.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2388.970 2145.495 2392.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 2145.495 2532.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 2691.540 292.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.970 2691.540 432.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 2691.540 572.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 2691.540 712.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.970 2691.540 852.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 988.970 2691.540 992.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.970 2691.540 1132.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 2691.540 1272.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 2691.540 1412.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.970 2691.540 1552.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 2691.540 1692.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 2691.540 1972.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 2691.540 2112.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.970 2691.540 2252.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2388.970 2691.540 2392.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 2691.540 2532.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 148.970 -9.470 152.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 3226.540 292.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.970 3226.540 432.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 3226.540 572.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 3226.540 712.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.970 3226.540 852.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 988.970 3226.540 992.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.970 3226.540 1132.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 3226.540 1272.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 3226.540 1412.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.970 3226.540 1552.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 3226.540 1692.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1828.970 2145.495 1832.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 3226.540 1972.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 3226.540 2112.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.970 3226.540 2252.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2388.970 3226.540 2392.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 3226.540 2532.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.970 -9.470 2672.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.970 -9.470 2812.070 3529.150 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 32.930 2944.050 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 172.930 2944.050 176.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 312.930 2944.050 316.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 452.930 2944.050 456.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 592.930 2944.050 596.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 732.930 2944.050 736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 872.930 2944.050 876.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1012.930 2944.050 1016.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1152.930 2944.050 1156.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1432.930 2944.050 1436.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1572.930 2944.050 1576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1712.930 2944.050 1716.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1852.930 2944.050 1856.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1992.930 2944.050 1996.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2132.930 2944.050 2136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 307.570 2198.230 730.670 2201.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1987.570 2198.230 2550.670 2201.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2272.930 2944.050 2276.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2412.930 2944.050 2416.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2692.930 2944.050 2696.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2832.930 2944.050 2836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2972.930 2944.050 2976.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3112.930 2944.050 3116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3252.930 2944.050 3256.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3392.930 2944.050 3396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 307.570 -19.070 310.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 447.570 -19.070 450.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 587.570 -19.070 590.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 -19.070 730.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 867.570 -19.070 870.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1147.570 -19.070 1150.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 -19.070 1290.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 -19.070 1430.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1567.570 -19.070 1570.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1707.570 -19.070 1710.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1987.570 -19.070 1990.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 -19.070 2130.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2267.570 -19.070 2270.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2407.570 -19.070 2410.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 -19.070 2550.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 307.570 726.540 310.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 447.570 726.540 450.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 587.570 726.540 590.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 726.540 730.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 867.570 726.540 870.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1147.570 726.540 1150.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 726.540 1290.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 726.540 1430.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1567.570 726.540 1570.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1707.570 726.540 1710.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1987.570 726.540 1990.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 726.540 2130.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2267.570 726.540 2270.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2407.570 726.540 2410.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 726.540 2550.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.570 -19.070 1010.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1147.570 1261.540 1150.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 1261.540 1290.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 1261.540 1430.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1567.570 1261.540 1570.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1847.570 -19.070 1850.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1987.570 1261.540 1990.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2407.570 1261.540 2410.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 1261.540 2550.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 307.570 1261.540 310.670 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 447.570 1261.540 450.670 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 587.570 1261.540 590.670 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 1261.540 730.670 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1847.570 1710.495 1850.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1987.570 1710.495 1990.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2267.570 1261.540 2270.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2407.570 1645.000 2410.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 1645.000 2550.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 307.570 2135.165 310.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 447.570 2135.165 450.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 587.570 2135.165 590.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 2135.165 730.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 867.570 1261.540 870.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1147.570 2130.000 1150.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 2130.000 1290.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 2130.000 1430.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1567.570 2130.000 1570.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1707.570 1261.540 1710.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1987.570 2145.495 1990.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 1261.540 2130.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2267.570 2145.495 2270.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2407.570 2145.495 2410.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 2145.495 2550.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 307.570 2691.540 310.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 447.570 2691.540 450.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 587.570 2691.540 590.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 2691.540 730.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 867.570 2691.540 870.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1147.570 2691.540 1150.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 2691.540 1290.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 2691.540 1430.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1567.570 2691.540 1570.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1707.570 2691.540 1710.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1987.570 2691.540 1990.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 2691.540 2130.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2267.570 2691.540 2270.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2407.570 2691.540 2410.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 2691.540 2550.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 167.570 -19.070 170.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 307.570 3226.540 310.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 447.570 3226.540 450.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 587.570 3226.540 590.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 3226.540 730.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 867.570 3226.540 870.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.570 2130.000 1010.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1147.570 3226.540 1150.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 3226.540 1290.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 3226.540 1430.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1567.570 3226.540 1570.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1707.570 3226.540 1710.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1847.570 2145.495 1850.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1987.570 3226.540 1990.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 3226.540 2130.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2267.570 3226.540 2270.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2407.570 3226.540 2410.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 3226.540 2550.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2687.570 -19.070 2690.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2827.570 -19.070 2830.670 3538.750 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 51.530 2953.650 54.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 191.530 2953.650 194.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 331.530 2953.650 334.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 471.530 2953.650 474.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 611.530 2953.650 614.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 751.530 2953.650 754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 891.530 2953.650 894.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1031.530 2953.650 1034.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1171.530 2953.650 1174.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1451.530 2953.650 1454.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1591.530 2953.650 1594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1731.530 2953.650 1734.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1871.530 2953.650 1874.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2011.530 2953.650 2014.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2151.530 2953.650 2154.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2291.530 2953.650 2294.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2431.530 2953.650 2434.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2711.530 2953.650 2714.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2851.530 2953.650 2854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2991.530 2953.650 2994.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3131.530 2953.650 3134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3271.530 2953.650 3274.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3411.530 2953.650 3414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.170 -28.670 329.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.170 -28.670 469.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.170 -28.670 609.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 -28.670 749.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.170 -28.670 889.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1166.170 -28.670 1169.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 -28.670 1309.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 -28.670 1449.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1586.170 -28.670 1589.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1726.170 -28.670 1729.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.170 -28.670 2009.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 -28.670 2149.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2286.170 -28.670 2289.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.170 -28.670 2429.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 -28.670 2569.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.170 726.540 329.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.170 726.540 469.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.170 726.540 609.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 726.540 749.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.170 726.540 889.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1166.170 726.540 1169.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 726.540 1309.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 726.540 1449.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1586.170 726.540 1589.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1726.170 726.540 1729.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.170 726.540 2009.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 726.540 2149.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2286.170 726.540 2289.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.170 726.540 2429.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 726.540 2569.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.170 -28.670 1029.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1166.170 1261.540 1169.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 1261.540 1309.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 1261.540 1449.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1586.170 1261.540 1589.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1866.170 -28.670 1869.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.170 1261.540 2009.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.170 1261.540 2429.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.170 1261.540 329.270 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.170 1261.540 469.270 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.170 1261.540 609.270 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 1261.540 749.270 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1866.170 1710.495 1869.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.170 1710.495 2009.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2286.170 1261.540 2289.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.170 1645.000 2429.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.170 2135.165 329.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.170 2135.165 469.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.170 2135.165 609.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 2135.165 749.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.170 1261.540 889.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1166.170 2130.000 1169.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 2130.000 1309.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 2130.000 1449.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1586.170 2130.000 1589.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1726.170 1261.540 1729.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.170 2145.495 2009.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 1261.540 2149.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2286.170 2145.495 2289.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.170 2145.495 2429.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 1261.540 2569.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.170 2691.540 329.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.170 2691.540 469.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.170 2691.540 609.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 2691.540 749.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.170 2691.540 889.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1166.170 2691.540 1169.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 2691.540 1309.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 2691.540 1449.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1586.170 2691.540 1589.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1726.170 2691.540 1729.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.170 2691.540 2009.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 2691.540 2149.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2286.170 2691.540 2289.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.170 2691.540 2429.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 2691.540 2569.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.170 -28.670 189.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.170 3226.540 329.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.170 3226.540 469.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.170 3226.540 609.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 3226.540 749.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.170 3226.540 889.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.170 2130.000 1029.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1166.170 3226.540 1169.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 3226.540 1309.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 3226.540 1449.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1586.170 3226.540 1589.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1726.170 3226.540 1729.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1866.170 2145.495 1869.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2006.170 3226.540 2009.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 3226.540 2149.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2286.170 3226.540 2289.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.170 3226.540 2429.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 3226.540 2569.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2706.170 -28.670 2709.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2846.170 -28.670 2849.270 3548.350 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 210.130 2963.250 213.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 350.130 2963.250 353.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 490.130 2963.250 493.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 630.130 2963.250 633.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 770.130 2963.250 773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 910.130 2963.250 913.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1050.130 2963.250 1053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1190.130 2963.250 1193.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1470.130 2963.250 1473.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1610.130 2963.250 1613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1750.130 2963.250 1753.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1890.130 2963.250 1893.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2030.130 2963.250 2033.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2170.130 2963.250 2173.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2310.130 2963.250 2313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2450.130 2963.250 2453.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2730.130 2963.250 2733.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2870.130 2963.250 2873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3010.130 2963.250 3013.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3150.130 2963.250 3153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3290.130 2963.250 3293.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3430.130 2963.250 3433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.770 -38.270 347.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.770 -38.270 487.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.770 -38.270 627.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 -38.270 767.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.770 -38.270 907.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.770 -38.270 1187.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 -38.270 1327.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 -38.270 1467.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.770 -38.270 1607.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1744.770 -38.270 1747.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.770 -38.270 2027.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 -38.270 2167.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.770 -38.270 2307.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2444.770 -38.270 2447.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 -38.270 2587.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.770 726.540 347.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.770 726.540 487.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.770 726.540 627.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 726.540 767.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.770 726.540 907.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.770 726.540 1187.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 726.540 1327.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 726.540 1467.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.770 726.540 1607.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1744.770 726.540 1747.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.770 726.540 2027.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 726.540 2167.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.770 726.540 2307.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2444.770 726.540 2447.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 726.540 2587.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1044.770 -38.270 1047.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.770 1261.540 1187.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 1261.540 1327.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 1261.540 1467.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.770 1261.540 1607.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1884.770 -38.270 1887.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.770 1261.540 2027.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.770 1261.540 2307.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2444.770 1261.540 2447.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.770 1261.540 347.870 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.770 1261.540 487.870 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.770 1261.540 627.870 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 1261.540 767.870 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1884.770 1710.495 1887.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.770 1710.495 2027.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.770 1645.000 2307.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2444.770 1645.000 2447.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.770 2135.165 347.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.770 2135.165 487.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.770 2135.165 627.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 2135.165 767.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.770 1261.540 907.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.770 2130.000 1187.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 2130.000 1327.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 2130.000 1467.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.770 2130.000 1607.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1744.770 1261.540 1747.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.770 2145.495 2027.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 1261.540 2167.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.770 2145.495 2307.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2444.770 2145.495 2447.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 1261.540 2587.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.770 2691.540 347.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.770 2691.540 487.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.770 2691.540 627.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 2691.540 767.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.770 2691.540 907.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.770 2691.540 1187.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 2691.540 1327.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 2691.540 1467.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.770 2691.540 1607.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1744.770 2691.540 1747.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.770 2691.540 2027.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 2691.540 2167.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.770 2691.540 2307.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2444.770 2691.540 2447.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 2691.540 2587.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.770 -38.270 207.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.770 3226.540 347.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.770 3226.540 487.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.770 3226.540 627.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 3226.540 767.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.770 3226.540 907.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1044.770 2130.000 1047.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.770 3226.540 1187.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 3226.540 1327.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 3226.540 1467.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.770 3226.540 1607.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1744.770 3226.540 1747.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1884.770 2145.495 1887.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.770 3226.540 2027.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 3226.540 2167.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.770 3226.540 2307.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2444.770 3226.540 2447.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 3226.540 2587.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2724.770 -38.270 2727.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2864.770 -38.270 2867.870 3557.950 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 121.530 2953.650 124.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 261.530 2953.650 264.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 401.530 2953.650 404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 541.530 2953.650 544.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 681.530 2953.650 684.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 821.530 2953.650 824.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 961.530 2953.650 964.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1101.530 2953.650 1104.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1241.530 2953.650 1244.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 1096.170 1316.230 1519.270 1319.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1936.170 1316.230 2499.270 1319.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1381.530 2953.650 1384.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1521.530 2953.650 1524.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1661.530 2953.650 1664.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1801.530 2953.650 1804.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2081.530 2953.650 2084.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2221.530 2953.650 2224.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2361.530 2953.650 2364.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2501.530 2953.650 2504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2641.530 2953.650 2644.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2781.530 2953.650 2784.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2921.530 2953.650 2924.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3061.530 2953.650 3064.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3341.530 2953.650 3344.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3481.530 2953.650 3484.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 -28.670 399.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.170 -28.670 539.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 -28.670 679.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.170 -28.670 819.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.170 -28.670 959.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 -28.670 1099.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1236.170 -28.670 1239.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1376.170 -28.670 1379.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.170 -28.670 1519.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1656.170 -28.670 1659.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 -28.670 1939.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2076.170 -28.670 2079.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.170 -28.670 2219.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.170 -28.670 2359.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 -28.670 2499.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 726.540 399.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.170 726.540 539.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 726.540 679.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.170 726.540 819.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.170 726.540 959.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 726.540 1099.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1236.170 726.540 1239.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1376.170 726.540 1379.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.170 726.540 1519.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1656.170 726.540 1659.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 726.540 1939.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2076.170 726.540 2079.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.170 726.540 2219.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.170 726.540 2359.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 726.540 2499.270 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 1261.540 1099.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1236.170 1261.540 1239.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1376.170 1261.540 1379.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.170 1261.540 1519.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1796.170 -28.670 1799.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 1261.540 1939.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2076.170 1261.540 2079.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.170 1261.540 2359.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 1261.540 2499.270 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 1261.540 399.270 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.170 1261.540 539.270 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 1261.540 679.270 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.170 1261.540 819.270 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1796.170 1710.495 1799.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 1710.495 1939.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2076.170 1710.495 2079.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.170 1645.000 2359.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 1645.000 2499.270 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 2135.165 399.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.170 2135.165 539.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 2135.165 679.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.170 2135.165 819.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.170 1261.540 959.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 2130.000 1099.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1236.170 2130.000 1239.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1376.170 2130.000 1379.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.170 2130.000 1519.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1656.170 1261.540 1659.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 2145.495 1939.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2076.170 2145.495 2079.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.170 1261.540 2219.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.170 2145.495 2359.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 2145.495 2499.270 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 2691.540 399.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.170 2691.540 539.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 2691.540 679.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.170 2691.540 819.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.170 2691.540 959.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 2691.540 1099.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1236.170 2691.540 1239.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1376.170 2691.540 1379.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.170 2691.540 1519.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1656.170 2691.540 1659.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 2691.540 1939.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2076.170 2691.540 2079.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.170 2691.540 2219.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.170 2691.540 2359.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 2691.540 2499.270 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.170 -28.670 119.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.170 -28.670 259.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 3226.540 399.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.170 3226.540 539.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 3226.540 679.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.170 3226.540 819.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.170 3226.540 959.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 3226.540 1099.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1236.170 3226.540 1239.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1376.170 3226.540 1379.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.170 3226.540 1519.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1656.170 3226.540 1659.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1796.170 2145.495 1799.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 3226.540 1939.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2076.170 3226.540 2079.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.170 3226.540 2219.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.170 3226.540 2359.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 3226.540 2499.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2636.170 -28.670 2639.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2776.170 -28.670 2779.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 140.130 2963.250 143.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 280.130 2963.250 283.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 420.130 2963.250 423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 560.130 2963.250 563.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 700.130 2963.250 703.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 414.770 774.830 2517.870 777.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 840.130 2963.250 843.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 980.130 2963.250 983.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1120.130 2963.250 1123.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1260.130 2963.250 1263.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 1114.770 1325.430 1537.870 1328.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 1954.770 1325.430 2517.870 1328.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1400.130 2963.250 1403.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1540.130 2963.250 1543.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1680.130 2963.250 1683.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 1814.770 1754.830 2097.870 1757.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1820.130 2963.250 1823.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2100.130 2963.250 2103.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2240.130 2963.250 2243.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2380.130 2963.250 2383.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2520.130 2963.250 2523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2660.130 2963.250 2663.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 414.770 2734.830 2517.870 2737.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2800.130 2963.250 2803.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2940.130 2963.250 2943.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3080.130 2963.250 3083.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3360.130 2963.250 3363.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3500.130 2963.250 3503.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 -38.270 417.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.770 -38.270 557.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 -38.270 697.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.770 -38.270 837.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.770 -38.270 977.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 -38.270 1117.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.770 -38.270 1257.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1394.770 -38.270 1397.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.770 -38.270 1537.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1674.770 -38.270 1677.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 -38.270 1957.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.770 -38.270 2097.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2234.770 -38.270 2237.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.770 -38.270 2377.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 -38.270 2517.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 726.540 417.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.770 726.540 557.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 726.540 697.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.770 726.540 837.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.770 726.540 977.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 726.540 1117.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.770 726.540 1257.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1394.770 726.540 1397.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.770 726.540 1537.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1674.770 726.540 1677.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 726.540 1957.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.770 726.540 2097.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2234.770 726.540 2237.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.770 726.540 2377.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 726.540 2517.870 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 1261.540 1117.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.770 1261.540 1257.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1394.770 1261.540 1397.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.770 1261.540 1537.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.770 -38.270 1817.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 1261.540 1957.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.770 1261.540 2097.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.770 1261.540 2377.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 1261.540 2517.870 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 1261.540 417.870 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.770 1261.540 557.870 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 1261.540 697.870 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.770 1261.540 837.870 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.770 1710.495 1817.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 1710.495 1957.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.770 1710.495 2097.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.770 1645.000 2377.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 1645.000 2517.870 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 2135.165 417.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.770 2135.165 557.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 2135.165 697.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.770 2135.165 837.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.770 1261.540 977.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 2130.000 1117.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.770 2130.000 1257.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1394.770 2130.000 1397.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.770 2130.000 1537.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1674.770 1261.540 1677.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 2145.495 1957.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.770 2145.495 2097.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2234.770 1261.540 2237.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.770 2145.495 2377.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 2145.495 2517.870 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 2691.540 417.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.770 2691.540 557.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 2691.540 697.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.770 2691.540 837.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.770 2691.540 977.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 2691.540 1117.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.770 2691.540 1257.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1394.770 2691.540 1397.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.770 2691.540 1537.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1674.770 2691.540 1677.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 2691.540 1957.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.770 2691.540 2097.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2234.770 2691.540 2237.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.770 2691.540 2377.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 2691.540 2517.870 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.770 -38.270 137.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.770 -38.270 277.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 3226.540 417.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.770 3226.540 557.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 3226.540 697.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.770 3226.540 837.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.770 3226.540 977.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 3226.540 1117.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.770 3226.540 1257.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1394.770 3226.540 1397.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.770 3226.540 1537.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1674.770 3226.540 1677.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.770 2145.495 1817.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 3226.540 1957.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.770 3226.540 2097.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2234.770 3226.540 2237.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.770 3226.540 2377.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 3226.540 2517.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.770 -38.270 2657.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2794.770 -38.270 2797.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 84.330 2934.450 87.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 224.330 2934.450 227.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 364.330 2934.450 367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 504.330 2934.450 507.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 644.330 2934.450 647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 784.330 2934.450 787.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 924.330 2934.450 927.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1064.330 2934.450 1067.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1204.330 2934.450 1207.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1344.330 2934.450 1347.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1484.330 2934.450 1487.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1624.330 2934.450 1627.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1764.330 2934.450 1767.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1904.330 2934.450 1907.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2044.330 2934.450 2047.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2184.330 2934.450 2187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2324.330 2934.450 2327.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2464.330 2934.450 2467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2604.330 2934.450 2607.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2744.330 2934.450 2747.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2884.330 2934.450 2887.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3024.330 2934.450 3027.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3164.330 2934.450 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3304.330 2934.450 3307.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3444.330 2934.450 3447.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 -9.470 362.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.970 -9.470 502.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 -9.470 642.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 778.970 -9.470 782.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 918.970 -9.470 922.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.970 -9.470 1202.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1338.970 -9.470 1342.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1478.970 -9.470 1482.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1618.970 -9.470 1622.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.970 -9.470 1762.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 -9.470 1902.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2038.970 -9.470 2042.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2178.970 -9.470 2182.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2318.970 -9.470 2322.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 -9.470 2462.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 726.540 362.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.970 726.540 502.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 726.540 642.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 778.970 726.540 782.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 918.970 726.540 922.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.970 726.540 1202.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1338.970 726.540 1342.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1478.970 726.540 1482.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1618.970 726.540 1622.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.970 726.540 1762.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 726.540 1902.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2038.970 726.540 2042.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2178.970 726.540 2182.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2318.970 726.540 2322.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 726.540 2462.070 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.970 -9.470 1062.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.970 1261.540 1202.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1338.970 1261.540 1342.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1478.970 1261.540 1482.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 1261.540 1902.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2038.970 1261.540 2042.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2318.970 1261.540 2322.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 1261.540 2462.070 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 1261.540 362.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.970 1261.540 502.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1261.540 642.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 778.970 1261.540 782.070 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 1710.495 1902.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2038.970 1710.495 2042.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2318.970 1645.000 2322.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 1645.000 2462.070 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 2135.165 362.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.970 2135.165 502.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2135.165 642.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 778.970 2135.165 782.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 918.970 1261.540 922.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.970 2130.000 1202.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1338.970 2130.000 1342.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1478.970 2130.000 1482.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1618.970 1261.540 1622.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.970 1261.540 1762.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 2145.495 1902.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2038.970 2145.495 2042.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2178.970 1261.540 2182.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2318.970 2145.495 2322.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 2145.495 2462.070 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 2691.540 362.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.970 2691.540 502.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2691.540 642.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 778.970 2691.540 782.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 918.970 2691.540 922.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.970 2691.540 1202.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1338.970 2691.540 1342.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1478.970 2691.540 1482.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1618.970 2691.540 1622.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.970 2691.540 1762.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 2691.540 1902.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2038.970 2691.540 2042.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2178.970 2691.540 2182.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2318.970 2691.540 2322.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 2691.540 2462.070 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 -9.470 82.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.970 -9.470 222.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 3226.540 362.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.970 3226.540 502.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 3226.540 642.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 778.970 3226.540 782.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 918.970 3226.540 922.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.970 2130.000 1062.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.970 3226.540 1202.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1338.970 3226.540 1342.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1478.970 3226.540 1482.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1618.970 3226.540 1622.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.970 3226.540 1762.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 3226.540 1902.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2038.970 3226.540 2042.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2178.970 3226.540 2182.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2318.970 3226.540 2322.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 3226.540 2462.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2598.970 -9.470 2602.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2738.970 -9.470 2742.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2878.970 -9.470 2882.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 102.930 2944.050 106.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 242.930 2944.050 246.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 382.930 2944.050 386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 522.930 2944.050 526.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 662.930 2944.050 666.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 802.930 2944.050 806.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 942.930 2944.050 946.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1082.930 2944.050 1086.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1222.930 2944.050 1226.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1362.930 2944.050 1366.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1502.930 2944.050 1506.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1642.930 2944.050 1646.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1782.930 2944.050 1786.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2062.930 2944.050 2066.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2202.930 2944.050 2206.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2342.930 2944.050 2346.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2482.930 2944.050 2486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2622.930 2944.050 2626.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2762.930 2944.050 2766.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2902.930 2944.050 2906.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3042.930 2944.050 3046.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3322.930 2944.050 3326.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3462.930 2944.050 3466.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 -19.070 380.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 517.570 -19.070 520.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 -19.070 660.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.570 -19.070 800.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 937.570 -19.070 940.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.570 -19.070 1220.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1357.570 -19.070 1360.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1497.570 -19.070 1500.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1637.570 -19.070 1640.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1777.570 -19.070 1780.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 -19.070 1920.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.570 -19.070 2060.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2197.570 -19.070 2200.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.570 -19.070 2340.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 -19.070 2480.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 726.540 380.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 517.570 726.540 520.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 726.540 660.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.570 726.540 800.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 937.570 726.540 940.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.570 726.540 1220.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1357.570 726.540 1360.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1497.570 726.540 1500.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1637.570 726.540 1640.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1777.570 726.540 1780.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 726.540 1920.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.570 726.540 2060.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2197.570 726.540 2200.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.570 726.540 2340.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 726.540 2480.670 825.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1077.570 -19.070 1080.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.570 1261.540 1220.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1357.570 1261.540 1360.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1497.570 1261.540 1500.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 1261.540 1920.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.570 1261.540 2060.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.570 1261.540 2340.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 1261.540 2480.670 1375.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 1261.540 380.670 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 517.570 1261.540 520.670 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 1261.540 660.670 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.570 1261.540 800.670 1560.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 1710.495 1920.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.570 1710.495 2060.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.570 1645.000 2340.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 1645.000 2480.670 1810.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 2135.165 380.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 517.570 2135.165 520.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 2135.165 660.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.570 2135.165 800.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 937.570 1261.540 940.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.570 2130.000 1220.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1357.570 2130.000 1360.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1497.570 2130.000 1500.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1637.570 1261.540 1640.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1777.570 1261.540 1780.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 2145.495 1920.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.570 2145.495 2060.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2197.570 1261.540 2200.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.570 2145.495 2340.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 2145.495 2480.670 2255.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 2691.540 380.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 517.570 2691.540 520.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 2691.540 660.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.570 2691.540 800.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 937.570 2691.540 940.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.570 2691.540 1220.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1357.570 2691.540 1360.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1497.570 2691.540 1500.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1637.570 2691.540 1640.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1777.570 2691.540 1780.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 2691.540 1920.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.570 2691.540 2060.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2197.570 2691.540 2200.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.570 2691.540 2340.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 2691.540 2480.670 2790.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.570 -19.070 100.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.570 -19.070 240.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 3226.540 380.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 517.570 3226.540 520.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 3226.540 660.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.570 3226.540 800.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 937.570 3226.540 940.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1077.570 2130.000 1080.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.570 3226.540 1220.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1357.570 3226.540 1360.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1497.570 3226.540 1500.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1637.570 3226.540 1640.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1777.570 3226.540 1780.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 3226.540 1920.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.570 3226.540 2060.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2197.570 3226.540 2200.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.570 3226.540 2340.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 3226.540 2480.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2617.570 -19.070 2620.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2757.570 -19.070 2760.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2897.570 -19.070 2900.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 305.520 1395.795 2549.000 2122.005 ;
      LAYER met1 ;
        RECT 2.830 17.040 2902.070 3501.960 ;
      LAYER met2 ;
        RECT 2.860 3517.320 40.150 3518.050 ;
        RECT 41.270 3517.320 121.110 3518.050 ;
        RECT 122.230 3517.320 202.070 3518.050 ;
        RECT 203.190 3517.320 283.490 3518.050 ;
        RECT 284.610 3517.320 364.450 3518.050 ;
        RECT 365.570 3517.320 445.410 3518.050 ;
        RECT 446.530 3517.320 526.830 3518.050 ;
        RECT 527.950 3517.320 607.790 3518.050 ;
        RECT 608.910 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 770.170 3518.050 ;
        RECT 771.290 3517.320 851.130 3518.050 ;
        RECT 852.250 3517.320 932.090 3518.050 ;
        RECT 933.210 3517.320 1013.510 3518.050 ;
        RECT 1014.630 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1175.430 3518.050 ;
        RECT 1176.550 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1500.190 3518.050 ;
        RECT 1501.310 3517.320 1581.150 3518.050 ;
        RECT 1582.270 3517.320 1662.110 3518.050 ;
        RECT 1663.230 3517.320 1743.530 3518.050 ;
        RECT 1744.650 3517.320 1824.490 3518.050 ;
        RECT 1825.610 3517.320 1905.450 3518.050 ;
        RECT 1906.570 3517.320 1986.870 3518.050 ;
        RECT 1987.990 3517.320 2067.830 3518.050 ;
        RECT 2068.950 3517.320 2148.790 3518.050 ;
        RECT 2149.910 3517.320 2230.210 3518.050 ;
        RECT 2231.330 3517.320 2311.170 3518.050 ;
        RECT 2312.290 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2554.510 3518.050 ;
        RECT 2555.630 3517.320 2635.470 3518.050 ;
        RECT 2636.590 3517.320 2716.890 3518.050 ;
        RECT 2718.010 3517.320 2797.850 3518.050 ;
        RECT 2798.970 3517.320 2878.810 3518.050 ;
        RECT 2879.930 3517.320 2902.050 3518.050 ;
        RECT 2.860 2.680 2902.050 3517.320 ;
        RECT 3.550 2.400 7.950 2.680 ;
        RECT 9.070 2.400 13.930 2.680 ;
        RECT 15.050 2.400 19.910 2.680 ;
        RECT 21.030 2.400 25.890 2.680 ;
        RECT 27.010 2.400 31.870 2.680 ;
        RECT 32.990 2.400 37.850 2.680 ;
        RECT 38.970 2.400 43.370 2.680 ;
        RECT 44.490 2.400 49.350 2.680 ;
        RECT 50.470 2.400 55.330 2.680 ;
        RECT 56.450 2.400 61.310 2.680 ;
        RECT 62.430 2.400 67.290 2.680 ;
        RECT 68.410 2.400 73.270 2.680 ;
        RECT 74.390 2.400 79.250 2.680 ;
        RECT 80.370 2.400 84.770 2.680 ;
        RECT 85.890 2.400 90.750 2.680 ;
        RECT 91.870 2.400 96.730 2.680 ;
        RECT 97.850 2.400 102.710 2.680 ;
        RECT 103.830 2.400 108.690 2.680 ;
        RECT 109.810 2.400 114.670 2.680 ;
        RECT 115.790 2.400 120.650 2.680 ;
        RECT 121.770 2.400 126.170 2.680 ;
        RECT 127.290 2.400 132.150 2.680 ;
        RECT 133.270 2.400 138.130 2.680 ;
        RECT 139.250 2.400 144.110 2.680 ;
        RECT 145.230 2.400 150.090 2.680 ;
        RECT 151.210 2.400 156.070 2.680 ;
        RECT 157.190 2.400 161.590 2.680 ;
        RECT 162.710 2.400 167.570 2.680 ;
        RECT 168.690 2.400 173.550 2.680 ;
        RECT 174.670 2.400 179.530 2.680 ;
        RECT 180.650 2.400 185.510 2.680 ;
        RECT 186.630 2.400 191.490 2.680 ;
        RECT 192.610 2.400 197.470 2.680 ;
        RECT 198.590 2.400 202.990 2.680 ;
        RECT 204.110 2.400 208.970 2.680 ;
        RECT 210.090 2.400 214.950 2.680 ;
        RECT 216.070 2.400 220.930 2.680 ;
        RECT 222.050 2.400 226.910 2.680 ;
        RECT 228.030 2.400 232.890 2.680 ;
        RECT 234.010 2.400 238.870 2.680 ;
        RECT 239.990 2.400 244.390 2.680 ;
        RECT 245.510 2.400 250.370 2.680 ;
        RECT 251.490 2.400 256.350 2.680 ;
        RECT 257.470 2.400 262.330 2.680 ;
        RECT 263.450 2.400 268.310 2.680 ;
        RECT 269.430 2.400 274.290 2.680 ;
        RECT 275.410 2.400 279.810 2.680 ;
        RECT 280.930 2.400 285.790 2.680 ;
        RECT 286.910 2.400 291.770 2.680 ;
        RECT 292.890 2.400 297.750 2.680 ;
        RECT 298.870 2.400 303.730 2.680 ;
        RECT 304.850 2.400 309.710 2.680 ;
        RECT 310.830 2.400 315.690 2.680 ;
        RECT 316.810 2.400 321.210 2.680 ;
        RECT 322.330 2.400 327.190 2.680 ;
        RECT 328.310 2.400 333.170 2.680 ;
        RECT 334.290 2.400 339.150 2.680 ;
        RECT 340.270 2.400 345.130 2.680 ;
        RECT 346.250 2.400 351.110 2.680 ;
        RECT 352.230 2.400 357.090 2.680 ;
        RECT 358.210 2.400 362.610 2.680 ;
        RECT 363.730 2.400 368.590 2.680 ;
        RECT 369.710 2.400 374.570 2.680 ;
        RECT 375.690 2.400 380.550 2.680 ;
        RECT 381.670 2.400 386.530 2.680 ;
        RECT 387.650 2.400 392.510 2.680 ;
        RECT 393.630 2.400 398.030 2.680 ;
        RECT 399.150 2.400 404.010 2.680 ;
        RECT 405.130 2.400 409.990 2.680 ;
        RECT 411.110 2.400 415.970 2.680 ;
        RECT 417.090 2.400 421.950 2.680 ;
        RECT 423.070 2.400 427.930 2.680 ;
        RECT 429.050 2.400 433.910 2.680 ;
        RECT 435.030 2.400 439.430 2.680 ;
        RECT 440.550 2.400 445.410 2.680 ;
        RECT 446.530 2.400 451.390 2.680 ;
        RECT 452.510 2.400 457.370 2.680 ;
        RECT 458.490 2.400 463.350 2.680 ;
        RECT 464.470 2.400 469.330 2.680 ;
        RECT 470.450 2.400 475.310 2.680 ;
        RECT 476.430 2.400 480.830 2.680 ;
        RECT 481.950 2.400 486.810 2.680 ;
        RECT 487.930 2.400 492.790 2.680 ;
        RECT 493.910 2.400 498.770 2.680 ;
        RECT 499.890 2.400 504.750 2.680 ;
        RECT 505.870 2.400 510.730 2.680 ;
        RECT 511.850 2.400 516.250 2.680 ;
        RECT 517.370 2.400 522.230 2.680 ;
        RECT 523.350 2.400 528.210 2.680 ;
        RECT 529.330 2.400 534.190 2.680 ;
        RECT 535.310 2.400 540.170 2.680 ;
        RECT 541.290 2.400 546.150 2.680 ;
        RECT 547.270 2.400 552.130 2.680 ;
        RECT 553.250 2.400 557.650 2.680 ;
        RECT 558.770 2.400 563.630 2.680 ;
        RECT 564.750 2.400 569.610 2.680 ;
        RECT 570.730 2.400 575.590 2.680 ;
        RECT 576.710 2.400 581.570 2.680 ;
        RECT 582.690 2.400 587.550 2.680 ;
        RECT 588.670 2.400 593.530 2.680 ;
        RECT 594.650 2.400 599.050 2.680 ;
        RECT 600.170 2.400 605.030 2.680 ;
        RECT 606.150 2.400 611.010 2.680 ;
        RECT 612.130 2.400 616.990 2.680 ;
        RECT 618.110 2.400 622.970 2.680 ;
        RECT 624.090 2.400 628.950 2.680 ;
        RECT 630.070 2.400 634.470 2.680 ;
        RECT 635.590 2.400 640.450 2.680 ;
        RECT 641.570 2.400 646.430 2.680 ;
        RECT 647.550 2.400 652.410 2.680 ;
        RECT 653.530 2.400 658.390 2.680 ;
        RECT 659.510 2.400 664.370 2.680 ;
        RECT 665.490 2.400 670.350 2.680 ;
        RECT 671.470 2.400 675.870 2.680 ;
        RECT 676.990 2.400 681.850 2.680 ;
        RECT 682.970 2.400 687.830 2.680 ;
        RECT 688.950 2.400 693.810 2.680 ;
        RECT 694.930 2.400 699.790 2.680 ;
        RECT 700.910 2.400 705.770 2.680 ;
        RECT 706.890 2.400 711.750 2.680 ;
        RECT 712.870 2.400 717.270 2.680 ;
        RECT 718.390 2.400 723.250 2.680 ;
        RECT 724.370 2.400 729.230 2.680 ;
        RECT 730.350 2.400 735.210 2.680 ;
        RECT 736.330 2.400 741.190 2.680 ;
        RECT 742.310 2.400 747.170 2.680 ;
        RECT 748.290 2.400 752.690 2.680 ;
        RECT 753.810 2.400 758.670 2.680 ;
        RECT 759.790 2.400 764.650 2.680 ;
        RECT 765.770 2.400 770.630 2.680 ;
        RECT 771.750 2.400 776.610 2.680 ;
        RECT 777.730 2.400 782.590 2.680 ;
        RECT 783.710 2.400 788.570 2.680 ;
        RECT 789.690 2.400 794.090 2.680 ;
        RECT 795.210 2.400 800.070 2.680 ;
        RECT 801.190 2.400 806.050 2.680 ;
        RECT 807.170 2.400 812.030 2.680 ;
        RECT 813.150 2.400 818.010 2.680 ;
        RECT 819.130 2.400 823.990 2.680 ;
        RECT 825.110 2.400 829.970 2.680 ;
        RECT 831.090 2.400 835.490 2.680 ;
        RECT 836.610 2.400 841.470 2.680 ;
        RECT 842.590 2.400 847.450 2.680 ;
        RECT 848.570 2.400 853.430 2.680 ;
        RECT 854.550 2.400 859.410 2.680 ;
        RECT 860.530 2.400 865.390 2.680 ;
        RECT 866.510 2.400 870.910 2.680 ;
        RECT 872.030 2.400 876.890 2.680 ;
        RECT 878.010 2.400 882.870 2.680 ;
        RECT 883.990 2.400 888.850 2.680 ;
        RECT 889.970 2.400 894.830 2.680 ;
        RECT 895.950 2.400 900.810 2.680 ;
        RECT 901.930 2.400 906.790 2.680 ;
        RECT 907.910 2.400 912.310 2.680 ;
        RECT 913.430 2.400 918.290 2.680 ;
        RECT 919.410 2.400 924.270 2.680 ;
        RECT 925.390 2.400 930.250 2.680 ;
        RECT 931.370 2.400 936.230 2.680 ;
        RECT 937.350 2.400 942.210 2.680 ;
        RECT 943.330 2.400 948.190 2.680 ;
        RECT 949.310 2.400 953.710 2.680 ;
        RECT 954.830 2.400 959.690 2.680 ;
        RECT 960.810 2.400 965.670 2.680 ;
        RECT 966.790 2.400 971.650 2.680 ;
        RECT 972.770 2.400 977.630 2.680 ;
        RECT 978.750 2.400 983.610 2.680 ;
        RECT 984.730 2.400 989.130 2.680 ;
        RECT 990.250 2.400 995.110 2.680 ;
        RECT 996.230 2.400 1001.090 2.680 ;
        RECT 1002.210 2.400 1007.070 2.680 ;
        RECT 1008.190 2.400 1013.050 2.680 ;
        RECT 1014.170 2.400 1019.030 2.680 ;
        RECT 1020.150 2.400 1025.010 2.680 ;
        RECT 1026.130 2.400 1030.530 2.680 ;
        RECT 1031.650 2.400 1036.510 2.680 ;
        RECT 1037.630 2.400 1042.490 2.680 ;
        RECT 1043.610 2.400 1048.470 2.680 ;
        RECT 1049.590 2.400 1054.450 2.680 ;
        RECT 1055.570 2.400 1060.430 2.680 ;
        RECT 1061.550 2.400 1066.410 2.680 ;
        RECT 1067.530 2.400 1071.930 2.680 ;
        RECT 1073.050 2.400 1077.910 2.680 ;
        RECT 1079.030 2.400 1083.890 2.680 ;
        RECT 1085.010 2.400 1089.870 2.680 ;
        RECT 1090.990 2.400 1095.850 2.680 ;
        RECT 1096.970 2.400 1101.830 2.680 ;
        RECT 1102.950 2.400 1107.350 2.680 ;
        RECT 1108.470 2.400 1113.330 2.680 ;
        RECT 1114.450 2.400 1119.310 2.680 ;
        RECT 1120.430 2.400 1125.290 2.680 ;
        RECT 1126.410 2.400 1131.270 2.680 ;
        RECT 1132.390 2.400 1137.250 2.680 ;
        RECT 1138.370 2.400 1143.230 2.680 ;
        RECT 1144.350 2.400 1148.750 2.680 ;
        RECT 1149.870 2.400 1154.730 2.680 ;
        RECT 1155.850 2.400 1160.710 2.680 ;
        RECT 1161.830 2.400 1166.690 2.680 ;
        RECT 1167.810 2.400 1172.670 2.680 ;
        RECT 1173.790 2.400 1178.650 2.680 ;
        RECT 1179.770 2.400 1184.630 2.680 ;
        RECT 1185.750 2.400 1190.150 2.680 ;
        RECT 1191.270 2.400 1196.130 2.680 ;
        RECT 1197.250 2.400 1202.110 2.680 ;
        RECT 1203.230 2.400 1208.090 2.680 ;
        RECT 1209.210 2.400 1214.070 2.680 ;
        RECT 1215.190 2.400 1220.050 2.680 ;
        RECT 1221.170 2.400 1225.570 2.680 ;
        RECT 1226.690 2.400 1231.550 2.680 ;
        RECT 1232.670 2.400 1237.530 2.680 ;
        RECT 1238.650 2.400 1243.510 2.680 ;
        RECT 1244.630 2.400 1249.490 2.680 ;
        RECT 1250.610 2.400 1255.470 2.680 ;
        RECT 1256.590 2.400 1261.450 2.680 ;
        RECT 1262.570 2.400 1266.970 2.680 ;
        RECT 1268.090 2.400 1272.950 2.680 ;
        RECT 1274.070 2.400 1278.930 2.680 ;
        RECT 1280.050 2.400 1284.910 2.680 ;
        RECT 1286.030 2.400 1290.890 2.680 ;
        RECT 1292.010 2.400 1296.870 2.680 ;
        RECT 1297.990 2.400 1302.850 2.680 ;
        RECT 1303.970 2.400 1308.370 2.680 ;
        RECT 1309.490 2.400 1314.350 2.680 ;
        RECT 1315.470 2.400 1320.330 2.680 ;
        RECT 1321.450 2.400 1326.310 2.680 ;
        RECT 1327.430 2.400 1332.290 2.680 ;
        RECT 1333.410 2.400 1338.270 2.680 ;
        RECT 1339.390 2.400 1343.790 2.680 ;
        RECT 1344.910 2.400 1349.770 2.680 ;
        RECT 1350.890 2.400 1355.750 2.680 ;
        RECT 1356.870 2.400 1361.730 2.680 ;
        RECT 1362.850 2.400 1367.710 2.680 ;
        RECT 1368.830 2.400 1373.690 2.680 ;
        RECT 1374.810 2.400 1379.670 2.680 ;
        RECT 1380.790 2.400 1385.190 2.680 ;
        RECT 1386.310 2.400 1391.170 2.680 ;
        RECT 1392.290 2.400 1397.150 2.680 ;
        RECT 1398.270 2.400 1403.130 2.680 ;
        RECT 1404.250 2.400 1409.110 2.680 ;
        RECT 1410.230 2.400 1415.090 2.680 ;
        RECT 1416.210 2.400 1421.070 2.680 ;
        RECT 1422.190 2.400 1426.590 2.680 ;
        RECT 1427.710 2.400 1432.570 2.680 ;
        RECT 1433.690 2.400 1438.550 2.680 ;
        RECT 1439.670 2.400 1444.530 2.680 ;
        RECT 1445.650 2.400 1450.510 2.680 ;
        RECT 1451.630 2.400 1456.490 2.680 ;
        RECT 1457.610 2.400 1462.470 2.680 ;
        RECT 1463.590 2.400 1467.990 2.680 ;
        RECT 1469.110 2.400 1473.970 2.680 ;
        RECT 1475.090 2.400 1479.950 2.680 ;
        RECT 1481.070 2.400 1485.930 2.680 ;
        RECT 1487.050 2.400 1491.910 2.680 ;
        RECT 1493.030 2.400 1497.890 2.680 ;
        RECT 1499.010 2.400 1503.410 2.680 ;
        RECT 1504.530 2.400 1509.390 2.680 ;
        RECT 1510.510 2.400 1515.370 2.680 ;
        RECT 1516.490 2.400 1521.350 2.680 ;
        RECT 1522.470 2.400 1527.330 2.680 ;
        RECT 1528.450 2.400 1533.310 2.680 ;
        RECT 1534.430 2.400 1539.290 2.680 ;
        RECT 1540.410 2.400 1544.810 2.680 ;
        RECT 1545.930 2.400 1550.790 2.680 ;
        RECT 1551.910 2.400 1556.770 2.680 ;
        RECT 1557.890 2.400 1562.750 2.680 ;
        RECT 1563.870 2.400 1568.730 2.680 ;
        RECT 1569.850 2.400 1574.710 2.680 ;
        RECT 1575.830 2.400 1580.690 2.680 ;
        RECT 1581.810 2.400 1586.210 2.680 ;
        RECT 1587.330 2.400 1592.190 2.680 ;
        RECT 1593.310 2.400 1598.170 2.680 ;
        RECT 1599.290 2.400 1604.150 2.680 ;
        RECT 1605.270 2.400 1610.130 2.680 ;
        RECT 1611.250 2.400 1616.110 2.680 ;
        RECT 1617.230 2.400 1621.630 2.680 ;
        RECT 1622.750 2.400 1627.610 2.680 ;
        RECT 1628.730 2.400 1633.590 2.680 ;
        RECT 1634.710 2.400 1639.570 2.680 ;
        RECT 1640.690 2.400 1645.550 2.680 ;
        RECT 1646.670 2.400 1651.530 2.680 ;
        RECT 1652.650 2.400 1657.510 2.680 ;
        RECT 1658.630 2.400 1663.030 2.680 ;
        RECT 1664.150 2.400 1669.010 2.680 ;
        RECT 1670.130 2.400 1674.990 2.680 ;
        RECT 1676.110 2.400 1680.970 2.680 ;
        RECT 1682.090 2.400 1686.950 2.680 ;
        RECT 1688.070 2.400 1692.930 2.680 ;
        RECT 1694.050 2.400 1698.910 2.680 ;
        RECT 1700.030 2.400 1704.430 2.680 ;
        RECT 1705.550 2.400 1710.410 2.680 ;
        RECT 1711.530 2.400 1716.390 2.680 ;
        RECT 1717.510 2.400 1722.370 2.680 ;
        RECT 1723.490 2.400 1728.350 2.680 ;
        RECT 1729.470 2.400 1734.330 2.680 ;
        RECT 1735.450 2.400 1739.850 2.680 ;
        RECT 1740.970 2.400 1745.830 2.680 ;
        RECT 1746.950 2.400 1751.810 2.680 ;
        RECT 1752.930 2.400 1757.790 2.680 ;
        RECT 1758.910 2.400 1763.770 2.680 ;
        RECT 1764.890 2.400 1769.750 2.680 ;
        RECT 1770.870 2.400 1775.730 2.680 ;
        RECT 1776.850 2.400 1781.250 2.680 ;
        RECT 1782.370 2.400 1787.230 2.680 ;
        RECT 1788.350 2.400 1793.210 2.680 ;
        RECT 1794.330 2.400 1799.190 2.680 ;
        RECT 1800.310 2.400 1805.170 2.680 ;
        RECT 1806.290 2.400 1811.150 2.680 ;
        RECT 1812.270 2.400 1817.130 2.680 ;
        RECT 1818.250 2.400 1822.650 2.680 ;
        RECT 1823.770 2.400 1828.630 2.680 ;
        RECT 1829.750 2.400 1834.610 2.680 ;
        RECT 1835.730 2.400 1840.590 2.680 ;
        RECT 1841.710 2.400 1846.570 2.680 ;
        RECT 1847.690 2.400 1852.550 2.680 ;
        RECT 1853.670 2.400 1858.070 2.680 ;
        RECT 1859.190 2.400 1864.050 2.680 ;
        RECT 1865.170 2.400 1870.030 2.680 ;
        RECT 1871.150 2.400 1876.010 2.680 ;
        RECT 1877.130 2.400 1881.990 2.680 ;
        RECT 1883.110 2.400 1887.970 2.680 ;
        RECT 1889.090 2.400 1893.950 2.680 ;
        RECT 1895.070 2.400 1899.470 2.680 ;
        RECT 1900.590 2.400 1905.450 2.680 ;
        RECT 1906.570 2.400 1911.430 2.680 ;
        RECT 1912.550 2.400 1917.410 2.680 ;
        RECT 1918.530 2.400 1923.390 2.680 ;
        RECT 1924.510 2.400 1929.370 2.680 ;
        RECT 1930.490 2.400 1935.350 2.680 ;
        RECT 1936.470 2.400 1940.870 2.680 ;
        RECT 1941.990 2.400 1946.850 2.680 ;
        RECT 1947.970 2.400 1952.830 2.680 ;
        RECT 1953.950 2.400 1958.810 2.680 ;
        RECT 1959.930 2.400 1964.790 2.680 ;
        RECT 1965.910 2.400 1970.770 2.680 ;
        RECT 1971.890 2.400 1976.290 2.680 ;
        RECT 1977.410 2.400 1982.270 2.680 ;
        RECT 1983.390 2.400 1988.250 2.680 ;
        RECT 1989.370 2.400 1994.230 2.680 ;
        RECT 1995.350 2.400 2000.210 2.680 ;
        RECT 2001.330 2.400 2006.190 2.680 ;
        RECT 2007.310 2.400 2012.170 2.680 ;
        RECT 2013.290 2.400 2017.690 2.680 ;
        RECT 2018.810 2.400 2023.670 2.680 ;
        RECT 2024.790 2.400 2029.650 2.680 ;
        RECT 2030.770 2.400 2035.630 2.680 ;
        RECT 2036.750 2.400 2041.610 2.680 ;
        RECT 2042.730 2.400 2047.590 2.680 ;
        RECT 2048.710 2.400 2053.570 2.680 ;
        RECT 2054.690 2.400 2059.090 2.680 ;
        RECT 2060.210 2.400 2065.070 2.680 ;
        RECT 2066.190 2.400 2071.050 2.680 ;
        RECT 2072.170 2.400 2077.030 2.680 ;
        RECT 2078.150 2.400 2083.010 2.680 ;
        RECT 2084.130 2.400 2088.990 2.680 ;
        RECT 2090.110 2.400 2094.510 2.680 ;
        RECT 2095.630 2.400 2100.490 2.680 ;
        RECT 2101.610 2.400 2106.470 2.680 ;
        RECT 2107.590 2.400 2112.450 2.680 ;
        RECT 2113.570 2.400 2118.430 2.680 ;
        RECT 2119.550 2.400 2124.410 2.680 ;
        RECT 2125.530 2.400 2130.390 2.680 ;
        RECT 2131.510 2.400 2135.910 2.680 ;
        RECT 2137.030 2.400 2141.890 2.680 ;
        RECT 2143.010 2.400 2147.870 2.680 ;
        RECT 2148.990 2.400 2153.850 2.680 ;
        RECT 2154.970 2.400 2159.830 2.680 ;
        RECT 2160.950 2.400 2165.810 2.680 ;
        RECT 2166.930 2.400 2171.790 2.680 ;
        RECT 2172.910 2.400 2177.310 2.680 ;
        RECT 2178.430 2.400 2183.290 2.680 ;
        RECT 2184.410 2.400 2189.270 2.680 ;
        RECT 2190.390 2.400 2195.250 2.680 ;
        RECT 2196.370 2.400 2201.230 2.680 ;
        RECT 2202.350 2.400 2207.210 2.680 ;
        RECT 2208.330 2.400 2212.730 2.680 ;
        RECT 2213.850 2.400 2218.710 2.680 ;
        RECT 2219.830 2.400 2224.690 2.680 ;
        RECT 2225.810 2.400 2230.670 2.680 ;
        RECT 2231.790 2.400 2236.650 2.680 ;
        RECT 2237.770 2.400 2242.630 2.680 ;
        RECT 2243.750 2.400 2248.610 2.680 ;
        RECT 2249.730 2.400 2254.130 2.680 ;
        RECT 2255.250 2.400 2260.110 2.680 ;
        RECT 2261.230 2.400 2266.090 2.680 ;
        RECT 2267.210 2.400 2272.070 2.680 ;
        RECT 2273.190 2.400 2278.050 2.680 ;
        RECT 2279.170 2.400 2284.030 2.680 ;
        RECT 2285.150 2.400 2290.010 2.680 ;
        RECT 2291.130 2.400 2295.530 2.680 ;
        RECT 2296.650 2.400 2301.510 2.680 ;
        RECT 2302.630 2.400 2307.490 2.680 ;
        RECT 2308.610 2.400 2313.470 2.680 ;
        RECT 2314.590 2.400 2319.450 2.680 ;
        RECT 2320.570 2.400 2325.430 2.680 ;
        RECT 2326.550 2.400 2330.950 2.680 ;
        RECT 2332.070 2.400 2336.930 2.680 ;
        RECT 2338.050 2.400 2342.910 2.680 ;
        RECT 2344.030 2.400 2348.890 2.680 ;
        RECT 2350.010 2.400 2354.870 2.680 ;
        RECT 2355.990 2.400 2360.850 2.680 ;
        RECT 2361.970 2.400 2366.830 2.680 ;
        RECT 2367.950 2.400 2372.350 2.680 ;
        RECT 2373.470 2.400 2378.330 2.680 ;
        RECT 2379.450 2.400 2384.310 2.680 ;
        RECT 2385.430 2.400 2390.290 2.680 ;
        RECT 2391.410 2.400 2396.270 2.680 ;
        RECT 2397.390 2.400 2402.250 2.680 ;
        RECT 2403.370 2.400 2408.230 2.680 ;
        RECT 2409.350 2.400 2413.750 2.680 ;
        RECT 2414.870 2.400 2419.730 2.680 ;
        RECT 2420.850 2.400 2425.710 2.680 ;
        RECT 2426.830 2.400 2431.690 2.680 ;
        RECT 2432.810 2.400 2437.670 2.680 ;
        RECT 2438.790 2.400 2443.650 2.680 ;
        RECT 2444.770 2.400 2449.170 2.680 ;
        RECT 2450.290 2.400 2455.150 2.680 ;
        RECT 2456.270 2.400 2461.130 2.680 ;
        RECT 2462.250 2.400 2467.110 2.680 ;
        RECT 2468.230 2.400 2473.090 2.680 ;
        RECT 2474.210 2.400 2479.070 2.680 ;
        RECT 2480.190 2.400 2485.050 2.680 ;
        RECT 2486.170 2.400 2490.570 2.680 ;
        RECT 2491.690 2.400 2496.550 2.680 ;
        RECT 2497.670 2.400 2502.530 2.680 ;
        RECT 2503.650 2.400 2508.510 2.680 ;
        RECT 2509.630 2.400 2514.490 2.680 ;
        RECT 2515.610 2.400 2520.470 2.680 ;
        RECT 2521.590 2.400 2526.450 2.680 ;
        RECT 2527.570 2.400 2531.970 2.680 ;
        RECT 2533.090 2.400 2537.950 2.680 ;
        RECT 2539.070 2.400 2543.930 2.680 ;
        RECT 2545.050 2.400 2549.910 2.680 ;
        RECT 2551.030 2.400 2555.890 2.680 ;
        RECT 2557.010 2.400 2561.870 2.680 ;
        RECT 2562.990 2.400 2567.390 2.680 ;
        RECT 2568.510 2.400 2573.370 2.680 ;
        RECT 2574.490 2.400 2579.350 2.680 ;
        RECT 2580.470 2.400 2585.330 2.680 ;
        RECT 2586.450 2.400 2591.310 2.680 ;
        RECT 2592.430 2.400 2597.290 2.680 ;
        RECT 2598.410 2.400 2603.270 2.680 ;
        RECT 2604.390 2.400 2608.790 2.680 ;
        RECT 2609.910 2.400 2614.770 2.680 ;
        RECT 2615.890 2.400 2620.750 2.680 ;
        RECT 2621.870 2.400 2626.730 2.680 ;
        RECT 2627.850 2.400 2632.710 2.680 ;
        RECT 2633.830 2.400 2638.690 2.680 ;
        RECT 2639.810 2.400 2644.670 2.680 ;
        RECT 2645.790 2.400 2650.190 2.680 ;
        RECT 2651.310 2.400 2656.170 2.680 ;
        RECT 2657.290 2.400 2662.150 2.680 ;
        RECT 2663.270 2.400 2668.130 2.680 ;
        RECT 2669.250 2.400 2674.110 2.680 ;
        RECT 2675.230 2.400 2680.090 2.680 ;
        RECT 2681.210 2.400 2685.610 2.680 ;
        RECT 2686.730 2.400 2691.590 2.680 ;
        RECT 2692.710 2.400 2697.570 2.680 ;
        RECT 2698.690 2.400 2703.550 2.680 ;
        RECT 2704.670 2.400 2709.530 2.680 ;
        RECT 2710.650 2.400 2715.510 2.680 ;
        RECT 2716.630 2.400 2721.490 2.680 ;
        RECT 2722.610 2.400 2727.010 2.680 ;
        RECT 2728.130 2.400 2732.990 2.680 ;
        RECT 2734.110 2.400 2738.970 2.680 ;
        RECT 2740.090 2.400 2744.950 2.680 ;
        RECT 2746.070 2.400 2750.930 2.680 ;
        RECT 2752.050 2.400 2756.910 2.680 ;
        RECT 2758.030 2.400 2762.890 2.680 ;
        RECT 2764.010 2.400 2768.410 2.680 ;
        RECT 2769.530 2.400 2774.390 2.680 ;
        RECT 2775.510 2.400 2780.370 2.680 ;
        RECT 2781.490 2.400 2786.350 2.680 ;
        RECT 2787.470 2.400 2792.330 2.680 ;
        RECT 2793.450 2.400 2798.310 2.680 ;
        RECT 2799.430 2.400 2803.830 2.680 ;
        RECT 2804.950 2.400 2809.810 2.680 ;
        RECT 2810.930 2.400 2815.790 2.680 ;
        RECT 2816.910 2.400 2821.770 2.680 ;
        RECT 2822.890 2.400 2827.750 2.680 ;
        RECT 2828.870 2.400 2833.730 2.680 ;
        RECT 2834.850 2.400 2839.710 2.680 ;
        RECT 2840.830 2.400 2845.230 2.680 ;
        RECT 2846.350 2.400 2851.210 2.680 ;
        RECT 2852.330 2.400 2857.190 2.680 ;
        RECT 2858.310 2.400 2863.170 2.680 ;
        RECT 2864.290 2.400 2869.150 2.680 ;
        RECT 2870.270 2.400 2875.130 2.680 ;
        RECT 2876.250 2.400 2881.110 2.680 ;
        RECT 2882.230 2.400 2886.630 2.680 ;
        RECT 2887.750 2.400 2892.610 2.680 ;
        RECT 2893.730 2.400 2898.590 2.680 ;
        RECT 2899.710 2.400 2902.050 2.680 ;
      LAYER met3 ;
        RECT 2.400 3487.700 2917.930 3501.825 ;
        RECT 2.800 3487.020 2917.930 3487.700 ;
        RECT 2.800 3485.700 2917.200 3487.020 ;
        RECT 2.400 3485.020 2917.200 3485.700 ;
        RECT 2.400 3422.420 2917.930 3485.020 ;
        RECT 2.800 3420.420 2917.930 3422.420 ;
        RECT 2.400 3420.380 2917.930 3420.420 ;
        RECT 2.400 3418.380 2917.200 3420.380 ;
        RECT 2.400 3357.140 2917.930 3418.380 ;
        RECT 2.800 3355.140 2917.930 3357.140 ;
        RECT 2.400 3354.420 2917.930 3355.140 ;
        RECT 2.400 3352.420 2917.200 3354.420 ;
        RECT 2.400 3291.860 2917.930 3352.420 ;
        RECT 2.800 3289.860 2917.930 3291.860 ;
        RECT 2.400 3287.780 2917.930 3289.860 ;
        RECT 2.400 3285.780 2917.200 3287.780 ;
        RECT 2.400 3226.580 2917.930 3285.780 ;
        RECT 2.800 3224.580 2917.930 3226.580 ;
        RECT 2.400 3221.140 2917.930 3224.580 ;
        RECT 2.400 3219.140 2917.200 3221.140 ;
        RECT 2.400 3161.300 2917.930 3219.140 ;
        RECT 2.800 3159.300 2917.930 3161.300 ;
        RECT 2.400 3155.180 2917.930 3159.300 ;
        RECT 2.400 3153.180 2917.200 3155.180 ;
        RECT 2.400 3096.700 2917.930 3153.180 ;
        RECT 2.800 3094.700 2917.930 3096.700 ;
        RECT 2.400 3088.540 2917.930 3094.700 ;
        RECT 2.400 3086.540 2917.200 3088.540 ;
        RECT 2.400 3031.420 2917.930 3086.540 ;
        RECT 2.800 3029.420 2917.930 3031.420 ;
        RECT 2.400 3021.900 2917.930 3029.420 ;
        RECT 2.400 3019.900 2917.200 3021.900 ;
        RECT 2.400 2966.140 2917.930 3019.900 ;
        RECT 2.800 2964.140 2917.930 2966.140 ;
        RECT 2.400 2955.940 2917.930 2964.140 ;
        RECT 2.400 2953.940 2917.200 2955.940 ;
        RECT 2.400 2900.860 2917.930 2953.940 ;
        RECT 2.800 2898.860 2917.930 2900.860 ;
        RECT 2.400 2889.300 2917.930 2898.860 ;
        RECT 2.400 2887.300 2917.200 2889.300 ;
        RECT 2.400 2835.580 2917.930 2887.300 ;
        RECT 2.800 2833.580 2917.930 2835.580 ;
        RECT 2.400 2822.660 2917.930 2833.580 ;
        RECT 2.400 2820.660 2917.200 2822.660 ;
        RECT 2.400 2770.300 2917.930 2820.660 ;
        RECT 2.800 2768.300 2917.930 2770.300 ;
        RECT 2.400 2756.700 2917.930 2768.300 ;
        RECT 2.400 2754.700 2917.200 2756.700 ;
        RECT 2.400 2705.020 2917.930 2754.700 ;
        RECT 2.800 2703.020 2917.930 2705.020 ;
        RECT 2.400 2690.060 2917.930 2703.020 ;
        RECT 2.400 2688.060 2917.200 2690.060 ;
        RECT 2.400 2640.420 2917.930 2688.060 ;
        RECT 2.800 2638.420 2917.930 2640.420 ;
        RECT 2.400 2623.420 2917.930 2638.420 ;
        RECT 2.400 2621.420 2917.200 2623.420 ;
        RECT 2.400 2575.140 2917.930 2621.420 ;
        RECT 2.800 2573.140 2917.930 2575.140 ;
        RECT 2.400 2557.460 2917.930 2573.140 ;
        RECT 2.400 2555.460 2917.200 2557.460 ;
        RECT 2.400 2509.860 2917.930 2555.460 ;
        RECT 2.800 2507.860 2917.930 2509.860 ;
        RECT 2.400 2490.820 2917.930 2507.860 ;
        RECT 2.400 2488.820 2917.200 2490.820 ;
        RECT 2.400 2444.580 2917.930 2488.820 ;
        RECT 2.800 2442.580 2917.930 2444.580 ;
        RECT 2.400 2424.180 2917.930 2442.580 ;
        RECT 2.400 2422.180 2917.200 2424.180 ;
        RECT 2.400 2379.300 2917.930 2422.180 ;
        RECT 2.800 2377.300 2917.930 2379.300 ;
        RECT 2.400 2358.220 2917.930 2377.300 ;
        RECT 2.400 2356.220 2917.200 2358.220 ;
        RECT 2.400 2314.020 2917.930 2356.220 ;
        RECT 2.800 2312.020 2917.930 2314.020 ;
        RECT 2.400 2291.580 2917.930 2312.020 ;
        RECT 2.400 2289.580 2917.200 2291.580 ;
        RECT 2.400 2248.740 2917.930 2289.580 ;
        RECT 2.800 2246.740 2917.930 2248.740 ;
        RECT 2.400 2224.940 2917.930 2246.740 ;
        RECT 2.400 2222.940 2917.200 2224.940 ;
        RECT 2.400 2184.140 2917.930 2222.940 ;
        RECT 2.800 2182.140 2917.930 2184.140 ;
        RECT 2.400 2158.980 2917.930 2182.140 ;
        RECT 2.400 2156.980 2917.200 2158.980 ;
        RECT 2.400 2118.860 2917.930 2156.980 ;
        RECT 2.800 2116.860 2917.930 2118.860 ;
        RECT 2.400 2092.340 2917.930 2116.860 ;
        RECT 2.400 2090.340 2917.200 2092.340 ;
        RECT 2.400 2053.580 2917.930 2090.340 ;
        RECT 2.800 2051.580 2917.930 2053.580 ;
        RECT 2.400 2025.700 2917.930 2051.580 ;
        RECT 2.400 2023.700 2917.200 2025.700 ;
        RECT 2.400 1988.300 2917.930 2023.700 ;
        RECT 2.800 1986.300 2917.930 1988.300 ;
        RECT 2.400 1959.740 2917.930 1986.300 ;
        RECT 2.400 1957.740 2917.200 1959.740 ;
        RECT 2.400 1923.020 2917.930 1957.740 ;
        RECT 2.800 1921.020 2917.930 1923.020 ;
        RECT 2.400 1893.100 2917.930 1921.020 ;
        RECT 2.400 1891.100 2917.200 1893.100 ;
        RECT 2.400 1857.740 2917.930 1891.100 ;
        RECT 2.800 1855.740 2917.930 1857.740 ;
        RECT 2.400 1826.460 2917.930 1855.740 ;
        RECT 2.400 1824.460 2917.200 1826.460 ;
        RECT 2.400 1793.140 2917.930 1824.460 ;
        RECT 2.800 1791.140 2917.930 1793.140 ;
        RECT 2.400 1760.500 2917.930 1791.140 ;
        RECT 2.400 1758.500 2917.200 1760.500 ;
        RECT 2.400 1727.860 2917.930 1758.500 ;
        RECT 2.800 1725.860 2917.930 1727.860 ;
        RECT 2.400 1693.860 2917.930 1725.860 ;
        RECT 2.400 1691.860 2917.200 1693.860 ;
        RECT 2.400 1662.580 2917.930 1691.860 ;
        RECT 2.800 1660.580 2917.930 1662.580 ;
        RECT 2.400 1627.220 2917.930 1660.580 ;
        RECT 2.400 1625.220 2917.200 1627.220 ;
        RECT 2.400 1597.300 2917.930 1625.220 ;
        RECT 2.800 1595.300 2917.930 1597.300 ;
        RECT 2.400 1561.260 2917.930 1595.300 ;
        RECT 2.400 1559.260 2917.200 1561.260 ;
        RECT 2.400 1532.020 2917.930 1559.260 ;
        RECT 2.800 1530.020 2917.930 1532.020 ;
        RECT 2.400 1494.620 2917.930 1530.020 ;
        RECT 2.400 1492.620 2917.200 1494.620 ;
        RECT 2.400 1466.740 2917.930 1492.620 ;
        RECT 2.800 1464.740 2917.930 1466.740 ;
        RECT 2.400 1427.980 2917.930 1464.740 ;
        RECT 2.400 1425.980 2917.200 1427.980 ;
        RECT 2.400 1401.460 2917.930 1425.980 ;
        RECT 2.800 1399.460 2917.930 1401.460 ;
        RECT 2.400 1362.020 2917.930 1399.460 ;
        RECT 2.400 1360.020 2917.200 1362.020 ;
        RECT 2.400 1336.860 2917.930 1360.020 ;
        RECT 2.800 1334.860 2917.930 1336.860 ;
        RECT 2.400 1295.380 2917.930 1334.860 ;
        RECT 2.400 1293.380 2917.200 1295.380 ;
        RECT 2.400 1271.580 2917.930 1293.380 ;
        RECT 2.800 1269.580 2917.930 1271.580 ;
        RECT 2.400 1228.740 2917.930 1269.580 ;
        RECT 2.400 1226.740 2917.200 1228.740 ;
        RECT 2.400 1206.300 2917.930 1226.740 ;
        RECT 2.800 1204.300 2917.930 1206.300 ;
        RECT 2.400 1162.780 2917.930 1204.300 ;
        RECT 2.400 1160.780 2917.200 1162.780 ;
        RECT 2.400 1141.020 2917.930 1160.780 ;
        RECT 2.800 1139.020 2917.930 1141.020 ;
        RECT 2.400 1096.140 2917.930 1139.020 ;
        RECT 2.400 1094.140 2917.200 1096.140 ;
        RECT 2.400 1075.740 2917.930 1094.140 ;
        RECT 2.800 1073.740 2917.930 1075.740 ;
        RECT 2.400 1029.500 2917.930 1073.740 ;
        RECT 2.400 1027.500 2917.200 1029.500 ;
        RECT 2.400 1010.460 2917.930 1027.500 ;
        RECT 2.800 1008.460 2917.930 1010.460 ;
        RECT 2.400 963.540 2917.930 1008.460 ;
        RECT 2.400 961.540 2917.200 963.540 ;
        RECT 2.400 945.180 2917.930 961.540 ;
        RECT 2.800 943.180 2917.930 945.180 ;
        RECT 2.400 896.900 2917.930 943.180 ;
        RECT 2.400 894.900 2917.200 896.900 ;
        RECT 2.400 880.580 2917.930 894.900 ;
        RECT 2.800 878.580 2917.930 880.580 ;
        RECT 2.400 830.260 2917.930 878.580 ;
        RECT 2.400 828.260 2917.200 830.260 ;
        RECT 2.400 815.300 2917.930 828.260 ;
        RECT 2.800 813.300 2917.930 815.300 ;
        RECT 2.400 764.300 2917.930 813.300 ;
        RECT 2.400 762.300 2917.200 764.300 ;
        RECT 2.400 750.020 2917.930 762.300 ;
        RECT 2.800 748.020 2917.930 750.020 ;
        RECT 2.400 697.660 2917.930 748.020 ;
        RECT 2.400 695.660 2917.200 697.660 ;
        RECT 2.400 684.740 2917.930 695.660 ;
        RECT 2.800 682.740 2917.930 684.740 ;
        RECT 2.400 631.020 2917.930 682.740 ;
        RECT 2.400 629.020 2917.200 631.020 ;
        RECT 2.400 619.460 2917.930 629.020 ;
        RECT 2.800 617.460 2917.930 619.460 ;
        RECT 2.400 565.060 2917.930 617.460 ;
        RECT 2.400 563.060 2917.200 565.060 ;
        RECT 2.400 554.180 2917.930 563.060 ;
        RECT 2.800 552.180 2917.930 554.180 ;
        RECT 2.400 498.420 2917.930 552.180 ;
        RECT 2.400 496.420 2917.200 498.420 ;
        RECT 2.400 488.900 2917.930 496.420 ;
        RECT 2.800 486.900 2917.930 488.900 ;
        RECT 2.400 431.780 2917.930 486.900 ;
        RECT 2.400 429.780 2917.200 431.780 ;
        RECT 2.400 424.300 2917.930 429.780 ;
        RECT 2.800 422.300 2917.930 424.300 ;
        RECT 2.400 365.820 2917.930 422.300 ;
        RECT 2.400 363.820 2917.200 365.820 ;
        RECT 2.400 359.020 2917.930 363.820 ;
        RECT 2.800 357.020 2917.930 359.020 ;
        RECT 2.400 299.180 2917.930 357.020 ;
        RECT 2.400 297.180 2917.200 299.180 ;
        RECT 2.400 293.740 2917.930 297.180 ;
        RECT 2.800 291.740 2917.930 293.740 ;
        RECT 2.400 232.540 2917.930 291.740 ;
        RECT 2.400 230.540 2917.200 232.540 ;
        RECT 2.400 228.460 2917.930 230.540 ;
        RECT 2.800 226.460 2917.930 228.460 ;
        RECT 2.400 166.580 2917.930 226.460 ;
        RECT 2.400 164.580 2917.200 166.580 ;
        RECT 2.400 163.180 2917.930 164.580 ;
        RECT 2.800 161.180 2917.930 163.180 ;
        RECT 2.400 99.940 2917.930 161.180 ;
        RECT 2.400 97.940 2917.200 99.940 ;
        RECT 2.400 97.900 2917.930 97.940 ;
        RECT 2.800 95.900 2917.930 97.900 ;
        RECT 2.400 57.975 2917.930 95.900 ;
      LAYER met4 ;
        RECT 285.495 3226.140 288.570 3501.825 ;
        RECT 292.470 3226.140 307.170 3501.825 ;
        RECT 311.070 3226.140 325.770 3501.825 ;
        RECT 329.670 3226.140 344.370 3501.825 ;
        RECT 348.270 3226.140 358.570 3501.825 ;
        RECT 362.470 3226.140 377.170 3501.825 ;
        RECT 381.070 3226.140 395.770 3501.825 ;
        RECT 399.670 3226.140 414.370 3501.825 ;
        RECT 418.270 3226.140 428.570 3501.825 ;
        RECT 432.470 3226.140 447.170 3501.825 ;
        RECT 451.070 3226.140 465.770 3501.825 ;
        RECT 469.670 3226.140 484.370 3501.825 ;
        RECT 488.270 3226.140 498.570 3501.825 ;
        RECT 502.470 3226.140 517.170 3501.825 ;
        RECT 521.070 3226.140 535.770 3501.825 ;
        RECT 539.670 3226.140 554.370 3501.825 ;
        RECT 558.270 3226.140 568.570 3501.825 ;
        RECT 572.470 3226.140 587.170 3501.825 ;
        RECT 591.070 3226.140 605.770 3501.825 ;
        RECT 609.670 3226.140 624.370 3501.825 ;
        RECT 628.270 3226.140 638.570 3501.825 ;
        RECT 642.470 3226.140 657.170 3501.825 ;
        RECT 661.070 3226.140 675.770 3501.825 ;
        RECT 679.670 3226.140 694.370 3501.825 ;
        RECT 698.270 3226.140 708.570 3501.825 ;
        RECT 712.470 3226.140 727.170 3501.825 ;
        RECT 731.070 3226.140 745.770 3501.825 ;
        RECT 749.670 3226.140 764.370 3501.825 ;
        RECT 768.270 3226.140 778.570 3501.825 ;
        RECT 782.470 3226.140 797.170 3501.825 ;
        RECT 801.070 3226.140 815.770 3501.825 ;
        RECT 819.670 3226.140 834.370 3501.825 ;
        RECT 838.270 3226.140 848.570 3501.825 ;
        RECT 852.470 3226.140 867.170 3501.825 ;
        RECT 871.070 3226.140 885.770 3501.825 ;
        RECT 889.670 3226.140 904.370 3501.825 ;
        RECT 908.270 3226.140 918.570 3501.825 ;
        RECT 922.470 3226.140 937.170 3501.825 ;
        RECT 941.070 3226.140 955.770 3501.825 ;
        RECT 959.670 3226.140 974.370 3501.825 ;
        RECT 978.270 3226.140 988.570 3501.825 ;
        RECT 992.470 3226.140 1007.170 3501.825 ;
        RECT 285.495 2790.400 1007.170 3226.140 ;
        RECT 285.495 2691.140 288.570 2790.400 ;
        RECT 292.470 2691.140 307.170 2790.400 ;
        RECT 311.070 2691.140 325.770 2790.400 ;
        RECT 329.670 2691.140 344.370 2790.400 ;
        RECT 348.270 2691.140 358.570 2790.400 ;
        RECT 362.470 2691.140 377.170 2790.400 ;
        RECT 381.070 2691.140 395.770 2790.400 ;
        RECT 399.670 2691.140 414.370 2790.400 ;
        RECT 418.270 2691.140 428.570 2790.400 ;
        RECT 432.470 2691.140 447.170 2790.400 ;
        RECT 451.070 2691.140 465.770 2790.400 ;
        RECT 469.670 2691.140 484.370 2790.400 ;
        RECT 488.270 2691.140 498.570 2790.400 ;
        RECT 502.470 2691.140 517.170 2790.400 ;
        RECT 521.070 2691.140 535.770 2790.400 ;
        RECT 539.670 2691.140 554.370 2790.400 ;
        RECT 558.270 2691.140 568.570 2790.400 ;
        RECT 572.470 2691.140 587.170 2790.400 ;
        RECT 591.070 2691.140 605.770 2790.400 ;
        RECT 609.670 2691.140 624.370 2790.400 ;
        RECT 628.270 2691.140 638.570 2790.400 ;
        RECT 642.470 2691.140 657.170 2790.400 ;
        RECT 661.070 2691.140 675.770 2790.400 ;
        RECT 679.670 2691.140 694.370 2790.400 ;
        RECT 698.270 2691.140 708.570 2790.400 ;
        RECT 712.470 2691.140 727.170 2790.400 ;
        RECT 731.070 2691.140 745.770 2790.400 ;
        RECT 749.670 2691.140 764.370 2790.400 ;
        RECT 768.270 2691.140 778.570 2790.400 ;
        RECT 782.470 2691.140 797.170 2790.400 ;
        RECT 801.070 2691.140 815.770 2790.400 ;
        RECT 819.670 2691.140 834.370 2790.400 ;
        RECT 838.270 2691.140 848.570 2790.400 ;
        RECT 852.470 2691.140 867.170 2790.400 ;
        RECT 871.070 2691.140 885.770 2790.400 ;
        RECT 889.670 2691.140 904.370 2790.400 ;
        RECT 908.270 2691.140 918.570 2790.400 ;
        RECT 922.470 2691.140 937.170 2790.400 ;
        RECT 941.070 2691.140 955.770 2790.400 ;
        RECT 959.670 2691.140 974.370 2790.400 ;
        RECT 978.270 2691.140 988.570 2790.400 ;
        RECT 992.470 2691.140 1007.170 2790.400 ;
        RECT 285.495 2255.400 1007.170 2691.140 ;
        RECT 285.495 2134.765 288.570 2255.400 ;
        RECT 292.470 2134.765 307.170 2255.400 ;
        RECT 311.070 2134.765 325.770 2255.400 ;
        RECT 329.670 2134.765 344.370 2255.400 ;
        RECT 348.270 2134.765 358.570 2255.400 ;
        RECT 362.470 2134.765 377.170 2255.400 ;
        RECT 381.070 2134.765 395.770 2255.400 ;
        RECT 399.670 2134.765 414.370 2255.400 ;
        RECT 418.270 2134.765 428.570 2255.400 ;
        RECT 432.470 2134.765 447.170 2255.400 ;
        RECT 451.070 2134.765 465.770 2255.400 ;
        RECT 469.670 2134.765 484.370 2255.400 ;
        RECT 488.270 2134.765 498.570 2255.400 ;
        RECT 502.470 2134.765 517.170 2255.400 ;
        RECT 521.070 2134.765 535.770 2255.400 ;
        RECT 539.670 2134.765 554.370 2255.400 ;
        RECT 558.270 2134.765 568.570 2255.400 ;
        RECT 572.470 2134.765 587.170 2255.400 ;
        RECT 591.070 2134.765 605.770 2255.400 ;
        RECT 609.670 2134.765 624.370 2255.400 ;
        RECT 628.270 2134.765 638.570 2255.400 ;
        RECT 642.470 2134.765 657.170 2255.400 ;
        RECT 661.070 2134.765 675.770 2255.400 ;
        RECT 679.670 2134.765 694.370 2255.400 ;
        RECT 698.270 2134.765 708.570 2255.400 ;
        RECT 712.470 2134.765 727.170 2255.400 ;
        RECT 731.070 2134.765 745.770 2255.400 ;
        RECT 749.670 2134.765 764.370 2255.400 ;
        RECT 768.270 2134.765 778.570 2255.400 ;
        RECT 782.470 2134.765 797.170 2255.400 ;
        RECT 801.070 2134.765 815.770 2255.400 ;
        RECT 819.670 2134.765 834.370 2255.400 ;
        RECT 838.270 2134.765 848.570 2255.400 ;
        RECT 852.470 2134.765 867.170 2255.400 ;
        RECT 285.495 1560.400 867.170 2134.765 ;
        RECT 285.495 1261.140 288.570 1560.400 ;
        RECT 292.470 1261.140 307.170 1560.400 ;
        RECT 311.070 1261.140 325.770 1560.400 ;
        RECT 329.670 1261.140 344.370 1560.400 ;
        RECT 348.270 1261.140 358.570 1560.400 ;
        RECT 362.470 1261.140 377.170 1560.400 ;
        RECT 381.070 1261.140 395.770 1560.400 ;
        RECT 399.670 1261.140 414.370 1560.400 ;
        RECT 418.270 1261.140 428.570 1560.400 ;
        RECT 432.470 1261.140 447.170 1560.400 ;
        RECT 451.070 1261.140 465.770 1560.400 ;
        RECT 469.670 1261.140 484.370 1560.400 ;
        RECT 488.270 1261.140 498.570 1560.400 ;
        RECT 502.470 1261.140 517.170 1560.400 ;
        RECT 521.070 1261.140 535.770 1560.400 ;
        RECT 539.670 1261.140 554.370 1560.400 ;
        RECT 558.270 1261.140 568.570 1560.400 ;
        RECT 572.470 1261.140 587.170 1560.400 ;
        RECT 591.070 1261.140 605.770 1560.400 ;
        RECT 609.670 1261.140 624.370 1560.400 ;
        RECT 628.270 1261.140 638.570 1560.400 ;
        RECT 642.470 1261.140 657.170 1560.400 ;
        RECT 661.070 1261.140 675.770 1560.400 ;
        RECT 679.670 1261.140 694.370 1560.400 ;
        RECT 698.270 1261.140 708.570 1560.400 ;
        RECT 712.470 1261.140 727.170 1560.400 ;
        RECT 731.070 1261.140 745.770 1560.400 ;
        RECT 749.670 1261.140 764.370 1560.400 ;
        RECT 768.270 1261.140 778.570 1560.400 ;
        RECT 782.470 1261.140 797.170 1560.400 ;
        RECT 801.070 1261.140 815.770 1560.400 ;
        RECT 819.670 1261.140 834.370 1560.400 ;
        RECT 838.270 1261.140 848.570 1560.400 ;
        RECT 852.470 1261.140 867.170 1560.400 ;
        RECT 871.070 1261.140 885.770 2255.400 ;
        RECT 889.670 1261.140 904.370 2255.400 ;
        RECT 908.270 1261.140 918.570 2255.400 ;
        RECT 922.470 1261.140 937.170 2255.400 ;
        RECT 941.070 1261.140 955.770 2255.400 ;
        RECT 959.670 1261.140 974.370 2255.400 ;
        RECT 978.270 2129.600 988.570 2255.400 ;
        RECT 992.470 2129.600 1007.170 2255.400 ;
        RECT 1011.070 2129.600 1025.770 3501.825 ;
        RECT 1029.670 2129.600 1044.370 3501.825 ;
        RECT 1048.270 2129.600 1058.570 3501.825 ;
        RECT 1062.470 2129.600 1077.170 3501.825 ;
        RECT 1081.070 3226.140 1095.770 3501.825 ;
        RECT 1099.670 3226.140 1114.370 3501.825 ;
        RECT 1118.270 3226.140 1128.570 3501.825 ;
        RECT 1132.470 3226.140 1147.170 3501.825 ;
        RECT 1151.070 3226.140 1165.770 3501.825 ;
        RECT 1169.670 3226.140 1184.370 3501.825 ;
        RECT 1188.270 3226.140 1198.570 3501.825 ;
        RECT 1202.470 3226.140 1217.170 3501.825 ;
        RECT 1221.070 3226.140 1235.770 3501.825 ;
        RECT 1239.670 3226.140 1254.370 3501.825 ;
        RECT 1258.270 3226.140 1268.570 3501.825 ;
        RECT 1272.470 3226.140 1287.170 3501.825 ;
        RECT 1291.070 3226.140 1305.770 3501.825 ;
        RECT 1309.670 3226.140 1324.370 3501.825 ;
        RECT 1328.270 3226.140 1338.570 3501.825 ;
        RECT 1342.470 3226.140 1357.170 3501.825 ;
        RECT 1361.070 3226.140 1375.770 3501.825 ;
        RECT 1379.670 3226.140 1394.370 3501.825 ;
        RECT 1398.270 3226.140 1408.570 3501.825 ;
        RECT 1412.470 3226.140 1427.170 3501.825 ;
        RECT 1431.070 3226.140 1445.770 3501.825 ;
        RECT 1449.670 3226.140 1464.370 3501.825 ;
        RECT 1468.270 3226.140 1478.570 3501.825 ;
        RECT 1482.470 3226.140 1497.170 3501.825 ;
        RECT 1501.070 3226.140 1515.770 3501.825 ;
        RECT 1519.670 3226.140 1534.370 3501.825 ;
        RECT 1538.270 3226.140 1548.570 3501.825 ;
        RECT 1552.470 3226.140 1567.170 3501.825 ;
        RECT 1571.070 3226.140 1585.770 3501.825 ;
        RECT 1589.670 3226.140 1604.370 3501.825 ;
        RECT 1608.270 3226.140 1618.570 3501.825 ;
        RECT 1622.470 3226.140 1637.170 3501.825 ;
        RECT 1641.070 3226.140 1655.770 3501.825 ;
        RECT 1659.670 3226.140 1674.370 3501.825 ;
        RECT 1678.270 3226.140 1688.570 3501.825 ;
        RECT 1692.470 3226.140 1707.170 3501.825 ;
        RECT 1711.070 3226.140 1725.770 3501.825 ;
        RECT 1729.670 3226.140 1744.370 3501.825 ;
        RECT 1748.270 3226.140 1758.570 3501.825 ;
        RECT 1762.470 3226.140 1777.170 3501.825 ;
        RECT 1781.070 3226.140 1795.770 3501.825 ;
        RECT 1081.070 2790.400 1795.770 3226.140 ;
        RECT 1081.070 2691.140 1095.770 2790.400 ;
        RECT 1099.670 2691.140 1114.370 2790.400 ;
        RECT 1118.270 2691.140 1128.570 2790.400 ;
        RECT 1132.470 2691.140 1147.170 2790.400 ;
        RECT 1151.070 2691.140 1165.770 2790.400 ;
        RECT 1169.670 2691.140 1184.370 2790.400 ;
        RECT 1188.270 2691.140 1198.570 2790.400 ;
        RECT 1202.470 2691.140 1217.170 2790.400 ;
        RECT 1221.070 2691.140 1235.770 2790.400 ;
        RECT 1239.670 2691.140 1254.370 2790.400 ;
        RECT 1258.270 2691.140 1268.570 2790.400 ;
        RECT 1272.470 2691.140 1287.170 2790.400 ;
        RECT 1291.070 2691.140 1305.770 2790.400 ;
        RECT 1309.670 2691.140 1324.370 2790.400 ;
        RECT 1328.270 2691.140 1338.570 2790.400 ;
        RECT 1342.470 2691.140 1357.170 2790.400 ;
        RECT 1361.070 2691.140 1375.770 2790.400 ;
        RECT 1379.670 2691.140 1394.370 2790.400 ;
        RECT 1398.270 2691.140 1408.570 2790.400 ;
        RECT 1412.470 2691.140 1427.170 2790.400 ;
        RECT 1431.070 2691.140 1445.770 2790.400 ;
        RECT 1449.670 2691.140 1464.370 2790.400 ;
        RECT 1468.270 2691.140 1478.570 2790.400 ;
        RECT 1482.470 2691.140 1497.170 2790.400 ;
        RECT 1501.070 2691.140 1515.770 2790.400 ;
        RECT 1519.670 2691.140 1534.370 2790.400 ;
        RECT 1538.270 2691.140 1548.570 2790.400 ;
        RECT 1552.470 2691.140 1567.170 2790.400 ;
        RECT 1571.070 2691.140 1585.770 2790.400 ;
        RECT 1589.670 2691.140 1604.370 2790.400 ;
        RECT 1608.270 2691.140 1618.570 2790.400 ;
        RECT 1622.470 2691.140 1637.170 2790.400 ;
        RECT 1641.070 2691.140 1655.770 2790.400 ;
        RECT 1659.670 2691.140 1674.370 2790.400 ;
        RECT 1678.270 2691.140 1688.570 2790.400 ;
        RECT 1692.470 2691.140 1707.170 2790.400 ;
        RECT 1711.070 2691.140 1725.770 2790.400 ;
        RECT 1729.670 2691.140 1744.370 2790.400 ;
        RECT 1748.270 2691.140 1758.570 2790.400 ;
        RECT 1762.470 2691.140 1777.170 2790.400 ;
        RECT 1781.070 2691.140 1795.770 2790.400 ;
        RECT 1081.070 2255.400 1795.770 2691.140 ;
        RECT 1081.070 2129.600 1095.770 2255.400 ;
        RECT 1099.670 2129.600 1114.370 2255.400 ;
        RECT 1118.270 2129.600 1128.570 2255.400 ;
        RECT 1132.470 2129.600 1147.170 2255.400 ;
        RECT 1151.070 2129.600 1165.770 2255.400 ;
        RECT 1169.670 2129.600 1184.370 2255.400 ;
        RECT 1188.270 2129.600 1198.570 2255.400 ;
        RECT 1202.470 2129.600 1217.170 2255.400 ;
        RECT 1221.070 2129.600 1235.770 2255.400 ;
        RECT 1239.670 2129.600 1254.370 2255.400 ;
        RECT 1258.270 2129.600 1268.570 2255.400 ;
        RECT 1272.470 2129.600 1287.170 2255.400 ;
        RECT 1291.070 2129.600 1305.770 2255.400 ;
        RECT 1309.670 2129.600 1324.370 2255.400 ;
        RECT 1328.270 2129.600 1338.570 2255.400 ;
        RECT 1342.470 2129.600 1357.170 2255.400 ;
        RECT 1361.070 2129.600 1375.770 2255.400 ;
        RECT 1379.670 2129.600 1394.370 2255.400 ;
        RECT 1398.270 2129.600 1408.570 2255.400 ;
        RECT 1412.470 2129.600 1427.170 2255.400 ;
        RECT 1431.070 2129.600 1445.770 2255.400 ;
        RECT 1449.670 2129.600 1464.370 2255.400 ;
        RECT 1468.270 2129.600 1478.570 2255.400 ;
        RECT 1482.470 2129.600 1497.170 2255.400 ;
        RECT 1501.070 2129.600 1515.770 2255.400 ;
        RECT 1519.670 2129.600 1534.370 2255.400 ;
        RECT 1538.270 2129.600 1548.570 2255.400 ;
        RECT 1552.470 2129.600 1567.170 2255.400 ;
        RECT 1571.070 2129.600 1585.770 2255.400 ;
        RECT 1589.670 2129.600 1604.370 2255.400 ;
        RECT 1608.270 2129.600 1618.570 2255.400 ;
        RECT 978.270 1375.400 1618.570 2129.600 ;
        RECT 978.270 1261.140 988.570 1375.400 ;
        RECT 992.470 1261.140 1007.170 1375.400 ;
        RECT 285.495 825.400 1007.170 1261.140 ;
        RECT 285.495 726.140 288.570 825.400 ;
        RECT 292.470 726.140 307.170 825.400 ;
        RECT 311.070 726.140 325.770 825.400 ;
        RECT 329.670 726.140 344.370 825.400 ;
        RECT 348.270 726.140 358.570 825.400 ;
        RECT 362.470 726.140 377.170 825.400 ;
        RECT 381.070 726.140 395.770 825.400 ;
        RECT 399.670 726.140 414.370 825.400 ;
        RECT 418.270 726.140 428.570 825.400 ;
        RECT 432.470 726.140 447.170 825.400 ;
        RECT 451.070 726.140 465.770 825.400 ;
        RECT 469.670 726.140 484.370 825.400 ;
        RECT 488.270 726.140 498.570 825.400 ;
        RECT 502.470 726.140 517.170 825.400 ;
        RECT 521.070 726.140 535.770 825.400 ;
        RECT 539.670 726.140 554.370 825.400 ;
        RECT 558.270 726.140 568.570 825.400 ;
        RECT 572.470 726.140 587.170 825.400 ;
        RECT 591.070 726.140 605.770 825.400 ;
        RECT 609.670 726.140 624.370 825.400 ;
        RECT 628.270 726.140 638.570 825.400 ;
        RECT 642.470 726.140 657.170 825.400 ;
        RECT 661.070 726.140 675.770 825.400 ;
        RECT 679.670 726.140 694.370 825.400 ;
        RECT 698.270 726.140 708.570 825.400 ;
        RECT 712.470 726.140 727.170 825.400 ;
        RECT 731.070 726.140 745.770 825.400 ;
        RECT 749.670 726.140 764.370 825.400 ;
        RECT 768.270 726.140 778.570 825.400 ;
        RECT 782.470 726.140 797.170 825.400 ;
        RECT 801.070 726.140 815.770 825.400 ;
        RECT 819.670 726.140 834.370 825.400 ;
        RECT 838.270 726.140 848.570 825.400 ;
        RECT 852.470 726.140 867.170 825.400 ;
        RECT 871.070 726.140 885.770 825.400 ;
        RECT 889.670 726.140 904.370 825.400 ;
        RECT 908.270 726.140 918.570 825.400 ;
        RECT 922.470 726.140 937.170 825.400 ;
        RECT 941.070 726.140 955.770 825.400 ;
        RECT 959.670 726.140 974.370 825.400 ;
        RECT 978.270 726.140 988.570 825.400 ;
        RECT 992.470 726.140 1007.170 825.400 ;
        RECT 285.495 290.400 1007.170 726.140 ;
        RECT 285.495 57.975 288.570 290.400 ;
        RECT 292.470 57.975 307.170 290.400 ;
        RECT 311.070 57.975 325.770 290.400 ;
        RECT 329.670 57.975 344.370 290.400 ;
        RECT 348.270 57.975 358.570 290.400 ;
        RECT 362.470 57.975 377.170 290.400 ;
        RECT 381.070 57.975 395.770 290.400 ;
        RECT 399.670 57.975 414.370 290.400 ;
        RECT 418.270 57.975 428.570 290.400 ;
        RECT 432.470 57.975 447.170 290.400 ;
        RECT 451.070 57.975 465.770 290.400 ;
        RECT 469.670 57.975 484.370 290.400 ;
        RECT 488.270 57.975 498.570 290.400 ;
        RECT 502.470 57.975 517.170 290.400 ;
        RECT 521.070 57.975 535.770 290.400 ;
        RECT 539.670 57.975 554.370 290.400 ;
        RECT 558.270 57.975 568.570 290.400 ;
        RECT 572.470 57.975 587.170 290.400 ;
        RECT 591.070 57.975 605.770 290.400 ;
        RECT 609.670 57.975 624.370 290.400 ;
        RECT 628.270 57.975 638.570 290.400 ;
        RECT 642.470 57.975 657.170 290.400 ;
        RECT 661.070 57.975 675.770 290.400 ;
        RECT 679.670 57.975 694.370 290.400 ;
        RECT 698.270 57.975 708.570 290.400 ;
        RECT 712.470 57.975 727.170 290.400 ;
        RECT 731.070 57.975 745.770 290.400 ;
        RECT 749.670 57.975 764.370 290.400 ;
        RECT 768.270 57.975 778.570 290.400 ;
        RECT 782.470 57.975 797.170 290.400 ;
        RECT 801.070 57.975 815.770 290.400 ;
        RECT 819.670 57.975 834.370 290.400 ;
        RECT 838.270 57.975 848.570 290.400 ;
        RECT 852.470 57.975 867.170 290.400 ;
        RECT 871.070 57.975 885.770 290.400 ;
        RECT 889.670 57.975 904.370 290.400 ;
        RECT 908.270 57.975 918.570 290.400 ;
        RECT 922.470 57.975 937.170 290.400 ;
        RECT 941.070 57.975 955.770 290.400 ;
        RECT 959.670 57.975 974.370 290.400 ;
        RECT 978.270 57.975 988.570 290.400 ;
        RECT 992.470 57.975 1007.170 290.400 ;
        RECT 1011.070 57.975 1025.770 1375.400 ;
        RECT 1029.670 57.975 1044.370 1375.400 ;
        RECT 1048.270 57.975 1058.570 1375.400 ;
        RECT 1062.470 57.975 1077.170 1375.400 ;
        RECT 1081.070 1261.140 1095.770 1375.400 ;
        RECT 1099.670 1261.140 1114.370 1375.400 ;
        RECT 1118.270 1261.140 1128.570 1375.400 ;
        RECT 1132.470 1261.140 1147.170 1375.400 ;
        RECT 1151.070 1261.140 1165.770 1375.400 ;
        RECT 1169.670 1261.140 1184.370 1375.400 ;
        RECT 1188.270 1261.140 1198.570 1375.400 ;
        RECT 1202.470 1261.140 1217.170 1375.400 ;
        RECT 1221.070 1261.140 1235.770 1375.400 ;
        RECT 1239.670 1261.140 1254.370 1375.400 ;
        RECT 1258.270 1261.140 1268.570 1375.400 ;
        RECT 1272.470 1261.140 1287.170 1375.400 ;
        RECT 1291.070 1261.140 1305.770 1375.400 ;
        RECT 1309.670 1261.140 1324.370 1375.400 ;
        RECT 1328.270 1261.140 1338.570 1375.400 ;
        RECT 1342.470 1261.140 1357.170 1375.400 ;
        RECT 1361.070 1261.140 1375.770 1375.400 ;
        RECT 1379.670 1261.140 1394.370 1375.400 ;
        RECT 1398.270 1261.140 1408.570 1375.400 ;
        RECT 1412.470 1261.140 1427.170 1375.400 ;
        RECT 1431.070 1261.140 1445.770 1375.400 ;
        RECT 1449.670 1261.140 1464.370 1375.400 ;
        RECT 1468.270 1261.140 1478.570 1375.400 ;
        RECT 1482.470 1261.140 1497.170 1375.400 ;
        RECT 1501.070 1261.140 1515.770 1375.400 ;
        RECT 1519.670 1261.140 1534.370 1375.400 ;
        RECT 1538.270 1261.140 1548.570 1375.400 ;
        RECT 1552.470 1261.140 1567.170 1375.400 ;
        RECT 1571.070 1261.140 1585.770 1375.400 ;
        RECT 1589.670 1261.140 1604.370 1375.400 ;
        RECT 1608.270 1261.140 1618.570 1375.400 ;
        RECT 1622.470 1261.140 1637.170 2255.400 ;
        RECT 1641.070 1261.140 1655.770 2255.400 ;
        RECT 1659.670 1261.140 1674.370 2255.400 ;
        RECT 1678.270 1261.140 1688.570 2255.400 ;
        RECT 1692.470 1261.140 1707.170 2255.400 ;
        RECT 1711.070 1261.140 1725.770 2255.400 ;
        RECT 1729.670 1261.140 1744.370 2255.400 ;
        RECT 1748.270 1261.140 1758.570 2255.400 ;
        RECT 1762.470 1261.140 1777.170 2255.400 ;
        RECT 1781.070 2145.095 1795.770 2255.400 ;
        RECT 1799.670 2145.095 1814.370 3501.825 ;
        RECT 1818.270 2145.095 1828.570 3501.825 ;
        RECT 1832.470 2145.095 1847.170 3501.825 ;
        RECT 1851.070 2145.095 1865.770 3501.825 ;
        RECT 1869.670 2145.095 1884.370 3501.825 ;
        RECT 1888.270 3226.140 1898.570 3501.825 ;
        RECT 1902.470 3226.140 1917.170 3501.825 ;
        RECT 1921.070 3226.140 1935.770 3501.825 ;
        RECT 1939.670 3226.140 1954.370 3501.825 ;
        RECT 1958.270 3226.140 1968.570 3501.825 ;
        RECT 1972.470 3226.140 1987.170 3501.825 ;
        RECT 1991.070 3226.140 2005.770 3501.825 ;
        RECT 2009.670 3226.140 2024.370 3501.825 ;
        RECT 2028.270 3226.140 2038.570 3501.825 ;
        RECT 2042.470 3226.140 2057.170 3501.825 ;
        RECT 2061.070 3226.140 2075.770 3501.825 ;
        RECT 2079.670 3226.140 2094.370 3501.825 ;
        RECT 2098.270 3226.140 2108.570 3501.825 ;
        RECT 2112.470 3226.140 2127.170 3501.825 ;
        RECT 2131.070 3226.140 2145.770 3501.825 ;
        RECT 2149.670 3226.140 2164.370 3501.825 ;
        RECT 2168.270 3226.140 2178.570 3501.825 ;
        RECT 2182.470 3226.140 2197.170 3501.825 ;
        RECT 2201.070 3226.140 2215.770 3501.825 ;
        RECT 2219.670 3226.140 2234.370 3501.825 ;
        RECT 2238.270 3226.140 2248.570 3501.825 ;
        RECT 2252.470 3226.140 2267.170 3501.825 ;
        RECT 2271.070 3226.140 2285.770 3501.825 ;
        RECT 2289.670 3226.140 2304.370 3501.825 ;
        RECT 2308.270 3226.140 2318.570 3501.825 ;
        RECT 2322.470 3226.140 2337.170 3501.825 ;
        RECT 2341.070 3226.140 2355.770 3501.825 ;
        RECT 2359.670 3226.140 2374.370 3501.825 ;
        RECT 2378.270 3226.140 2388.570 3501.825 ;
        RECT 2392.470 3226.140 2407.170 3501.825 ;
        RECT 2411.070 3226.140 2425.770 3501.825 ;
        RECT 2429.670 3226.140 2444.370 3501.825 ;
        RECT 2448.270 3226.140 2458.570 3501.825 ;
        RECT 2462.470 3226.140 2477.170 3501.825 ;
        RECT 2481.070 3226.140 2495.770 3501.825 ;
        RECT 2499.670 3226.140 2514.370 3501.825 ;
        RECT 2518.270 3226.140 2528.570 3501.825 ;
        RECT 2532.470 3226.140 2547.170 3501.825 ;
        RECT 2551.070 3226.140 2565.770 3501.825 ;
        RECT 2569.670 3226.140 2582.480 3501.825 ;
        RECT 1888.270 2790.400 2582.480 3226.140 ;
        RECT 1888.270 2691.140 1898.570 2790.400 ;
        RECT 1902.470 2691.140 1917.170 2790.400 ;
        RECT 1921.070 2691.140 1935.770 2790.400 ;
        RECT 1939.670 2691.140 1954.370 2790.400 ;
        RECT 1958.270 2691.140 1968.570 2790.400 ;
        RECT 1972.470 2691.140 1987.170 2790.400 ;
        RECT 1991.070 2691.140 2005.770 2790.400 ;
        RECT 2009.670 2691.140 2024.370 2790.400 ;
        RECT 2028.270 2691.140 2038.570 2790.400 ;
        RECT 2042.470 2691.140 2057.170 2790.400 ;
        RECT 2061.070 2691.140 2075.770 2790.400 ;
        RECT 2079.670 2691.140 2094.370 2790.400 ;
        RECT 2098.270 2691.140 2108.570 2790.400 ;
        RECT 2112.470 2691.140 2127.170 2790.400 ;
        RECT 2131.070 2691.140 2145.770 2790.400 ;
        RECT 2149.670 2691.140 2164.370 2790.400 ;
        RECT 2168.270 2691.140 2178.570 2790.400 ;
        RECT 2182.470 2691.140 2197.170 2790.400 ;
        RECT 2201.070 2691.140 2215.770 2790.400 ;
        RECT 2219.670 2691.140 2234.370 2790.400 ;
        RECT 2238.270 2691.140 2248.570 2790.400 ;
        RECT 2252.470 2691.140 2267.170 2790.400 ;
        RECT 2271.070 2691.140 2285.770 2790.400 ;
        RECT 2289.670 2691.140 2304.370 2790.400 ;
        RECT 2308.270 2691.140 2318.570 2790.400 ;
        RECT 2322.470 2691.140 2337.170 2790.400 ;
        RECT 2341.070 2691.140 2355.770 2790.400 ;
        RECT 2359.670 2691.140 2374.370 2790.400 ;
        RECT 2378.270 2691.140 2388.570 2790.400 ;
        RECT 2392.470 2691.140 2407.170 2790.400 ;
        RECT 2411.070 2691.140 2425.770 2790.400 ;
        RECT 2429.670 2691.140 2444.370 2790.400 ;
        RECT 2448.270 2691.140 2458.570 2790.400 ;
        RECT 2462.470 2691.140 2477.170 2790.400 ;
        RECT 2481.070 2691.140 2495.770 2790.400 ;
        RECT 2499.670 2691.140 2514.370 2790.400 ;
        RECT 2518.270 2691.140 2528.570 2790.400 ;
        RECT 2532.470 2691.140 2547.170 2790.400 ;
        RECT 2551.070 2691.140 2565.770 2790.400 ;
        RECT 2569.670 2691.140 2582.480 2790.400 ;
        RECT 1888.270 2255.400 2582.480 2691.140 ;
        RECT 1888.270 2145.095 1898.570 2255.400 ;
        RECT 1902.470 2145.095 1917.170 2255.400 ;
        RECT 1921.070 2145.095 1935.770 2255.400 ;
        RECT 1939.670 2145.095 1954.370 2255.400 ;
        RECT 1958.270 2145.095 1968.570 2255.400 ;
        RECT 1972.470 2145.095 1987.170 2255.400 ;
        RECT 1991.070 2145.095 2005.770 2255.400 ;
        RECT 2009.670 2145.095 2024.370 2255.400 ;
        RECT 2028.270 2145.095 2038.570 2255.400 ;
        RECT 2042.470 2145.095 2057.170 2255.400 ;
        RECT 2061.070 2145.095 2075.770 2255.400 ;
        RECT 2079.670 2145.095 2094.370 2255.400 ;
        RECT 2098.270 2145.095 2108.570 2255.400 ;
        RECT 2112.470 2145.095 2127.170 2255.400 ;
        RECT 1781.070 1810.400 2127.170 2145.095 ;
        RECT 1781.070 1710.095 1795.770 1810.400 ;
        RECT 1799.670 1710.095 1814.370 1810.400 ;
        RECT 1818.270 1710.095 1828.570 1810.400 ;
        RECT 1832.470 1710.095 1847.170 1810.400 ;
        RECT 1851.070 1710.095 1865.770 1810.400 ;
        RECT 1869.670 1710.095 1884.370 1810.400 ;
        RECT 1888.270 1710.095 1898.570 1810.400 ;
        RECT 1902.470 1710.095 1917.170 1810.400 ;
        RECT 1921.070 1710.095 1935.770 1810.400 ;
        RECT 1939.670 1710.095 1954.370 1810.400 ;
        RECT 1958.270 1710.095 1968.570 1810.400 ;
        RECT 1972.470 1710.095 1987.170 1810.400 ;
        RECT 1991.070 1710.095 2005.770 1810.400 ;
        RECT 2009.670 1710.095 2024.370 1810.400 ;
        RECT 2028.270 1710.095 2038.570 1810.400 ;
        RECT 2042.470 1710.095 2057.170 1810.400 ;
        RECT 2061.070 1710.095 2075.770 1810.400 ;
        RECT 2079.670 1710.095 2094.370 1810.400 ;
        RECT 2098.270 1710.095 2108.570 1810.400 ;
        RECT 2112.470 1710.095 2127.170 1810.400 ;
        RECT 1781.070 1375.400 2127.170 1710.095 ;
        RECT 1781.070 1261.140 1795.770 1375.400 ;
        RECT 1081.070 825.400 1795.770 1261.140 ;
        RECT 1081.070 726.140 1095.770 825.400 ;
        RECT 1099.670 726.140 1114.370 825.400 ;
        RECT 1118.270 726.140 1128.570 825.400 ;
        RECT 1132.470 726.140 1147.170 825.400 ;
        RECT 1151.070 726.140 1165.770 825.400 ;
        RECT 1169.670 726.140 1184.370 825.400 ;
        RECT 1188.270 726.140 1198.570 825.400 ;
        RECT 1202.470 726.140 1217.170 825.400 ;
        RECT 1221.070 726.140 1235.770 825.400 ;
        RECT 1239.670 726.140 1254.370 825.400 ;
        RECT 1258.270 726.140 1268.570 825.400 ;
        RECT 1272.470 726.140 1287.170 825.400 ;
        RECT 1291.070 726.140 1305.770 825.400 ;
        RECT 1309.670 726.140 1324.370 825.400 ;
        RECT 1328.270 726.140 1338.570 825.400 ;
        RECT 1342.470 726.140 1357.170 825.400 ;
        RECT 1361.070 726.140 1375.770 825.400 ;
        RECT 1379.670 726.140 1394.370 825.400 ;
        RECT 1398.270 726.140 1408.570 825.400 ;
        RECT 1412.470 726.140 1427.170 825.400 ;
        RECT 1431.070 726.140 1445.770 825.400 ;
        RECT 1449.670 726.140 1464.370 825.400 ;
        RECT 1468.270 726.140 1478.570 825.400 ;
        RECT 1482.470 726.140 1497.170 825.400 ;
        RECT 1501.070 726.140 1515.770 825.400 ;
        RECT 1519.670 726.140 1534.370 825.400 ;
        RECT 1538.270 726.140 1548.570 825.400 ;
        RECT 1552.470 726.140 1567.170 825.400 ;
        RECT 1571.070 726.140 1585.770 825.400 ;
        RECT 1589.670 726.140 1604.370 825.400 ;
        RECT 1608.270 726.140 1618.570 825.400 ;
        RECT 1622.470 726.140 1637.170 825.400 ;
        RECT 1641.070 726.140 1655.770 825.400 ;
        RECT 1659.670 726.140 1674.370 825.400 ;
        RECT 1678.270 726.140 1688.570 825.400 ;
        RECT 1692.470 726.140 1707.170 825.400 ;
        RECT 1711.070 726.140 1725.770 825.400 ;
        RECT 1729.670 726.140 1744.370 825.400 ;
        RECT 1748.270 726.140 1758.570 825.400 ;
        RECT 1762.470 726.140 1777.170 825.400 ;
        RECT 1781.070 726.140 1795.770 825.400 ;
        RECT 1081.070 290.400 1795.770 726.140 ;
        RECT 1081.070 57.975 1095.770 290.400 ;
        RECT 1099.670 57.975 1114.370 290.400 ;
        RECT 1118.270 57.975 1128.570 290.400 ;
        RECT 1132.470 57.975 1147.170 290.400 ;
        RECT 1151.070 57.975 1165.770 290.400 ;
        RECT 1169.670 57.975 1184.370 290.400 ;
        RECT 1188.270 57.975 1198.570 290.400 ;
        RECT 1202.470 57.975 1217.170 290.400 ;
        RECT 1221.070 57.975 1235.770 290.400 ;
        RECT 1239.670 57.975 1254.370 290.400 ;
        RECT 1258.270 57.975 1268.570 290.400 ;
        RECT 1272.470 57.975 1287.170 290.400 ;
        RECT 1291.070 57.975 1305.770 290.400 ;
        RECT 1309.670 57.975 1324.370 290.400 ;
        RECT 1328.270 57.975 1338.570 290.400 ;
        RECT 1342.470 57.975 1357.170 290.400 ;
        RECT 1361.070 57.975 1375.770 290.400 ;
        RECT 1379.670 57.975 1394.370 290.400 ;
        RECT 1398.270 57.975 1408.570 290.400 ;
        RECT 1412.470 57.975 1427.170 290.400 ;
        RECT 1431.070 57.975 1445.770 290.400 ;
        RECT 1449.670 57.975 1464.370 290.400 ;
        RECT 1468.270 57.975 1478.570 290.400 ;
        RECT 1482.470 57.975 1497.170 290.400 ;
        RECT 1501.070 57.975 1515.770 290.400 ;
        RECT 1519.670 57.975 1534.370 290.400 ;
        RECT 1538.270 57.975 1548.570 290.400 ;
        RECT 1552.470 57.975 1567.170 290.400 ;
        RECT 1571.070 57.975 1585.770 290.400 ;
        RECT 1589.670 57.975 1604.370 290.400 ;
        RECT 1608.270 57.975 1618.570 290.400 ;
        RECT 1622.470 57.975 1637.170 290.400 ;
        RECT 1641.070 57.975 1655.770 290.400 ;
        RECT 1659.670 57.975 1674.370 290.400 ;
        RECT 1678.270 57.975 1688.570 290.400 ;
        RECT 1692.470 57.975 1707.170 290.400 ;
        RECT 1711.070 57.975 1725.770 290.400 ;
        RECT 1729.670 57.975 1744.370 290.400 ;
        RECT 1748.270 57.975 1758.570 290.400 ;
        RECT 1762.470 57.975 1777.170 290.400 ;
        RECT 1781.070 57.975 1795.770 290.400 ;
        RECT 1799.670 57.975 1814.370 1375.400 ;
        RECT 1818.270 57.975 1828.570 1375.400 ;
        RECT 1832.470 57.975 1847.170 1375.400 ;
        RECT 1851.070 57.975 1865.770 1375.400 ;
        RECT 1869.670 57.975 1884.370 1375.400 ;
        RECT 1888.270 1261.140 1898.570 1375.400 ;
        RECT 1902.470 1261.140 1917.170 1375.400 ;
        RECT 1921.070 1261.140 1935.770 1375.400 ;
        RECT 1939.670 1261.140 1954.370 1375.400 ;
        RECT 1958.270 1261.140 1968.570 1375.400 ;
        RECT 1972.470 1261.140 1987.170 1375.400 ;
        RECT 1991.070 1261.140 2005.770 1375.400 ;
        RECT 2009.670 1261.140 2024.370 1375.400 ;
        RECT 2028.270 1261.140 2038.570 1375.400 ;
        RECT 2042.470 1261.140 2057.170 1375.400 ;
        RECT 2061.070 1261.140 2075.770 1375.400 ;
        RECT 2079.670 1261.140 2094.370 1375.400 ;
        RECT 2098.270 1261.140 2108.570 1375.400 ;
        RECT 2112.470 1261.140 2127.170 1375.400 ;
        RECT 2131.070 1261.140 2145.770 2255.400 ;
        RECT 2149.670 1261.140 2164.370 2255.400 ;
        RECT 2168.270 1261.140 2178.570 2255.400 ;
        RECT 2182.470 1261.140 2197.170 2255.400 ;
        RECT 2201.070 1261.140 2215.770 2255.400 ;
        RECT 2219.670 1261.140 2234.370 2255.400 ;
        RECT 2238.270 2145.095 2248.570 2255.400 ;
        RECT 2252.470 2145.095 2267.170 2255.400 ;
        RECT 2271.070 2145.095 2285.770 2255.400 ;
        RECT 2289.670 2145.095 2304.370 2255.400 ;
        RECT 2308.270 2145.095 2318.570 2255.400 ;
        RECT 2322.470 2145.095 2337.170 2255.400 ;
        RECT 2341.070 2145.095 2355.770 2255.400 ;
        RECT 2359.670 2145.095 2374.370 2255.400 ;
        RECT 2378.270 2145.095 2388.570 2255.400 ;
        RECT 2392.470 2145.095 2407.170 2255.400 ;
        RECT 2411.070 2145.095 2425.770 2255.400 ;
        RECT 2429.670 2145.095 2444.370 2255.400 ;
        RECT 2448.270 2145.095 2458.570 2255.400 ;
        RECT 2462.470 2145.095 2477.170 2255.400 ;
        RECT 2481.070 2145.095 2495.770 2255.400 ;
        RECT 2499.670 2145.095 2514.370 2255.400 ;
        RECT 2518.270 2145.095 2528.570 2255.400 ;
        RECT 2532.470 2145.095 2547.170 2255.400 ;
        RECT 2551.070 2145.095 2565.770 2255.400 ;
        RECT 2238.270 1810.400 2565.770 2145.095 ;
        RECT 2238.270 1261.140 2248.570 1810.400 ;
        RECT 2252.470 1261.140 2267.170 1810.400 ;
        RECT 2271.070 1261.140 2285.770 1810.400 ;
        RECT 2289.670 1644.600 2304.370 1810.400 ;
        RECT 2308.270 1644.600 2318.570 1810.400 ;
        RECT 2322.470 1644.600 2337.170 1810.400 ;
        RECT 2341.070 1644.600 2355.770 1810.400 ;
        RECT 2359.670 1644.600 2374.370 1810.400 ;
        RECT 2378.270 1644.600 2388.570 1810.400 ;
        RECT 2392.470 1644.600 2407.170 1810.400 ;
        RECT 2411.070 1644.600 2425.770 1810.400 ;
        RECT 2429.670 1644.600 2444.370 1810.400 ;
        RECT 2448.270 1644.600 2458.570 1810.400 ;
        RECT 2462.470 1644.600 2477.170 1810.400 ;
        RECT 2481.070 1644.600 2495.770 1810.400 ;
        RECT 2499.670 1644.600 2514.370 1810.400 ;
        RECT 2518.270 1644.600 2528.570 1810.400 ;
        RECT 2532.470 1644.600 2547.170 1810.400 ;
        RECT 2551.070 1644.600 2565.770 1810.400 ;
        RECT 2289.670 1375.400 2565.770 1644.600 ;
        RECT 2289.670 1261.140 2304.370 1375.400 ;
        RECT 2308.270 1261.140 2318.570 1375.400 ;
        RECT 2322.470 1261.140 2337.170 1375.400 ;
        RECT 2341.070 1261.140 2355.770 1375.400 ;
        RECT 2359.670 1261.140 2374.370 1375.400 ;
        RECT 2378.270 1261.140 2388.570 1375.400 ;
        RECT 2392.470 1261.140 2407.170 1375.400 ;
        RECT 2411.070 1261.140 2425.770 1375.400 ;
        RECT 2429.670 1261.140 2444.370 1375.400 ;
        RECT 2448.270 1261.140 2458.570 1375.400 ;
        RECT 2462.470 1261.140 2477.170 1375.400 ;
        RECT 2481.070 1261.140 2495.770 1375.400 ;
        RECT 2499.670 1261.140 2514.370 1375.400 ;
        RECT 2518.270 1261.140 2528.570 1375.400 ;
        RECT 2532.470 1261.140 2547.170 1375.400 ;
        RECT 2551.070 1261.140 2565.770 1375.400 ;
        RECT 2569.670 1261.140 2582.480 2255.400 ;
        RECT 1888.270 825.400 2582.480 1261.140 ;
        RECT 1888.270 726.140 1898.570 825.400 ;
        RECT 1902.470 726.140 1917.170 825.400 ;
        RECT 1921.070 726.140 1935.770 825.400 ;
        RECT 1939.670 726.140 1954.370 825.400 ;
        RECT 1958.270 726.140 1968.570 825.400 ;
        RECT 1972.470 726.140 1987.170 825.400 ;
        RECT 1991.070 726.140 2005.770 825.400 ;
        RECT 2009.670 726.140 2024.370 825.400 ;
        RECT 2028.270 726.140 2038.570 825.400 ;
        RECT 2042.470 726.140 2057.170 825.400 ;
        RECT 2061.070 726.140 2075.770 825.400 ;
        RECT 2079.670 726.140 2094.370 825.400 ;
        RECT 2098.270 726.140 2108.570 825.400 ;
        RECT 2112.470 726.140 2127.170 825.400 ;
        RECT 2131.070 726.140 2145.770 825.400 ;
        RECT 2149.670 726.140 2164.370 825.400 ;
        RECT 2168.270 726.140 2178.570 825.400 ;
        RECT 2182.470 726.140 2197.170 825.400 ;
        RECT 2201.070 726.140 2215.770 825.400 ;
        RECT 2219.670 726.140 2234.370 825.400 ;
        RECT 2238.270 726.140 2248.570 825.400 ;
        RECT 2252.470 726.140 2267.170 825.400 ;
        RECT 2271.070 726.140 2285.770 825.400 ;
        RECT 2289.670 726.140 2304.370 825.400 ;
        RECT 2308.270 726.140 2318.570 825.400 ;
        RECT 2322.470 726.140 2337.170 825.400 ;
        RECT 2341.070 726.140 2355.770 825.400 ;
        RECT 2359.670 726.140 2374.370 825.400 ;
        RECT 2378.270 726.140 2388.570 825.400 ;
        RECT 2392.470 726.140 2407.170 825.400 ;
        RECT 2411.070 726.140 2425.770 825.400 ;
        RECT 2429.670 726.140 2444.370 825.400 ;
        RECT 2448.270 726.140 2458.570 825.400 ;
        RECT 2462.470 726.140 2477.170 825.400 ;
        RECT 2481.070 726.140 2495.770 825.400 ;
        RECT 2499.670 726.140 2514.370 825.400 ;
        RECT 2518.270 726.140 2528.570 825.400 ;
        RECT 2532.470 726.140 2547.170 825.400 ;
        RECT 2551.070 726.140 2565.770 825.400 ;
        RECT 2569.670 726.140 2582.480 825.400 ;
        RECT 1888.270 290.400 2582.480 726.140 ;
        RECT 1888.270 57.975 1898.570 290.400 ;
        RECT 1902.470 57.975 1917.170 290.400 ;
        RECT 1921.070 57.975 1935.770 290.400 ;
        RECT 1939.670 57.975 1954.370 290.400 ;
        RECT 1958.270 57.975 1968.570 290.400 ;
        RECT 1972.470 57.975 1987.170 290.400 ;
        RECT 1991.070 57.975 2005.770 290.400 ;
        RECT 2009.670 57.975 2024.370 290.400 ;
        RECT 2028.270 57.975 2038.570 290.400 ;
        RECT 2042.470 57.975 2057.170 290.400 ;
        RECT 2061.070 57.975 2075.770 290.400 ;
        RECT 2079.670 57.975 2094.370 290.400 ;
        RECT 2098.270 57.975 2108.570 290.400 ;
        RECT 2112.470 57.975 2127.170 290.400 ;
        RECT 2131.070 57.975 2145.770 290.400 ;
        RECT 2149.670 57.975 2164.370 290.400 ;
        RECT 2168.270 57.975 2178.570 290.400 ;
        RECT 2182.470 57.975 2197.170 290.400 ;
        RECT 2201.070 57.975 2215.770 290.400 ;
        RECT 2219.670 57.975 2234.370 290.400 ;
        RECT 2238.270 57.975 2248.570 290.400 ;
        RECT 2252.470 57.975 2267.170 290.400 ;
        RECT 2271.070 57.975 2285.770 290.400 ;
        RECT 2289.670 57.975 2304.370 290.400 ;
        RECT 2308.270 57.975 2318.570 290.400 ;
        RECT 2322.470 57.975 2337.170 290.400 ;
        RECT 2341.070 57.975 2355.770 290.400 ;
        RECT 2359.670 57.975 2374.370 290.400 ;
        RECT 2378.270 57.975 2388.570 290.400 ;
        RECT 2392.470 57.975 2407.170 290.400 ;
        RECT 2411.070 57.975 2425.770 290.400 ;
        RECT 2429.670 57.975 2444.370 290.400 ;
        RECT 2448.270 57.975 2458.570 290.400 ;
        RECT 2462.470 57.975 2477.170 290.400 ;
        RECT 2481.070 57.975 2495.770 290.400 ;
        RECT 2499.670 57.975 2514.370 290.400 ;
        RECT 2518.270 57.975 2528.570 290.400 ;
        RECT 2532.470 57.975 2547.170 290.400 ;
        RECT 2551.070 57.975 2565.770 290.400 ;
        RECT 2569.670 57.975 2582.480 290.400 ;
  END
END user_project_wrapper
END LIBRARY

